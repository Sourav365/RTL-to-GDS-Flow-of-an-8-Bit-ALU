NAMESCASESENSITIVE ON ;
MACRO AN2
    CLASS CORE ;
    FOREIGN AN2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 2.790 2.310 3.190 ;
        RECT  2.030 1.180 2.310 3.300 ;
        RECT  2.000 1.380 2.310 1.780 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.110 2.650 ;
        RECT  0.790 2.100 1.070 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.650 0.550 2.180 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  1.340 -0.380 1.740 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.410 4.090 1.810 5.420 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.470 4.130 0.870 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.470 3.410 1.760 3.650 ;
        RECT  1.520 1.080 1.760 3.650 ;
        RECT  1.520 2.250 1.790 2.650 ;
        RECT  0.160 1.080 1.760 1.320 ;
    END
END AN2

MACRO AN2B1
    CLASS CORE ;
    FOREIGN AN2B1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.340 3.100 2.930 3.340 ;
        RECT  1.600 1.180 3.460 1.420 ;
        RECT  2.650 1.180 2.930 3.340 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.300 1.070 2.940 ;
        RECT  0.720 2.300 1.070 2.700 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.670 2.480 1.950 3.920 ;
        RECT  3.690 2.370 4.170 2.770 ;
        RECT  3.890 2.300 4.170 3.920 ;
        RECT  1.670 3.640 4.170 3.920 ;
        RECT  1.490 2.480 1.950 2.880 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.330 -0.380 2.730 0.820 ;
        RECT  3.780 -0.380 4.180 1.290 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.880 -0.380 1.280 1.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 4.160 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.880 3.910 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.620 4.160 3.460 4.400 ;
        RECT  0.190 3.670 0.480 4.070 ;
        RECT  0.190 1.100 0.430 4.070 ;
        RECT  2.170 1.810 2.410 2.210 ;
        RECT  0.190 1.810 2.410 2.050 ;
        RECT  0.190 1.100 0.480 1.500 ;
    END
END AN2B1

MACRO AN2B1P
    CLASS CORE ;
    FOREIGN AN2B1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.760 2.900 4.170 3.300 ;
        RECT  3.150 1.530 4.800 1.810 ;
        RECT  3.890 1.530 4.170 3.300 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.350 2.100 1.690 2.500 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.660 1.070 3.300 ;
        RECT  0.670 2.660 1.070 3.060 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 -0.380 4.180 1.020 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.020 -0.380 1.420 1.130 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 4.480 3.060 5.420 ;
        RECT  4.400 4.180 4.800 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  1.020 3.910 1.420 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.850 3.910 2.910 4.150 ;
        RECT  2.670 0.810 2.910 4.150 ;
        RECT  2.670 2.130 3.650 2.530 ;
        RECT  2.510 0.810 2.910 1.210 ;
        RECT  0.190 3.670 0.480 4.070 ;
        RECT  0.190 0.810 0.430 4.070 ;
        RECT  1.930 1.370 2.330 1.690 ;
        RECT  0.190 1.370 2.330 1.610 ;
        RECT  0.190 0.810 0.480 1.610 ;
    END
END AN2B1P

MACRO AN2B1S
    CLASS CORE ;
    FOREIGN AN2B1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.100 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.070 2.310 2.100 ;
        RECT  2.030 1.820 2.930 2.100 ;
        RECT  2.650 1.820 2.930 3.420 ;
        RECT  2.620 3.020 2.930 3.420 ;
        RECT  1.860 1.070 2.310 1.470 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.610 1.070 2.250 ;
        RECT  0.720 1.610 1.070 2.010 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.320 1.700 2.720 ;
        RECT  1.410 2.300 1.690 2.940 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.550 -0.380 2.940 1.210 ;
        RECT  0.000 -0.380 3.100 0.380 ;
        RECT  1.020 -0.380 1.420 1.230 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.100 5.420 ;
        RECT  1.010 4.480 1.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.190 4.000 2.380 4.240 ;
        RECT  2.140 2.480 2.380 4.240 ;
        RECT  0.190 3.830 0.480 4.240 ;
        RECT  0.190 1.070 0.430 4.240 ;
        RECT  2.140 2.480 2.410 2.880 ;
        RECT  0.190 1.070 0.480 1.470 ;
    END
END AN2B1S

MACRO AN2B1T
    CLASS CORE ;
    FOREIGN AN2B1T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.750 1.490 5.310 3.280 ;
        RECT  3.610 2.880 5.310 3.280 ;
        RECT  3.610 1.490 5.310 1.890 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.200 2.630 2.600 ;
        RECT  2.030 2.200 2.310 2.840 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.450 1.070 3.400 ;
        RECT  0.740 2.450 1.070 2.850 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.740 -0.380 3.140 0.560 ;
        RECT  4.260 -0.380 4.660 1.120 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.380 -0.380 0.780 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.910 4.260 3.310 5.420 ;
        RECT  4.260 4.180 4.660 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  1.400 3.750 1.800 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.120 3.780 3.370 4.020 ;
        RECT  3.130 0.890 3.370 4.020 ;
        RECT  3.130 2.170 3.510 2.570 ;
        RECT  1.400 0.890 3.370 1.130 ;
        RECT  0.240 1.370 0.480 3.390 ;
        RECT  1.430 1.370 1.670 2.310 ;
        RECT  0.240 1.370 1.670 1.610 ;
    END
END AN2B1T

MACRO AN2P
    CLASS CORE ;
    FOREIGN AN2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.520 2.790 2.930 3.190 ;
        RECT  2.650 1.180 2.930 3.300 ;
        RECT  2.520 1.320 2.930 1.720 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.360 2.250 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.540 0.530 1.940 ;
        RECT  0.170 1.540 0.450 2.180 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.160 -0.380 3.560 0.780 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  1.670 -0.380 2.070 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 4.260 2.070 5.420 ;
        RECT  3.160 4.260 3.560 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.160 3.780 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.780 2.280 4.020 ;
        RECT  2.040 1.020 2.280 4.020 ;
        RECT  0.160 1.020 2.280 1.260 ;
    END
END AN2P

MACRO AN2S
    CLASS CORE ;
    FOREIGN AN2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.300 2.310 3.400 ;
        RECT  2.000 3.000 2.310 3.400 ;
        RECT  2.000 1.300 2.310 1.700 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.540 1.070 3.300 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.840 0.490 2.240 ;
        RECT  0.170 1.740 0.450 2.380 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.900 -0.380 1.300 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.780 4.100 2.180 5.420 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.450 4.480 0.850 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.450 3.540 1.760 3.780 ;
        RECT  1.520 0.800 1.760 3.780 ;
        RECT  1.520 2.140 1.770 2.540 ;
        RECT  0.320 0.800 1.760 1.040 ;
        RECT  0.160 0.620 0.560 0.860 ;
    END
END AN2S

MACRO AN2T
    CLASS CORE ;
    FOREIGN AN2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.510 1.490 4.070 3.280 ;
        RECT  2.480 2.880 4.070 3.280 ;
        RECT  2.480 1.490 4.070 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.530 1.690 3.300 ;
        RECT  1.190 2.530 1.690 2.930 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.530 2.500 ;
        RECT  0.170 1.740 0.450 2.500 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.020 -0.380 3.420 1.120 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  1.540 -0.380 1.940 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 4.260 2.070 5.420 ;
        RECT  3.020 4.180 3.420 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.160 3.910 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.780 2.240 4.020 ;
        RECT  2.000 0.890 2.240 4.020 ;
        RECT  2.000 2.170 2.270 2.570 ;
        RECT  0.160 0.890 2.240 1.130 ;
    END
END AN2T

MACRO AN3
    CLASS CORE ;
    FOREIGN AN3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.240 2.790 3.550 3.190 ;
        RECT  3.270 1.180 3.550 3.300 ;
        RECT  3.240 1.490 3.550 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.540 1.690 2.180 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.300 0.530 2.700 ;
        RECT  0.170 2.300 0.450 2.940 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 2.940 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  2.370 -0.380 2.770 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.190 4.480 2.590 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.920 4.130 1.320 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.370 2.910 3.610 ;
        RECT  2.670 0.900 2.910 3.610 ;
        RECT  2.670 2.140 3.030 2.540 ;
        RECT  0.160 0.900 2.910 1.140 ;
        RECT  0.160 0.890 0.560 1.140 ;
    END
END AN3

MACRO AN3B1
    CLASS CORE ;
    FOREIGN AN3B1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 2.790 4.790 3.190 ;
        RECT  4.510 1.180 4.790 3.300 ;
        RECT  4.480 1.490 4.790 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.640 1.690 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.840 2.310 3.480 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.840 1.070 3.480 ;
        RECT  0.670 2.840 1.070 3.240 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 -0.380 4.010 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.130 4.480 2.530 5.420 ;
        RECT  3.680 4.260 4.080 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.540 3.720 4.150 3.960 ;
        RECT  3.910 1.020 4.150 3.960 ;
        RECT  3.030 1.020 4.150 1.260 ;
        RECT  3.030 0.860 3.270 1.260 ;
        RECT  0.190 3.570 0.480 3.970 ;
        RECT  0.190 0.940 0.430 3.970 ;
        RECT  2.550 1.500 3.030 1.740 ;
        RECT  2.550 0.940 2.790 1.740 ;
        RECT  0.160 0.940 2.790 1.180 ;
    END
END AN3B1

MACRO AN3B1P
    CLASS CORE ;
    FOREIGN AN3B1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.450 2.790 4.790 3.190 ;
        RECT  4.510 1.180 4.790 3.300 ;
        RECT  4.450 1.320 4.790 1.720 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.640 1.690 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.820 2.310 3.460 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.820 1.070 3.460 ;
        RECT  0.670 2.820 1.070 3.220 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.710 -0.380 4.110 0.860 ;
        RECT  5.020 -0.380 5.420 0.860 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 4.480 2.600 5.420 ;
        RECT  3.710 4.180 4.110 5.420 ;
        RECT  5.020 4.180 5.420 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  1.020 4.480 1.420 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.610 3.700 4.150 3.940 ;
        RECT  3.910 1.100 4.150 3.940 ;
        RECT  3.070 1.100 4.150 1.340 ;
        RECT  3.070 0.940 3.310 1.340 ;
        RECT  0.190 3.580 0.480 3.980 ;
        RECT  0.190 1.020 0.430 3.980 ;
        RECT  2.590 1.580 3.340 1.820 ;
        RECT  2.590 1.020 2.830 1.820 ;
        RECT  0.160 1.020 2.830 1.260 ;
    END
END AN3B1P

MACRO AN3B1S
    CLASS CORE ;
    FOREIGN AN3B1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.060 4.790 3.710 ;
        RECT  4.480 3.310 4.790 3.710 ;
        RECT  4.480 1.060 4.790 1.460 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.540 1.690 2.180 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 2.940 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.670 2.540 1.070 2.940 ;
        RECT  0.790 2.300 1.070 2.940 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.790 -0.380 4.190 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.610 4.480 2.010 5.420 ;
        RECT  2.270 4.480 2.670 5.420 ;
        RECT  3.610 4.480 4.010 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.540 3.330 4.150 3.570 ;
        RECT  3.910 1.020 4.150 3.570 ;
        RECT  3.150 1.020 4.150 1.260 ;
        RECT  3.150 0.860 3.390 1.260 ;
        RECT  0.190 3.250 0.480 3.650 ;
        RECT  0.190 0.800 0.430 3.650 ;
        RECT  2.670 1.500 3.070 1.740 ;
        RECT  2.670 0.800 2.910 1.740 ;
        RECT  0.160 0.940 0.560 1.180 ;
        RECT  0.190 0.800 2.910 1.040 ;
    END
END AN3B1S

MACRO AN3B1T
    CLASS CORE ;
    FOREIGN AN3B1T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.350 2.870 4.590 3.270 ;
        RECT  5.130 1.400 5.410 3.110 ;
        RECT  4.350 1.400 6.040 1.640 ;
        RECT  4.350 2.870 6.040 3.110 ;
        RECT  4.350 1.240 4.590 1.640 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.880 1.690 2.750 ;
        RECT  1.350 1.880 1.690 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.220 2.310 2.860 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.220 1.070 2.860 ;
        RECT  0.670 2.220 1.070 2.620 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.640 -0.380 4.040 0.860 ;
        RECT  5.020 -0.380 5.420 0.860 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.750 -0.380 1.150 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.130 4.480 2.530 5.420 ;
        RECT  3.640 4.180 4.040 5.420 ;
        RECT  5.020 4.180 5.420 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.750 4.480 1.150 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.540 3.440 4.080 3.680 ;
        RECT  3.840 1.100 4.080 3.680 ;
        RECT  3.000 1.100 4.080 1.340 ;
        RECT  3.000 0.940 3.240 1.340 ;
        RECT  0.190 3.020 0.480 3.420 ;
        RECT  0.190 1.220 0.430 3.420 ;
        RECT  2.500 1.820 3.090 2.060 ;
        RECT  2.500 1.220 2.740 2.060 ;
        RECT  0.160 1.280 0.560 1.520 ;
        RECT  0.190 1.220 2.740 1.460 ;
    END
END AN3B1T

MACRO AN3B2
    CLASS CORE ;
    FOREIGN AN3B2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.100 2.790 5.410 3.190 ;
        RECT  5.130 1.180 5.410 3.300 ;
        RECT  5.100 1.490 5.410 1.890 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.220 1.540 1.690 1.940 ;
        RECT  1.410 0.960 1.690 1.940 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.760 1.070 3.400 ;
        RECT  0.710 2.760 1.070 3.160 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.100 4.170 2.740 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.130 -0.380 4.530 0.560 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.230 4.480 2.630 5.420 ;
        RECT  4.250 4.480 4.650 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.750 4.480 1.150 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.620 4.000 4.770 4.240 ;
        RECT  4.530 0.800 4.770 4.240 ;
        RECT  3.000 3.640 3.240 4.240 ;
        RECT  1.620 3.640 1.860 4.240 ;
        RECT  4.530 2.140 4.870 2.540 ;
        RECT  2.650 0.800 4.770 1.040 ;
        RECT  3.050 1.490 3.290 3.190 ;
        RECT  2.950 2.030 3.290 2.430 ;
        RECT  3.050 1.490 3.340 1.890 ;
        RECT  0.190 3.580 0.480 3.980 ;
        RECT  0.190 0.860 0.430 3.980 ;
        RECT  0.190 2.280 2.130 2.520 ;
        RECT  0.190 0.860 0.480 1.260 ;
    END
END AN3B2

MACRO AN3B2P
    CLASS CORE ;
    FOREIGN AN3B2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.100 2.790 5.410 3.190 ;
        RECT  5.130 1.180 5.410 3.300 ;
        RECT  5.100 1.490 5.410 1.890 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 1.540 1.690 1.940 ;
        RECT  1.410 1.180 1.690 1.940 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.760 1.070 3.400 ;
        RECT  0.710 2.760 1.070 3.160 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.100 4.170 2.740 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.130 -0.380 4.530 0.560 ;
        RECT  5.640 -0.380 6.040 1.070 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.330 4.480 2.730 5.420 ;
        RECT  4.400 4.220 4.800 5.420 ;
        RECT  5.640 4.220 6.040 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.750 4.480 1.150 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.540 3.660 4.770 3.900 ;
        RECT  4.530 0.800 4.770 3.900 ;
        RECT  4.530 2.140 4.870 2.540 ;
        RECT  2.670 0.800 4.770 1.040 ;
        RECT  3.290 1.490 3.530 3.190 ;
        RECT  3.050 2.100 3.530 2.500 ;
        RECT  0.190 3.580 0.480 3.980 ;
        RECT  0.190 0.930 0.430 3.980 ;
        RECT  0.190 2.280 2.310 2.520 ;
        RECT  0.190 0.930 0.480 1.330 ;
    END
END AN3B2P

MACRO AN3B2S
    CLASS CORE ;
    FOREIGN AN3B2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.120 3.550 3.300 ;
        RECT  3.240 2.900 3.550 3.300 ;
        RECT  1.600 1.140 3.560 1.380 ;
        RECT  1.600 1.120 3.550 1.400 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.690 1.070 2.330 ;
        RECT  0.720 1.690 1.070 2.090 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.690 2.350 2.090 ;
        RECT  2.030 1.690 2.310 2.330 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.370 -0.380 2.770 0.560 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.880 -0.380 1.280 1.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  1.040 4.260 1.440 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.190 3.780 3.000 4.020 ;
        RECT  2.760 2.250 3.000 4.020 ;
        RECT  0.190 3.620 0.480 4.020 ;
        RECT  0.190 1.060 0.430 4.020 ;
        RECT  2.760 2.250 3.030 2.650 ;
        RECT  0.190 1.060 0.480 1.460 ;
    END
END AN3B2S

MACRO AN3B2T
    CLASS CORE ;
    FOREIGN AN3B2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.100 2.870 5.340 3.270 ;
        RECT  5.750 1.570 6.030 3.110 ;
        RECT  5.100 1.570 6.660 1.810 ;
        RECT  5.100 2.870 6.660 3.110 ;
        RECT  5.100 1.410 5.340 1.810 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 1.540 1.690 1.940 ;
        RECT  1.410 1.180 1.690 1.940 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.660 1.070 3.400 ;
        RECT  0.710 2.660 1.070 3.060 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.880 4.170 2.520 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.130 -0.380 4.530 0.560 ;
        RECT  5.640 -0.380 6.040 1.070 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.330 4.480 2.730 5.420 ;
        RECT  4.400 4.220 4.800 5.420 ;
        RECT  5.640 4.220 6.040 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  0.750 4.480 1.150 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.540 3.660 4.770 3.900 ;
        RECT  4.530 0.820 4.770 3.900 ;
        RECT  4.530 2.140 4.870 2.540 ;
        RECT  2.670 0.820 4.770 1.060 ;
        RECT  3.290 2.870 4.010 3.110 ;
        RECT  3.290 1.490 3.530 3.110 ;
        RECT  3.050 2.100 3.530 2.500 ;
        RECT  0.190 3.580 0.480 3.980 ;
        RECT  0.190 0.930 0.430 3.980 ;
        RECT  0.190 2.180 2.310 2.420 ;
        RECT  0.190 0.930 0.480 1.330 ;
    END
END AN3B2T

MACRO AN3P
    CLASS CORE ;
    FOREIGN AN3P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.140 2.790 3.550 3.190 ;
        RECT  3.270 1.180 3.550 3.300 ;
        RECT  3.140 1.490 3.550 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.300 1.690 2.940 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.540 0.530 1.940 ;
        RECT  0.170 1.540 0.450 2.180 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.540 2.310 2.180 ;
        RECT  1.980 1.540 2.310 1.940 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 -0.380 4.180 0.950 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  2.150 -0.380 2.550 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.330 4.260 2.730 5.420 ;
        RECT  3.780 4.260 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.850 4.130 1.250 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.360 2.900 3.600 ;
        RECT  2.660 0.890 2.900 3.600 ;
        RECT  0.160 0.890 2.900 1.130 ;
    END
END AN3P

MACRO AN3S
    CLASS CORE ;
    FOREIGN AN3S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 0.620 3.550 3.850 ;
        RECT  3.240 3.450 3.550 3.850 ;
        RECT  3.240 0.670 3.550 1.070 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.540 1.690 2.180 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.550 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  2.370 -0.380 2.770 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.370 4.130 2.770 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.920 4.130 1.320 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.370 2.910 3.610 ;
        RECT  2.670 0.800 2.910 3.610 ;
        RECT  2.670 2.140 3.030 2.540 ;
        RECT  0.160 0.800 0.560 1.130 ;
        RECT  0.160 0.800 2.910 1.040 ;
    END
END AN3S

MACRO AN3T
    CLASS CORE ;
    FOREIGN AN3T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.040 2.870 3.280 3.270 ;
        RECT  3.890 1.570 4.170 3.110 ;
        RECT  3.040 1.570 4.800 1.810 ;
        RECT  3.040 2.870 4.800 3.110 ;
        RECT  3.040 1.410 3.280 1.810 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.090 1.690 2.790 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.620 0.530 2.020 ;
        RECT  0.170 1.620 0.450 2.260 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.620 2.310 2.260 ;
        RECT  1.930 1.620 2.310 2.020 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.680 -0.380 4.080 0.950 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  2.150 -0.380 2.550 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 4.260 2.640 5.420 ;
        RECT  3.680 4.260 4.080 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.850 4.130 1.250 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.360 2.790 3.600 ;
        RECT  2.550 0.890 2.790 3.600 ;
        RECT  2.550 2.140 3.400 2.540 ;
        RECT  0.160 0.890 2.790 1.130 ;
    END
END AN3T

MACRO AN4
    CLASS CORE ;
    FOREIGN AN4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 1.420 5.410 3.260 ;
        RECT  4.500 2.860 5.410 3.260 ;
        RECT  4.800 1.420 5.410 1.660 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.400 1.260 2.800 ;
        RECT  0.790 2.160 1.070 2.800 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.910 0.500 2.310 ;
        RECT  0.170 1.540 0.450 2.310 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.930 1.910 2.310 2.310 ;
        RECT  2.030 1.540 2.310 2.310 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.160 2.930 2.800 ;
        RECT  2.610 2.260 2.930 2.660 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.910 -0.380 4.310 0.560 ;
        RECT  5.640 -0.380 6.040 0.810 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  1.450 -0.380 1.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.920 4.480 3.320 5.420 ;
        RECT  5.640 4.260 6.040 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.160 4.480 1.740 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.830 4.000 4.770 4.240 ;
        RECT  5.710 2.300 5.950 4.020 ;
        RECT  4.530 3.780 5.950 4.020 ;
        RECT  0.830 3.040 1.070 4.240 ;
        RECT  0.830 3.040 3.410 3.280 ;
        RECT  3.170 0.800 3.410 3.280 ;
        RECT  3.170 2.060 3.530 2.460 ;
        RECT  0.160 0.800 0.560 1.130 ;
        RECT  0.160 0.800 3.410 1.040 ;
        RECT  2.130 3.520 4.260 3.760 ;
        RECT  4.020 1.470 4.260 3.760 ;
        RECT  4.020 2.380 4.590 2.620 ;
        RECT  3.650 1.470 4.260 1.710 ;
        RECT  3.650 1.310 3.890 1.710 ;
    END
END AN4

MACRO AN4B1
    CLASS CORE ;
    FOREIGN AN4B1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.830 2.930 4.170 3.330 ;
        RECT  3.890 1.280 4.650 1.560 ;
        RECT  3.890 1.280 4.170 3.330 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.350 1.760 1.690 2.160 ;
        RECT  1.410 1.180 1.690 2.160 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 2.940 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.100 1.590 3.550 1.990 ;
        RECT  3.270 0.800 5.410 1.040 ;
        RECT  4.870 2.300 5.410 2.700 ;
        RECT  5.130 0.800 5.410 2.740 ;
        RECT  3.270 0.800 3.550 1.990 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.300 0.490 2.700 ;
        RECT  0.170 2.300 0.450 2.940 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.440 -0.380 3.840 0.560 ;
        RECT  5.020 -0.380 5.420 0.560 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.160 -0.380 0.560 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.190 4.480 2.590 5.420 ;
        RECT  5.020 4.260 5.420 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.830 4.480 1.230 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.690 2.800 3.930 ;
        RECT  2.560 1.220 2.800 3.930 ;
        RECT  3.410 2.290 3.650 2.690 ;
        RECT  2.560 2.350 3.650 2.590 ;
    END
END AN4B1

MACRO AN4B1P
    CLASS CORE ;
    FOREIGN AN4B1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.060 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.840 2.940 6.680 3.220 ;
        RECT  3.320 1.260 7.900 1.540 ;
        RECT  4.510 1.260 4.790 3.220 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.540 1.690 2.430 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.400 2.700 ;
        RECT  2.030 2.300 2.310 2.940 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.170 2.380 5.570 2.620 ;
        RECT  5.330 1.790 7.890 2.030 ;
        RECT  7.410 1.790 7.890 2.700 ;
        RECT  7.610 1.790 7.890 2.740 ;
        RECT  5.330 1.790 5.570 2.620 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.300 0.490 2.700 ;
        RECT  0.170 2.300 0.450 2.940 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.830 -0.380 4.230 0.560 ;
        RECT  5.410 -0.380 5.810 0.560 ;
        RECT  6.710 -0.380 7.110 0.560 ;
        RECT  0.000 -0.380 8.060 0.380 ;
        RECT  0.160 -0.380 0.560 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.640 4.260 3.040 5.420 ;
        RECT  5.060 4.260 5.460 5.420 ;
        RECT  7.500 4.260 7.900 5.420 ;
        RECT  0.000 4.660 8.060 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.780 3.080 4.020 ;
        RECT  2.840 0.620 3.080 4.020 ;
        RECT  6.920 2.380 7.160 3.780 ;
        RECT  2.840 3.540 7.160 3.780 ;
        RECT  6.330 2.380 7.160 2.620 ;
        RECT  2.840 2.370 4.010 2.610 ;
        RECT  2.390 0.620 3.080 1.020 ;
    END
END AN4B1P

MACRO AN4B1S
    CLASS CORE ;
    FOREIGN AN4B1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.860 0.640 4.170 1.040 ;
        RECT  2.130 0.800 4.170 1.040 ;
        RECT  3.860 3.220 4.170 3.620 ;
        RECT  3.890 0.640 4.170 3.860 ;
        RECT  2.130 0.720 2.530 1.040 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 0.920 1.690 1.620 ;
        RECT  1.330 0.920 1.690 1.320 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.680 3.050 3.080 ;
        RECT  2.650 2.680 2.930 3.300 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.550 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.990 -0.380 3.390 0.560 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.240 -0.380 0.480 1.190 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.370 4.480 2.770 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.720 4.480 1.120 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.650 3.530 3.890 ;
        RECT  3.290 1.280 3.530 3.890 ;
        RECT  2.450 1.280 2.690 1.860 ;
        RECT  3.290 1.280 3.650 1.680 ;
        RECT  2.450 1.280 3.650 1.520 ;
    END
END AN4B1S

MACRO AN4B1T
    CLASS CORE ;
    FOREIGN AN4B1T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.540 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.860 2.960 4.140 3.340 ;
        RECT  8.870 1.350 9.110 3.200 ;
        RECT  3.860 2.960 9.110 3.200 ;
        RECT  3.850 1.350 10.380 1.590 ;
        RECT  3.860 2.940 4.100 3.340 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.370 2.250 1.690 2.650 ;
        RECT  1.410 1.910 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.250 2.330 2.650 ;
        RECT  2.030 2.160 2.310 2.800 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.250 3.080 2.650 ;
        RECT  2.650 3.580 4.720 3.820 ;
        RECT  4.480 3.540 9.730 3.780 ;
        RECT  9.490 2.250 9.730 3.780 ;
        RECT  9.490 2.250 9.970 2.650 ;
        RECT  2.650 2.160 2.930 3.820 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.100 1.070 2.740 ;
        RECT  0.690 2.250 1.070 2.650 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.570 -0.380 4.970 1.030 ;
        RECT  6.010 -0.380 6.410 1.030 ;
        RECT  7.820 -0.380 8.220 1.030 ;
        RECT  9.260 -0.380 9.660 1.030 ;
        RECT  0.000 -0.380 10.540 0.380 ;
        RECT  0.160 -0.380 0.560 0.800 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.400 4.260 2.800 5.420 ;
        RECT  4.960 4.260 5.360 5.420 ;
        RECT  7.400 4.260 7.800 5.420 ;
        RECT  9.890 4.260 10.290 5.420 ;
        RECT  0.000 4.660 10.540 5.420 ;
        RECT  0.880 3.910 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.430 2.010 3.670 ;
        RECT  0.160 1.150 0.400 3.670 ;
        RECT  8.390 2.280 8.630 2.680 ;
        RECT  3.320 2.330 8.630 2.570 ;
        RECT  3.320 1.150 3.560 2.570 ;
        RECT  3.210 1.150 3.560 1.670 ;
        RECT  0.160 1.150 3.560 1.390 ;
    END
END AN4B1T

MACRO AN4P
    CLASS CORE ;
    FOREIGN AN4P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.490 2.940 4.790 3.340 ;
        RECT  4.110 0.800 4.770 1.040 ;
        RECT  4.530 0.800 4.770 1.540 ;
        RECT  4.510 2.940 4.790 3.860 ;
        RECT  7.610 1.260 7.890 3.220 ;
        RECT  4.490 2.940 7.890 3.220 ;
        RECT  4.530 1.260 8.520 1.540 ;
        RECT  3.800 0.620 4.350 0.860 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.310 2.250 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.880 0.500 2.280 ;
        RECT  0.170 1.540 0.450 2.280 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.990 1.880 2.310 2.280 ;
        RECT  2.030 1.540 2.310 2.280 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.250 2.950 2.650 ;
        RECT  2.650 2.160 2.930 2.800 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.590 -0.380 4.990 0.560 ;
        RECT  6.030 -0.380 6.430 0.560 ;
        RECT  7.330 -0.380 7.730 0.560 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  1.550 -0.380 1.950 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.930 4.480 3.330 5.420 ;
        RECT  5.590 4.260 5.990 5.420 ;
        RECT  8.030 4.260 8.430 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.910 4.160 5.350 4.400 ;
        RECT  5.110 3.540 5.350 4.400 ;
        RECT  1.590 4.000 4.150 4.240 ;
        RECT  1.590 3.040 1.830 4.240 ;
        RECT  5.110 3.540 8.370 3.780 ;
        RECT  8.130 2.300 8.370 3.780 ;
        RECT  0.750 3.040 3.530 3.280 ;
        RECT  3.290 0.800 3.530 3.280 ;
        RECT  3.290 2.030 3.670 2.430 ;
        RECT  0.160 0.800 3.530 1.040 ;
        RECT  2.140 3.520 4.150 3.760 ;
        RECT  3.910 1.340 4.150 3.760 ;
        RECT  3.910 2.380 7.260 2.620 ;
        RECT  3.830 1.340 4.150 1.740 ;
    END
END AN4P

MACRO AN4S
    CLASS CORE ;
    FOREIGN AN4S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.350 3.350 4.790 3.750 ;
        RECT  4.510 0.850 4.790 3.860 ;
        RECT  3.810 0.850 4.790 1.130 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.970 2.360 1.210 2.760 ;
        RECT  0.790 2.100 1.070 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.540 0.500 1.940 ;
        RECT  0.170 1.540 0.450 2.180 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.930 2.860 2.390 3.300 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.630 2.860 3.050 3.300 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.020 -0.380 3.420 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.410 -0.380 1.810 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.950 4.480 3.350 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.160 4.480 1.740 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.130 3.940 4.110 4.180 ;
        RECT  3.870 1.370 4.110 4.180 ;
        RECT  3.870 2.300 4.270 2.700 ;
        RECT  2.500 1.370 4.110 1.610 ;
        RECT  0.750 3.650 1.690 3.890 ;
        RECT  1.450 0.890 1.690 3.890 ;
        RECT  1.450 1.850 3.630 2.090 ;
        RECT  0.160 0.890 1.690 1.130 ;
    END
END AN4S

MACRO AN4T
    CLASS CORE ;
    FOREIGN AN4T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.520 2.960 4.760 3.860 ;
        RECT  9.490 1.350 9.730 3.200 ;
        RECT  4.480 2.960 9.730 3.200 ;
        RECT  4.470 1.350 11.000 1.590 ;
        RECT  4.480 2.940 4.720 3.340 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.310 2.250 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.880 0.500 2.280 ;
        RECT  0.170 1.540 0.450 2.280 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.990 1.880 2.310 2.280 ;
        RECT  2.030 1.540 2.310 2.280 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.250 2.950 2.650 ;
        RECT  2.650 2.160 2.930 2.800 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.190 -0.380 5.590 1.030 ;
        RECT  6.630 -0.380 7.030 1.030 ;
        RECT  8.440 -0.380 8.840 1.030 ;
        RECT  9.880 -0.380 10.280 1.030 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  1.550 -0.380 1.950 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.930 4.480 3.330 5.420 ;
        RECT  5.580 4.260 5.980 5.420 ;
        RECT  8.020 4.260 8.420 5.420 ;
        RECT  10.510 4.260 10.910 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.900 4.160 5.340 4.400 ;
        RECT  5.100 3.540 5.340 4.400 ;
        RECT  1.590 4.000 4.140 4.240 ;
        RECT  1.590 3.040 1.830 4.240 ;
        RECT  5.100 3.540 10.660 3.780 ;
        RECT  10.420 2.250 10.660 3.780 ;
        RECT  0.750 3.040 3.530 3.280 ;
        RECT  3.290 0.800 3.530 3.280 ;
        RECT  10.360 2.250 10.660 2.650 ;
        RECT  3.290 2.030 3.670 2.430 ;
        RECT  0.160 0.800 3.530 1.040 ;
        RECT  2.130 3.520 4.180 3.760 ;
        RECT  3.940 1.270 4.180 3.760 ;
        RECT  9.010 2.280 9.250 2.680 ;
        RECT  3.940 2.330 9.250 2.570 ;
        RECT  3.830 1.270 4.180 1.670 ;
    END
END AN4T

MACRO ANTENNA
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNA 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.240 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.180 1.070 1.620 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.240 0.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 1.240 5.420 ;
        END
    END VCC
END ANTENNA

MACRO AO112
    CLASS CORE ;
    FOREIGN AO112 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.300 0.480 1.700 ;
        RECT  0.170 2.790 0.480 3.190 ;
        RECT  0.170 1.300 0.450 3.190 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.240 3.650 2.640 ;
        RECT  3.270 2.160 3.550 2.740 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.530 4.790 2.180 ;
        RECT  4.470 1.530 4.790 1.930 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.160 1.690 2.810 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.570 2.360 1.970 ;
        RECT  2.030 1.530 2.310 2.180 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.460 -0.380 3.860 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.050 -0.380 1.450 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.450 4.480 2.850 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.740 4.480 1.140 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.910 3.910 4.800 4.150 ;
        RECT  3.910 0.890 4.150 4.150 ;
        RECT  0.700 2.150 1.050 2.550 ;
        RECT  0.810 0.890 1.050 2.550 ;
        RECT  0.810 0.890 4.790 1.130 ;
        RECT  1.530 3.910 3.590 4.150 ;
    END
END AO112

MACRO AO112P
    CLASS CORE ;
    FOREIGN AO112P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.960 1.220 1.200 1.620 ;
        RECT  0.170 1.380 1.200 1.620 ;
        RECT  0.170 2.870 1.280 3.110 ;
        RECT  0.170 1.380 0.450 3.110 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.240 4.280 2.640 ;
        RECT  3.890 1.950 4.170 2.880 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 1.950 5.410 2.880 ;
        RECT  5.090 2.250 5.410 2.650 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.950 2.310 2.890 ;
        RECT  1.950 2.250 2.310 2.650 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.950 2.930 2.890 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  4.230 -0.380 4.630 1.230 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.170 2.000 5.420 ;
        RECT  3.050 3.930 3.450 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.160 4.170 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.530 3.910 5.420 4.150 ;
        RECT  4.530 1.470 4.770 4.150 ;
        RECT  1.190 2.150 1.680 2.550 ;
        RECT  1.440 1.470 1.680 2.550 ;
        RECT  1.440 1.470 5.420 1.710 ;
        RECT  2.330 3.450 4.030 3.690 ;
        RECT  3.640 3.210 4.040 3.450 ;
    END
END AO112P

MACRO AO112S
    CLASS CORE ;
    FOREIGN AO112S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 0.810 0.480 1.210 ;
        RECT  0.170 3.330 0.510 3.730 ;
        RECT  0.170 0.810 0.450 3.730 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.790 3.560 3.190 ;
        RECT  3.270 2.720 3.550 3.370 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.090 4.790 2.740 ;
        RECT  4.410 2.180 4.790 2.580 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.720 1.690 3.370 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.640 2.310 2.290 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.460 -0.380 3.860 0.570 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.040 -0.380 1.440 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.470 4.480 2.870 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.890 4.480 1.290 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.910 3.870 4.800 4.110 ;
        RECT  3.910 0.890 4.150 4.110 ;
        RECT  0.720 1.350 1.050 1.750 ;
        RECT  0.810 0.890 1.050 1.750 ;
        RECT  0.810 0.890 4.800 1.130 ;
        RECT  1.680 3.870 3.590 4.110 ;
    END
END AO112S

MACRO AO112T
    CLASS CORE ;
    FOREIGN AO112T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.220 1.920 1.620 ;
        RECT  0.160 1.380 1.920 1.620 ;
        RECT  0.160 2.870 2.000 3.110 ;
        RECT  0.790 1.380 1.070 3.110 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.240 4.900 2.640 ;
        RECT  4.510 1.940 4.790 2.880 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.950 6.030 2.880 ;
        RECT  5.710 2.250 6.030 2.650 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.950 2.930 2.890 ;
        RECT  2.640 2.250 2.930 2.650 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.250 3.620 2.650 ;
        RECT  3.270 1.950 3.550 2.890 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 2.720 0.950 ;
        RECT  4.850 -0.380 5.250 1.170 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.170 2.720 5.420 ;
        RECT  3.770 3.930 4.170 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.880 4.170 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.150 3.910 6.040 4.150 ;
        RECT  5.150 1.410 5.390 4.150 ;
        RECT  1.910 2.150 2.400 2.550 ;
        RECT  2.160 1.410 2.400 2.550 ;
        RECT  2.160 1.410 6.040 1.650 ;
        RECT  3.050 3.450 4.750 3.690 ;
        RECT  4.340 3.210 4.740 3.690 ;
    END
END AO112T

MACRO AO12
    CLASS CORE ;
    FOREIGN AO12 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 0.620 3.550 3.290 ;
        RECT  3.170 2.890 3.550 3.290 ;
        RECT  3.240 1.260 3.550 1.660 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.510 0.490 1.910 ;
        RECT  0.170 1.090 0.450 1.910 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.890 ;
        RECT  1.310 2.100 1.690 2.500 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.020 2.120 2.310 2.520 ;
        RECT  2.030 1.730 2.310 2.520 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 -0.380 2.640 0.560 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  2.430 4.250 2.830 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.420 1.280 3.760 ;
        RECT  0.880 3.420 2.910 3.660 ;
        RECT  2.670 0.890 2.910 3.660 ;
        RECT  2.670 2.150 3.030 2.550 ;
        RECT  1.440 0.890 2.910 1.130 ;
        RECT  0.160 4.000 2.000 4.240 ;
        RECT  1.600 3.900 2.000 4.240 ;
        RECT  0.160 3.770 0.560 4.240 ;
    END
END AO12

MACRO AO12P
    CLASS CORE ;
    FOREIGN AO12P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.150 3.550 3.260 ;
        RECT  3.170 2.860 3.550 3.260 ;
        RECT  3.140 1.260 3.550 1.660 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.710 0.490 2.110 ;
        RECT  0.170 1.540 0.450 2.180 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.890 ;
        RECT  1.310 2.100 1.690 2.500 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.020 2.120 2.310 2.520 ;
        RECT  2.030 1.730 2.310 2.520 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 -0.380 2.640 0.560 ;
        RECT  3.780 -0.380 4.180 0.930 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 4.180 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  2.430 4.180 2.830 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.400 2.800 3.640 ;
        RECT  2.560 0.890 2.800 3.640 ;
        RECT  2.560 2.150 3.030 2.550 ;
        RECT  1.440 0.890 2.800 1.130 ;
        RECT  0.160 3.880 2.000 4.120 ;
    END
END AO12P

MACRO AO12S
    CLASS CORE ;
    FOREIGN AO12S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 0.810 3.550 3.770 ;
        RECT  3.240 3.370 3.550 3.770 ;
        RECT  3.240 0.810 3.550 1.210 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.350 0.490 1.750 ;
        RECT  0.170 1.060 0.450 1.750 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.970 1.690 2.740 ;
        RECT  1.390 1.970 1.690 2.370 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.730 2.310 2.370 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.370 -0.380 2.770 0.560 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  2.410 4.480 2.810 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.660 1.280 3.900 ;
        RECT  1.040 3.400 1.280 3.900 ;
        RECT  1.040 3.400 2.910 3.640 ;
        RECT  2.670 0.890 2.910 3.640 ;
        RECT  2.670 2.150 2.990 2.550 ;
        RECT  1.440 0.890 2.910 1.130 ;
        RECT  0.240 4.140 2.000 4.380 ;
        RECT  1.600 3.880 2.000 4.380 ;
        RECT  0.240 3.800 0.480 4.380 ;
    END
END AO12S

MACRO AO12T
    CLASS CORE ;
    FOREIGN AO12T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.370 3.550 3.260 ;
        RECT  3.130 2.860 3.550 3.260 ;
        RECT  4.400 1.340 4.800 1.610 ;
        RECT  3.030 1.370 4.800 1.610 ;
        RECT  3.130 2.940 4.800 3.180 ;
        RECT  3.030 1.370 3.550 1.770 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.030 0.490 2.430 ;
        RECT  0.170 1.860 0.450 2.700 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.890 ;
        RECT  1.310 2.100 1.690 2.500 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.910 ;
        RECT  2.020 2.120 2.310 2.520 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.170 -0.380 2.570 1.250 ;
        RECT  3.680 -0.380 4.080 1.130 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.160 -0.380 0.560 1.050 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.790 4.260 4.190 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  2.320 3.880 2.720 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.830 3.400 1.280 3.640 ;
        RECT  0.830 1.490 1.070 3.640 ;
        RECT  2.550 2.030 2.990 2.430 ;
        RECT  2.550 1.490 2.790 2.430 ;
        RECT  0.830 1.490 2.790 1.730 ;
        RECT  0.160 3.880 2.000 4.120 ;
    END
END AO12T

MACRO AO13
    CLASS CORE ;
    FOREIGN AO13 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 3.150 4.790 3.550 ;
        RECT  4.510 1.270 4.790 3.750 ;
        RECT  4.480 1.490 4.790 1.890 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 2.500 0.490 2.900 ;
        RECT  0.160 2.500 0.460 3.300 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.380 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 2.300 2.340 2.880 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.920 3.000 2.320 ;
        RECT  2.650 1.740 2.930 2.320 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.270 -0.380 3.670 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.180 -0.380 0.580 1.130 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.690 3.880 2.090 5.420 ;
        RECT  3.890 4.180 4.290 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.170 3.700 4.150 3.940 ;
        RECT  3.910 0.890 4.150 3.940 ;
        RECT  2.410 0.890 4.150 1.130 ;
        RECT  0.950 3.400 2.850 3.640 ;
    END
END AO13

MACRO AO13P
    CLASS CORE ;
    FOREIGN AO13P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.430 2.910 4.670 3.310 ;
        RECT  4.240 1.570 5.410 1.810 ;
        RECT  5.130 1.570 5.410 3.150 ;
        RECT  4.430 2.910 5.410 3.150 ;
        RECT  4.240 1.410 4.480 1.810 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 2.060 0.490 2.460 ;
        RECT  0.160 2.060 0.460 2.860 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.380 ;
        RECT  1.410 1.740 1.650 2.430 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 1.740 2.340 2.430 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.030 3.010 2.430 ;
        RECT  2.650 1.740 2.930 2.430 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.270 -0.380 3.670 0.950 ;
        RECT  5.020 -0.380 5.420 1.130 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 3.880 2.000 5.420 ;
        RECT  3.710 3.930 4.110 5.420 ;
        RECT  5.020 4.260 5.420 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.160 3.880 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.040 2.870 4.000 3.110 ;
        RECT  3.760 1.190 4.000 3.110 ;
        RECT  3.760 2.250 4.150 2.650 ;
        RECT  2.410 1.190 4.000 1.430 ;
        RECT  2.410 0.970 2.810 1.430 ;
        RECT  0.880 3.400 2.720 3.640 ;
    END
END AO13P

MACRO AO13S
    CLASS CORE ;
    FOREIGN AO13S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 0.970 4.170 4.300 ;
        RECT  3.860 3.900 4.170 4.300 ;
        RECT  3.850 0.970 4.170 1.370 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 1.920 0.490 2.320 ;
        RECT  0.160 1.740 0.460 2.320 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 2.480 1.690 2.880 ;
        RECT  1.410 2.300 1.690 2.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 1.740 2.340 2.320 ;
        RECT  1.970 1.740 2.340 2.140 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.630 2.300 2.950 2.880 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.970 -0.380 3.370 0.560 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.180 -0.380 0.580 1.130 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 4.480 2.060 5.420 ;
        RECT  3.020 4.250 3.420 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.060 3.180 3.530 3.580 ;
        RECT  3.290 0.890 3.530 3.580 ;
        RECT  3.290 2.490 3.650 2.890 ;
        RECT  2.100 0.890 3.530 1.130 ;
        RECT  0.760 3.260 2.540 3.500 ;
    END
END AO13S

MACRO AO13T
    CLASS CORE ;
    FOREIGN AO13T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.410 2.910 4.650 3.310 ;
        RECT  5.130 1.570 5.410 3.150 ;
        RECT  4.280 1.570 6.040 1.810 ;
        RECT  4.410 2.910 6.040 3.150 ;
        RECT  4.280 1.410 4.520 1.810 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 2.030 0.490 2.430 ;
        RECT  0.160 1.740 0.460 2.630 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.630 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 1.740 2.340 2.630 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.030 3.010 2.430 ;
        RECT  2.650 1.740 2.930 2.630 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.270 -0.380 3.670 0.950 ;
        RECT  4.920 -0.380 5.320 1.130 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.670 3.920 4.070 5.420 ;
        RECT  5.000 4.180 5.400 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.040 2.870 4.020 3.110 ;
        RECT  3.780 1.190 4.020 3.110 ;
        RECT  3.780 2.030 4.150 2.430 ;
        RECT  2.410 1.190 4.020 1.430 ;
        RECT  0.880 3.400 2.720 3.640 ;
    END
END AO13T

MACRO AO22
    CLASS CORE ;
    FOREIGN AO22 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.490 0.480 1.890 ;
        RECT  0.170 2.790 0.480 3.190 ;
        RECT  0.170 1.490 0.450 3.190 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.090 4.790 2.710 ;
        RECT  4.420 2.180 4.790 2.580 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.500 3.550 2.150 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.500 1.690 2.150 ;
        RECT  1.390 1.500 1.690 1.900 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 2.950 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.390 -0.380 4.790 0.580 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.050 -0.380 1.450 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.230 4.480 2.630 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.740 4.480 1.140 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.870 3.910 4.790 4.150 ;
        RECT  2.870 3.600 3.110 4.150 ;
        RECT  1.540 3.600 3.110 3.840 ;
        RECT  1.540 3.360 1.940 3.840 ;
        RECT  3.750 3.270 4.150 3.670 ;
        RECT  3.910 0.890 4.150 3.670 ;
        RECT  0.700 2.150 1.050 2.550 ;
        RECT  0.810 0.890 1.050 2.550 ;
        RECT  0.810 0.890 4.150 1.130 ;
    END
END AO22

MACRO AO222
    CLASS CORE ;
    FOREIGN AO222 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.420 6.030 3.300 ;
        RECT  5.720 2.900 6.030 3.300 ;
        RECT  5.720 1.490 6.030 1.890 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.040 2.310 2.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.680 3.120 2.080 ;
        RECT  2.650 1.480 2.930 2.180 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.680 4.800 2.080 ;
        RECT  4.510 1.540 4.790 2.180 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.070 4.170 2.740 ;
        RECT  3.730 2.250 4.170 2.650 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.480 1.690 2.180 ;
        RECT  1.300 1.580 1.690 1.980 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.180 0.530 2.580 ;
        RECT  0.170 2.090 0.450 2.740 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.780 -0.380 5.180 0.560 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  1.650 -0.380 2.050 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.040 4.100 5.480 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  3.570 3.860 3.970 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.810 2.910 1.200 3.310 ;
        RECT  0.810 0.890 1.050 3.310 ;
        RECT  5.150 2.180 5.510 2.580 ;
        RECT  5.150 0.890 5.390 2.580 ;
        RECT  0.160 0.890 5.390 1.130 ;
        RECT  2.260 2.980 4.600 3.220 ;
        RECT  0.240 3.870 3.240 4.110 ;
        RECT  0.240 3.000 0.480 4.110 ;
    END
END AO222

MACRO AO222P
    CLASS CORE ;
    FOREIGN AO222P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 1.530 6.650 3.220 ;
        RECT  5.640 2.940 6.650 3.220 ;
        RECT  5.740 1.530 6.650 1.810 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.040 2.310 2.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.620 2.970 2.020 ;
        RECT  2.650 1.480 2.930 2.180 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.480 4.790 2.180 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.070 4.170 2.740 ;
        RECT  3.860 2.250 4.170 2.650 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.480 1.690 2.180 ;
        RECT  1.290 1.610 1.690 2.010 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.180 0.530 2.580 ;
        RECT  0.170 2.090 0.450 2.740 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.820 -0.380 5.220 0.560 ;
        RECT  6.260 -0.380 6.660 0.880 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  1.650 -0.380 2.050 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.990 4.100 5.430 5.420 ;
        RECT  6.220 4.100 6.670 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  3.630 4.140 4.030 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.810 3.430 1.280 3.670 ;
        RECT  0.810 0.890 1.050 3.670 ;
        RECT  5.150 2.180 5.570 2.580 ;
        RECT  5.150 0.890 5.390 2.580 ;
        RECT  0.160 0.890 5.390 1.130 ;
        RECT  3.370 3.580 4.690 3.820 ;
        RECT  3.370 2.980 3.610 3.820 ;
        RECT  2.280 2.980 3.610 3.220 ;
        RECT  1.410 3.910 1.810 4.390 ;
        RECT  0.240 3.910 3.130 4.150 ;
        RECT  2.890 3.600 3.130 4.150 ;
        RECT  0.240 3.510 0.480 4.150 ;
    END
END AO222P

MACRO AO222S
    CLASS CORE ;
    FOREIGN AO222S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 0.810 6.030 3.570 ;
        RECT  5.720 3.170 6.030 3.570 ;
        RECT  5.720 0.810 6.030 1.210 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.240 2.310 2.940 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.480 2.930 2.180 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.240 4.800 2.640 ;
        RECT  4.510 2.100 4.790 2.740 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.510 4.170 2.180 ;
        RECT  3.880 1.510 4.170 1.910 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.480 1.690 2.180 ;
        RECT  1.300 1.580 1.690 1.980 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.180 0.530 2.580 ;
        RECT  0.170 2.090 0.450 2.740 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.820 -0.380 5.220 0.560 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  1.590 -0.380 1.990 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.050 4.480 5.450 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  3.610 3.830 4.010 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.810 3.250 1.280 3.520 ;
        RECT  0.810 0.800 1.050 3.520 ;
        RECT  5.150 1.350 5.480 1.750 ;
        RECT  5.150 0.800 5.390 1.750 ;
        RECT  3.210 0.800 3.610 1.130 ;
        RECT  0.160 0.800 1.050 1.130 ;
        RECT  0.160 0.800 5.390 1.040 ;
        RECT  2.270 3.250 4.650 3.490 ;
        RECT  0.160 3.860 3.290 4.100 ;
        RECT  1.540 3.840 1.940 4.100 ;
    END
END AO222S

MACRO AO222T
    CLASS CORE ;
    FOREIGN AO222T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.580 1.550 7.280 1.830 ;
        RECT  5.640 2.940 7.280 3.220 ;
        RECT  6.370 1.550 6.650 3.220 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.040 2.310 2.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.910 2.970 2.310 ;
        RECT  2.650 1.480 2.930 2.310 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.470 1.910 4.790 2.310 ;
        RECT  4.510 1.480 4.790 2.310 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.070 4.170 2.740 ;
        RECT  3.790 2.250 4.170 2.650 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.290 1.910 1.690 2.310 ;
        RECT  1.410 1.480 1.690 2.310 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.180 0.530 2.580 ;
        RECT  0.170 2.090 0.450 2.740 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.820 -0.380 5.220 0.560 ;
        RECT  6.290 -0.380 6.690 1.000 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  1.650 -0.380 2.050 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.990 4.100 5.430 5.420 ;
        RECT  6.220 4.100 6.670 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  3.630 4.140 4.030 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.810 3.430 1.280 3.670 ;
        RECT  0.810 0.890 1.050 3.670 ;
        RECT  5.100 2.180 5.570 2.580 ;
        RECT  5.100 0.890 5.340 2.580 ;
        RECT  0.160 0.890 5.340 1.130 ;
        RECT  3.370 3.460 4.660 3.700 ;
        RECT  3.370 2.980 3.610 3.700 ;
        RECT  2.280 2.980 3.610 3.220 ;
        RECT  1.410 3.910 1.810 4.390 ;
        RECT  0.240 3.910 3.130 4.150 ;
        RECT  2.890 3.610 3.130 4.150 ;
        RECT  0.240 3.510 0.480 4.150 ;
    END
END AO222T

MACRO AO22P
    CLASS CORE ;
    FOREIGN AO22P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.390 1.270 1.790 ;
        RECT  0.790 1.190 1.070 3.190 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.090 1.810 5.410 2.210 ;
        RECT  5.130 1.530 5.410 2.210 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.240 4.280 2.640 ;
        RECT  3.890 2.160 4.170 2.780 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.810 2.320 2.210 ;
        RECT  2.030 1.590 2.310 2.210 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.250 3.040 2.650 ;
        RECT  2.650 2.160 2.930 2.780 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.740 -0.380 2.140 0.580 ;
        RECT  5.020 -0.380 5.420 0.580 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.160 -0.380 0.560 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.150 4.100 0.600 5.420 ;
        RECT  1.530 4.130 1.930 5.420 ;
        RECT  3.240 4.100 3.640 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.250 4.090 0.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.870 3.540 5.390 3.780 ;
        RECT  5.090 3.000 5.390 3.780 ;
        RECT  2.230 3.380 4.110 3.620 ;
        RECT  4.380 2.900 4.770 3.300 ;
        RECT  4.530 0.820 4.770 3.300 ;
        RECT  1.310 2.030 1.750 2.430 ;
        RECT  1.510 0.820 1.750 2.430 ;
        RECT  3.210 0.820 3.610 1.130 ;
        RECT  1.510 0.820 4.770 1.060 ;
    END
END AO22P

MACRO AO22S
    CLASS CORE ;
    FOREIGN AO22S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 0.810 0.480 1.210 ;
        RECT  0.170 3.180 0.480 3.580 ;
        RECT  0.170 0.810 0.450 3.580 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.540 4.790 2.180 ;
        RECT  4.470 1.540 4.790 1.940 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.300 3.550 2.940 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.640 1.690 3.370 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.540 2.310 2.180 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.390 -0.380 4.790 0.580 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.950 -0.380 1.350 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.230 4.480 2.630 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.790 4.480 1.190 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.110 3.930 4.790 4.170 ;
        RECT  4.390 3.910 4.790 4.170 ;
        RECT  2.950 3.930 4.790 4.150 ;
        RECT  1.580 3.720 3.350 3.960 ;
        RECT  3.670 3.450 4.150 3.690 ;
        RECT  3.910 0.950 4.150 3.690 ;
        RECT  0.720 1.410 1.050 1.810 ;
        RECT  0.810 0.950 1.050 1.810 ;
        RECT  0.810 0.950 4.150 1.190 ;
    END
END AO22S

MACRO AO22T
    CLASS CORE ;
    FOREIGN AO22T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 2.870 1.900 3.110 ;
        RECT  1.690 1.310 1.930 1.710 ;
        RECT  0.160 1.470 1.930 1.710 ;
        RECT  0.790 1.470 1.070 3.110 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 2.240 6.030 2.640 ;
        RECT  5.750 1.910 6.030 2.640 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.240 4.900 2.640 ;
        RECT  4.510 2.160 4.790 2.780 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.250 2.980 2.650 ;
        RECT  2.650 2.030 2.930 2.650 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.250 3.700 2.650 ;
        RECT  3.270 2.160 3.550 2.780 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.400 -0.380 2.800 0.580 ;
        RECT  5.640 -0.380 6.040 0.950 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.880 -0.380 1.280 1.130 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.190 4.130 2.590 5.420 ;
        RECT  3.850 4.100 4.250 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.760 4.090 1.210 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.490 3.540 6.010 3.780 ;
        RECT  5.710 3.000 6.010 3.780 ;
        RECT  2.890 3.380 4.730 3.620 ;
        RECT  5.000 2.900 5.390 3.300 ;
        RECT  5.150 0.820 5.390 3.300 ;
        RECT  1.970 2.030 2.410 2.430 ;
        RECT  2.170 0.820 2.410 2.430 ;
        RECT  3.870 0.820 4.270 1.130 ;
        RECT  2.170 0.820 5.390 1.060 ;
    END
END AO22T

MACRO AOI112H
    CLASS CORE ;
    FOREIGN AOI112H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.540 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.490 8.510 3.450 ;
        RECT  5.360 1.490 9.660 1.730 ;
        RECT  8.230 3.170 10.380 3.450 ;
        RECT  3.040 1.570 5.600 1.810 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 2.150 7.270 2.790 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 2.150 9.750 2.790 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.150 1.690 2.790 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.150 3.560 2.550 ;
        RECT  3.270 2.150 3.550 2.790 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  5.200 -0.380 5.600 1.010 ;
        RECT  7.100 -0.380 7.500 1.250 ;
        RECT  8.540 -0.380 8.940 1.250 ;
        RECT  9.980 -0.380 10.380 1.250 ;
        RECT  0.000 -0.380 10.540 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.090 5.380 5.420 ;
        RECT  0.000 4.660 10.540 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.380 3.690 9.660 3.930 ;
        RECT  0.880 3.780 4.160 4.020 ;
        RECT  3.920 3.210 4.160 4.020 ;
        RECT  3.920 3.210 7.500 3.450 ;
        RECT  0.880 1.190 2.720 1.430 ;
        RECT  2.480 1.090 4.160 1.330 ;
    END
END AOI112H

MACRO AOI112HP
    CLASS CORE ;
    FOREIGN AOI112HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.220 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.050 1.490 15.330 3.450 ;
        RECT  9.680 1.490 18.330 1.730 ;
        RECT  15.050 3.170 18.330 3.450 ;
        RECT  5.200 1.570 9.920 1.810 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.150 12.230 2.790 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 2.150 16.570 2.790 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.310 2.790 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.650 2.790 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 2.720 0.950 ;
        RECT  3.760 -0.380 4.160 0.950 ;
        RECT  9.520 -0.380 9.920 1.250 ;
        RECT  11.450 -0.380 11.850 1.250 ;
        RECT  12.890 -0.380 13.290 1.250 ;
        RECT  14.330 -0.380 14.730 1.250 ;
        RECT  15.770 -0.380 16.170 1.250 ;
        RECT  17.210 -0.380 17.610 1.250 ;
        RECT  18.650 -0.380 19.050 1.250 ;
        RECT  0.000 -0.380 19.220 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  5.920 4.260 6.320 5.420 ;
        RECT  7.360 4.260 7.760 5.420 ;
        RECT  9.000 4.090 9.400 5.420 ;
        RECT  0.000 4.660 19.220 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.010 3.690 19.050 3.930 ;
        RECT  0.880 3.780 8.480 4.020 ;
        RECT  8.240 3.210 8.480 4.020 ;
        RECT  8.240 3.210 14.010 3.450 ;
        RECT  0.160 1.190 4.880 1.430 ;
        RECT  4.480 1.090 9.200 1.330 ;
    END
END AOI112HP

MACRO AOI112HS
    CLASS CORE ;
    FOREIGN AOI112HS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.490 6.030 3.450 ;
        RECT  3.920 1.490 6.560 1.730 ;
        RECT  5.750 3.170 6.560 3.450 ;
        RECT  2.320 1.570 4.160 1.810 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.810 2.550 ;
        RECT  4.510 2.150 4.790 2.790 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.650 2.790 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.150 1.070 2.800 ;
        RECT  0.730 2.150 1.070 2.550 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.410 2.550 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.760 -0.380 4.160 1.250 ;
        RECT  5.440 -0.380 5.840 1.250 ;
        RECT  6.880 -0.380 7.280 1.250 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.090 3.440 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.000 3.690 7.280 3.930 ;
        RECT  0.880 3.780 2.720 4.020 ;
        RECT  2.480 3.210 2.720 4.020 ;
        RECT  2.480 3.210 5.120 3.450 ;
        RECT  0.160 1.190 2.000 1.430 ;
        RECT  1.600 1.090 3.440 1.330 ;
    END
END AOI112HS

MACRO AOI112HT
    CLASS CORE ;
    FOREIGN AOI112HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.900 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  21.250 1.570 21.530 3.450 ;
        RECT  13.280 1.570 27.020 1.810 ;
        RECT  21.250 3.170 27.740 3.450 ;
        RECT  7.360 1.390 13.520 1.630 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  18.150 2.150 18.430 2.890 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  24.350 2.150 24.630 2.890 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.250 3.550 2.890 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.250 10.370 2.890 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  5.920 -0.380 6.320 0.950 ;
        RECT  13.840 -0.380 14.780 1.250 ;
        RECT  15.820 -0.380 16.220 1.250 ;
        RECT  17.260 -0.380 17.660 1.250 ;
        RECT  18.700 -0.380 19.100 1.250 ;
        RECT  20.140 -0.380 20.540 1.250 ;
        RECT  21.580 -0.380 21.980 1.250 ;
        RECT  23.020 -0.380 23.420 1.250 ;
        RECT  24.460 -0.380 24.860 1.250 ;
        RECT  25.900 -0.380 26.300 1.250 ;
        RECT  27.340 -0.380 27.740 1.250 ;
        RECT  0.000 -0.380 27.900 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  5.920 4.260 6.320 5.420 ;
        RECT  7.360 4.260 7.760 5.420 ;
        RECT  8.800 4.260 9.200 5.420 ;
        RECT  10.240 4.260 10.640 5.420 ;
        RECT  11.680 4.260 12.080 5.420 ;
        RECT  13.120 4.090 14.020 5.420 ;
        RECT  0.000 4.660 27.900 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  15.100 3.690 27.020 3.930 ;
        RECT  0.880 3.510 12.800 3.750 ;
        RECT  12.560 3.210 12.800 3.750 ;
        RECT  12.560 3.210 20.540 3.450 ;
        RECT  0.880 1.190 6.960 1.430 ;
        RECT  6.720 0.900 6.960 1.430 ;
        RECT  6.720 0.900 12.800 1.140 ;
    END
END AOI112HT

MACRO AOI12H
    CLASS CORE ;
    FOREIGN AOI12H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.280 6.030 3.930 ;
        RECT  3.760 3.690 6.030 3.930 ;
        RECT  2.320 1.280 6.030 1.520 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.150 1.070 2.800 ;
        RECT  0.730 2.150 1.070 2.550 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.410 2.550 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.810 2.550 ;
        RECT  4.510 2.150 4.790 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 -0.380 4.180 0.910 ;
        RECT  5.640 -0.380 6.040 0.910 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.090 3.440 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.780 2.720 4.020 ;
        RECT  2.480 3.210 2.720 4.020 ;
        RECT  2.480 3.210 5.120 3.450 ;
        RECT  0.160 1.190 1.920 1.430 ;
        RECT  1.680 0.720 1.920 1.430 ;
        RECT  1.680 0.720 3.440 0.960 ;
    END
END AOI12H

MACRO AOI12HP
    CLASS CORE ;
    FOREIGN AOI12HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.540 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.760 1.280 10.370 1.520 ;
        RECT  10.090 1.280 10.370 4.320 ;
        RECT  6.640 4.080 10.370 4.320 ;
        RECT  6.640 3.690 7.040 4.320 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.150 1.690 2.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.790 2.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.150 8.510 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 2.720 0.950 ;
        RECT  6.660 -0.380 7.060 0.880 ;
        RECT  8.400 -0.380 8.800 0.560 ;
        RECT  9.980 -0.380 10.380 0.560 ;
        RECT  0.000 -0.380 10.540 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  5.920 4.090 6.320 5.420 ;
        RECT  0.000 4.660 10.540 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.780 5.670 4.020 ;
        RECT  5.430 3.210 5.670 4.020 ;
        RECT  7.280 3.520 9.630 3.760 ;
        RECT  7.280 3.210 7.520 3.760 ;
        RECT  5.430 3.210 7.520 3.450 ;
        RECT  0.160 1.190 3.200 1.430 ;
        RECT  2.960 0.720 3.200 1.430 ;
        RECT  2.960 0.720 6.320 0.960 ;
    END
END AOI12HP

MACRO AOI12HS
    CLASS CORE ;
    FOREIGN AOI12HS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.260 4.170 3.310 ;
        RECT  3.830 2.910 4.170 3.310 ;
        RECT  1.600 1.260 4.170 1.540 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.240 0.540 2.640 ;
        RECT  0.170 2.080 0.450 2.750 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.110 1.690 2.750 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.100 3.550 2.740 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.890 -0.380 3.290 0.950 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.790 4.140 2.190 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.160 4.230 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.620 3.300 3.860 ;
    END
END AOI12HS

MACRO AOI12HT
    CLASS CORE ;
    FOREIGN AOI12HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.200 1.280 10.860 1.520 ;
        RECT  10.420 1.340 12.350 1.580 ;
        RECT  11.910 1.280 14.710 1.520 ;
        RECT  14.430 1.280 14.710 4.320 ;
        RECT  9.520 4.080 14.710 4.320 ;
        RECT  9.520 3.690 9.920 4.320 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 2.150 7.270 2.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.150 12.230 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 2.720 0.950 ;
        RECT  3.760 -0.380 4.160 0.950 ;
        RECT  9.540 -0.380 9.940 0.880 ;
        RECT  11.210 -0.380 11.610 1.100 ;
        RECT  12.740 -0.380 13.140 0.560 ;
        RECT  14.320 -0.380 14.720 0.560 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  5.920 4.260 6.320 5.420 ;
        RECT  7.360 4.260 7.760 5.420 ;
        RECT  8.800 4.090 9.200 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.780 8.550 4.020 ;
        RECT  8.310 3.210 8.550 4.020 ;
        RECT  10.160 3.520 13.980 3.760 ;
        RECT  10.160 3.210 10.400 3.760 ;
        RECT  8.310 3.210 10.400 3.450 ;
        RECT  0.160 1.190 4.670 1.430 ;
        RECT  4.430 0.720 4.670 1.430 ;
        RECT  4.430 0.720 9.200 0.960 ;
    END
END AOI12HT

MACRO AOI13H
    CLASS CORE ;
    FOREIGN AOI13H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.520 0.710 5.760 1.730 ;
        RECT  5.770 1.490 6.010 3.490 ;
        RECT  5.770 3.250 6.560 3.490 ;
        RECT  5.520 1.490 7.280 1.730 ;
        RECT  3.860 0.710 5.760 0.950 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.780 2.060 1.110 2.460 ;
        RECT  0.780 2.060 1.080 2.860 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.040 2.930 2.810 ;
        RECT  2.630 2.060 2.930 2.460 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 2.040 4.820 2.810 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.060 6.710 2.460 ;
        RECT  6.370 2.060 6.650 2.810 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.160 -0.380 6.560 1.250 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.650 4.260 5.050 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.780 7.280 4.020 ;
        RECT  2.320 1.210 5.120 1.450 ;
        RECT  0.160 1.190 1.920 1.430 ;
        RECT  1.680 0.710 1.920 1.430 ;
        RECT  1.680 0.710 3.540 0.950 ;
    END
END AOI13H

MACRO AOI13HP
    CLASS CORE ;
    FOREIGN AOI13HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.660 0.710 9.900 1.780 ;
        RECT  10.110 1.540 10.350 3.490 ;
        RECT  10.110 3.250 12.140 3.490 ;
        RECT  9.660 1.540 12.860 1.780 ;
        RECT  6.700 0.710 9.900 0.950 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 2.060 1.730 2.460 ;
        RECT  1.400 2.060 1.700 2.860 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.040 4.790 2.810 ;
        RECT  4.490 2.060 4.790 2.460 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.200 2.040 8.540 2.810 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.060 11.670 2.460 ;
        RECT  11.330 2.060 11.610 2.810 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 2.720 0.950 ;
        RECT  10.300 -0.380 10.700 1.300 ;
        RECT  11.740 -0.380 12.140 1.300 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  5.920 3.930 6.320 5.420 ;
        RECT  7.420 3.930 7.820 5.420 ;
        RECT  8.860 4.260 9.260 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.140 3.780 12.860 4.020 ;
        RECT  8.140 3.450 8.380 4.020 ;
        RECT  0.880 3.450 8.380 3.690 ;
        RECT  3.760 1.210 9.260 1.450 ;
        RECT  0.160 1.190 3.360 1.430 ;
        RECT  3.120 0.710 3.360 1.430 ;
        RECT  3.120 0.710 6.320 0.950 ;
    END
END AOI13HP

MACRO AOI13HS
    CLASS CORE ;
    FOREIGN AOI13HS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.810 1.010 2.580 1.250 ;
        RECT  0.810 3.250 3.560 3.490 ;
        RECT  0.810 1.010 1.050 3.490 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 2.060 0.490 2.460 ;
        RECT  0.160 2.060 0.460 2.860 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.810 ;
        RECT  1.290 2.060 1.690 2.460 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 1.740 2.340 2.810 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.060 3.010 2.460 ;
        RECT  2.650 1.740 2.930 2.810 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.160 -0.380 3.560 1.250 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.160 3.910 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.780 2.720 4.020 ;
    END
END AOI13HS

MACRO AOI13HT
    CLASS CORE ;
    FOREIGN AOI13HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.600 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.800 0.710 14.040 1.780 ;
        RECT  14.450 1.540 14.690 3.490 ;
        RECT  14.440 3.250 17.720 3.490 ;
        RECT  13.800 1.540 18.440 1.780 ;
        RECT  9.400 0.710 14.040 0.950 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.020 2.060 2.320 2.860 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.060 6.650 2.810 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 2.060 11.640 2.810 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 2.060 16.630 2.460 ;
        RECT  16.290 2.060 16.570 2.810 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 2.720 0.950 ;
        RECT  3.760 -0.380 4.160 1.130 ;
        RECT  14.440 -0.380 14.840 1.300 ;
        RECT  15.880 -0.380 16.280 1.300 ;
        RECT  17.320 -0.380 17.720 1.300 ;
        RECT  0.000 -0.380 18.600 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 3.910 4.880 5.420 ;
        RECT  5.920 4.260 6.320 5.420 ;
        RECT  7.360 4.260 7.760 5.420 ;
        RECT  8.800 4.260 9.200 5.420 ;
        RECT  10.120 4.260 10.520 5.420 ;
        RECT  11.560 4.260 11.960 5.420 ;
        RECT  13.000 3.910 13.400 5.420 ;
        RECT  0.000 4.660 18.600 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.720 3.780 18.440 4.020 ;
        RECT  13.720 3.430 13.960 4.020 ;
        RECT  0.880 3.430 13.960 3.670 ;
        RECT  8.240 1.910 9.840 2.150 ;
        RECT  9.600 1.570 9.840 2.150 ;
        RECT  8.240 1.570 8.480 2.150 ;
        RECT  9.600 1.570 13.400 1.810 ;
        RECT  5.200 1.570 8.480 1.810 ;
        RECT  8.800 1.090 9.200 1.670 ;
        RECT  0.160 1.370 4.800 1.610 ;
        RECT  4.560 1.090 4.800 1.610 ;
        RECT  4.560 1.090 9.200 1.330 ;
    END
END AOI13HT

MACRO AOI222H
    CLASS CORE ;
    FOREIGN AOI222H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.180 1.570 7.420 3.450 ;
        RECT  11.950 1.570 12.230 3.450 ;
        RECT  10.620 1.570 12.460 1.810 ;
        RECT  7.180 3.210 14.620 3.450 ;
        RECT  3.040 1.570 7.420 1.810 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 2.150 9.130 2.790 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.650 2.790 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.150 1.690 2.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.150 3.550 2.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 2.150 14.090 2.790 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.150 11.610 2.790 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 1.100 ;
        RECT  8.460 -0.380 8.860 0.950 ;
        RECT  9.900 -0.380 10.300 1.230 ;
        RECT  13.500 -0.380 13.900 0.950 ;
        RECT  14.940 -0.380 15.340 0.950 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.170 4.880 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.300 3.700 15.340 3.940 ;
        RECT  12.780 1.570 14.620 1.810 ;
        RECT  12.780 1.090 13.020 1.810 ;
        RECT  11.340 1.090 13.020 1.330 ;
        RECT  5.740 4.180 10.300 4.420 ;
        RECT  5.740 3.690 5.980 4.420 ;
        RECT  0.880 3.690 5.980 3.930 ;
        RECT  7.740 1.570 9.580 1.810 ;
        RECT  7.740 1.090 7.980 1.810 ;
        RECT  6.300 1.090 7.980 1.330 ;
        RECT  0.880 1.340 2.720 1.580 ;
        RECT  2.480 1.090 2.720 1.580 ;
        RECT  2.480 1.090 4.160 1.330 ;
    END
END AOI222H

MACRO AOI222HP
    CLASS CORE ;
    FOREIGN AOI222HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 28.520 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.620 1.670 20.280 1.910 ;
        RECT  22.490 1.570 22.770 3.450 ;
        RECT  20.040 1.570 23.320 1.810 ;
        RECT  20.040 3.210 27.640 3.450 ;
        RECT  5.200 1.570 13.860 1.810 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 2.150 16.570 2.790 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.150 12.230 2.790 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.310 2.790 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.650 2.790 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  25.590 2.150 25.870 2.790 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  21.250 2.150 21.530 2.790 ;
        RECT  21.250 2.140 21.490 2.790 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 2.720 0.950 ;
        RECT  3.760 -0.380 4.160 0.950 ;
        RECT  14.900 -0.380 15.300 0.950 ;
        RECT  16.340 -0.380 16.740 0.950 ;
        RECT  17.780 -0.380 18.180 0.950 ;
        RECT  24.360 -0.380 24.760 0.950 ;
        RECT  25.800 -0.380 26.200 0.950 ;
        RECT  27.240 -0.380 27.640 0.950 ;
        RECT  0.000 -0.380 28.520 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  5.920 4.260 6.320 5.420 ;
        RECT  7.360 4.260 7.760 5.420 ;
        RECT  9.000 4.170 9.400 5.420 ;
        RECT  0.000 4.660 28.520 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  23.820 1.190 28.360 1.430 ;
        RECT  19.320 1.090 24.060 1.330 ;
        RECT  19.400 3.700 28.360 3.940 ;
        RECT  19.400 3.030 19.640 3.940 ;
        RECT  10.580 3.030 19.640 3.270 ;
        RECT  14.360 1.190 18.900 1.430 ;
        RECT  9.860 1.090 14.600 1.330 ;
        RECT  0.880 3.690 18.900 3.930 ;
        RECT  0.160 1.190 4.880 1.430 ;
        RECT  4.480 1.090 9.200 1.330 ;
    END
END AOI222HP

MACRO AOI222HS
    CLASS CORE ;
    FOREIGN AOI222HS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.170 1.570 5.410 3.450 ;
        RECT  8.440 1.570 9.130 1.810 ;
        RECT  8.850 1.570 9.130 3.450 ;
        RECT  5.170 3.210 10.280 3.450 ;
        RECT  2.320 1.570 5.410 1.810 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.770 2.550 ;
        RECT  6.370 2.150 6.650 2.790 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.930 2.550 ;
        RECT  4.510 2.150 4.790 2.790 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.150 1.070 2.800 ;
        RECT  0.730 2.150 1.070 2.550 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.410 2.550 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.150 10.370 2.790 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.150 8.530 2.550 ;
        RECT  8.230 2.150 8.510 2.790 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.280 -0.380 6.680 1.100 ;
        RECT  9.880 -0.380 10.280 0.960 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.170 3.440 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.370 1.340 11.000 1.580 ;
        RECT  9.370 1.090 9.610 1.580 ;
        RECT  7.720 1.090 9.610 1.330 ;
        RECT  4.840 3.700 11.000 3.940 ;
        RECT  5.720 1.570 7.400 1.810 ;
        RECT  5.720 1.090 5.960 1.810 ;
        RECT  4.120 1.090 5.960 1.330 ;
        RECT  4.280 4.180 7.400 4.420 ;
        RECT  4.280 3.690 4.520 4.420 ;
        RECT  0.880 3.690 4.520 3.930 ;
        RECT  0.160 1.340 1.840 1.580 ;
        RECT  1.600 1.090 2.000 1.430 ;
        RECT  1.600 1.090 3.440 1.330 ;
    END
END AOI222HS

MACRO AOI22H
    CLASS CORE ;
    FOREIGN AOI22H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 1.570 5.410 3.450 ;
        RECT  4.720 3.210 6.560 3.450 ;
        RECT  2.320 1.570 5.410 1.810 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.650 2.790 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.810 2.550 ;
        RECT  4.510 2.150 4.790 2.790 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.150 1.070 2.800 ;
        RECT  0.730 2.150 1.070 2.550 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.410 2.550 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.160 -0.380 6.560 0.950 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.170 3.440 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.650 1.190 7.280 1.430 ;
        RECT  4.000 1.090 5.890 1.330 ;
        RECT  0.880 3.690 7.280 3.930 ;
        RECT  0.160 1.190 2.000 1.430 ;
        RECT  1.600 1.090 3.440 1.330 ;
    END
END AOI22H

MACRO AOI22HP
    CLASS CORE ;
    FOREIGN AOI22HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.760 1.570 9.250 1.810 ;
        RECT  7.410 3.210 12.130 3.450 ;
        RECT  8.850 1.570 9.130 3.450 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.150 11.610 2.790 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.610 2.150 7.890 2.790 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.150 1.690 2.790 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.790 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 2.720 0.950 ;
        RECT  10.290 -0.380 10.690 0.950 ;
        RECT  11.730 -0.380 12.130 0.950 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  5.940 3.930 6.340 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.750 1.190 12.850 1.430 ;
        RECT  6.690 1.090 9.990 1.330 ;
        RECT  6.630 3.690 12.850 3.930 ;
        RECT  6.630 3.030 6.870 3.930 ;
        RECT  0.880 3.030 6.870 3.270 ;
        RECT  0.160 1.190 3.280 1.430 ;
        RECT  3.040 1.090 6.320 1.330 ;
    END
END AOI22HP

MACRO AOI22HT
    CLASS CORE ;
    FOREIGN AOI22HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.220 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.200 1.570 14.010 1.810 ;
        RECT  10.730 3.210 18.330 3.450 ;
        RECT  13.190 1.570 13.470 3.450 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 2.150 16.570 2.790 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.150 12.230 2.790 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.310 2.790 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.650 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 2.720 0.950 ;
        RECT  3.760 -0.380 4.160 0.950 ;
        RECT  15.050 -0.380 15.450 0.950 ;
        RECT  16.490 -0.380 16.890 0.950 ;
        RECT  17.930 -0.380 18.330 0.950 ;
        RECT  0.000 -0.380 19.220 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  5.920 4.260 6.320 5.420 ;
        RECT  7.360 4.260 7.760 5.420 ;
        RECT  9.000 4.170 9.400 5.420 ;
        RECT  0.000 4.660 19.220 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  14.510 1.190 19.050 1.430 ;
        RECT  10.010 1.090 14.750 1.330 ;
        RECT  0.880 3.780 8.480 4.020 ;
        RECT  8.080 3.690 19.050 3.930 ;
        RECT  0.160 1.190 4.880 1.430 ;
        RECT  4.480 1.090 9.200 1.330 ;
    END
END AOI22HT

MACRO AOI22S
    CLASS CORE ;
    FOREIGN AOI22S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.360 1.170 1.760 ;
        RECT  0.790 2.970 1.730 3.250 ;
        RECT  1.490 2.970 1.730 3.370 ;
        RECT  0.790 1.190 1.070 3.250 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.650 2.310 2.370 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.840 1.690 2.730 ;
        RECT  1.310 2.290 1.690 2.690 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.900 2.970 2.300 ;
        RECT  2.650 1.740 2.930 2.350 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.220 0.550 2.740 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  2.290 -0.380 2.690 0.930 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.910 4.160 3.310 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.160 4.190 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.240 1.170 3.480 1.570 ;
        RECT  1.810 1.170 3.480 1.410 ;
        RECT  1.810 0.710 2.050 1.410 ;
        RECT  0.220 0.710 2.050 0.950 ;
        RECT  0.850 4.080 2.340 4.320 ;
        RECT  0.850 3.490 1.090 4.320 ;
        RECT  0.690 3.490 1.090 3.730 ;
    END
END AOI22S

MACRO BHD1
    CLASS CORE ;
    FOREIGN BHD1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.100 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN H
        DIRECTION INOUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.260 2.930 1.540 ;
        RECT  2.620 1.260 2.930 1.890 ;
        RECT  2.650 1.260 2.930 3.520 ;
        RECT  2.620 3.120 2.930 3.520 ;
        RECT  0.790 1.260 1.070 2.430 ;
        END
    END H
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.100 0.380 ;
        RECT  0.950 -0.380 1.350 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.100 5.420 ;
        RECT  1.110 4.480 1.510 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.240 1.490 0.480 3.520 ;
        RECT  0.240 2.670 2.370 2.910 ;
    END
END BHD1

MACRO BUF1
    CLASS CORE ;
    FOREIGN BUF1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.260 2.310 3.270 ;
        RECT  2.000 2.870 2.310 3.270 ;
        RECT  2.000 1.260 2.310 1.660 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.070 2.840 ;
        RECT  0.740 2.240 1.070 2.640 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.200 -0.380 1.600 0.940 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.320 -0.380 0.720 0.910 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  1.180 4.100 1.580 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.190 2.860 0.480 3.260 ;
        RECT  0.190 1.280 0.430 3.260 ;
        RECT  1.420 2.240 1.670 2.640 ;
        RECT  1.430 1.280 1.670 2.640 ;
        RECT  0.190 1.280 0.480 1.890 ;
        RECT  0.190 1.280 1.670 1.520 ;
    END
END BUF1

MACRO BUF12CK
    CLASS CORE ;
    FOREIGN BUF12CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.930 0.680 6.330 4.040 ;
        RECT  7.370 0.680 7.770 4.040 ;
        RECT  8.810 0.680 9.210 4.040 ;
        RECT  10.250 0.680 10.650 4.040 ;
        RECT  4.510 1.680 12.090 3.360 ;
        RECT  11.690 0.680 12.090 4.040 ;
        RECT  4.510 0.680 4.870 4.040 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.850 2.310 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.770 -0.380 4.170 0.780 ;
        RECT  5.210 -0.380 5.610 0.860 ;
        RECT  6.650 -0.380 7.050 0.860 ;
        RECT  8.090 -0.380 8.490 0.860 ;
        RECT  9.530 -0.380 9.930 0.860 ;
        RECT  10.970 -0.380 11.370 0.860 ;
        RECT  0.000 -0.380 12.400 0.380 ;
        RECT  2.320 -0.380 2.720 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.260 2.720 5.420 ;
        RECT  3.770 4.260 4.170 5.420 ;
        RECT  5.210 4.260 5.610 5.420 ;
        RECT  6.650 4.260 7.050 5.420 ;
        RECT  8.090 4.260 8.490 5.420 ;
        RECT  9.530 4.260 9.930 5.420 ;
        RECT  10.970 4.260 11.370 5.420 ;
        RECT  0.000 4.660 12.400 5.420 ;
        RECT  0.880 3.910 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.430 4.270 3.670 ;
        RECT  4.030 1.020 4.270 3.670 ;
        RECT  1.600 1.020 4.270 1.260 ;
    END
END BUF12CK

MACRO BUF1CK
    CLASS CORE ;
    FOREIGN BUF1CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 2.710 1.940 3.860 ;
        RECT  1.600 0.700 2.310 0.980 ;
        RECT  2.030 0.700 2.310 2.990 ;
        RECT  1.660 2.710 2.310 2.990 ;
        RECT  1.680 2.710 1.920 4.040 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.070 2.840 ;
        RECT  0.770 2.250 1.070 2.650 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.880 -0.380 1.280 1.140 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.880 3.730 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.240 0.820 0.480 4.010 ;
        RECT  0.240 1.440 1.470 1.680 ;
    END
END BUF1CK

MACRO BUF1S
    CLASS CORE ;
    FOREIGN BUF1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.050 0.670 2.290 4.020 ;
        RECT  2.000 3.620 2.290 4.020 ;
        RECT  2.000 0.670 2.290 1.070 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.480 2.650 ;
        RECT  0.170 2.250 0.450 3.400 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.300 -0.380 0.700 0.910 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.310 3.760 0.750 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.560 1.490 1.800 3.190 ;
    END
END BUF1S

MACRO BUF2
    CLASS CORE ;
    FOREIGN BUF2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.100 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.060 2.310 3.790 ;
        RECT  1.850 3.280 2.310 3.790 ;
        RECT  1.820 1.060 2.310 1.500 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.150 0.530 2.550 ;
        RECT  0.170 2.050 0.450 2.730 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.380 2.940 0.940 ;
        RECT  0.000 -0.380 3.100 0.380 ;
        RECT  1.100 -0.380 1.500 0.930 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 4.100 2.940 5.420 ;
        RECT  0.000 4.660 3.100 5.420 ;
        RECT  1.080 4.100 1.500 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.580 1.050 3.820 ;
        RECT  0.810 1.220 1.050 3.820 ;
        RECT  0.810 2.280 1.540 2.640 ;
        RECT  0.160 1.220 1.050 1.460 ;
    END
END BUF2

MACRO BUF2CK
    CLASS CORE ;
    FOREIGN BUF2CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.100 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 0.970 2.310 4.040 ;
        RECT  1.890 3.000 2.310 4.040 ;
        RECT  1.810 0.970 2.310 1.250 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.070 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.610 -0.380 2.930 0.950 ;
        RECT  0.000 -0.380 3.100 0.380 ;
        RECT  1.090 -0.380 1.490 0.870 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.530 4.260 2.930 5.420 ;
        RECT  0.000 4.660 3.100 5.420 ;
        RECT  1.090 4.260 1.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.300 3.520 1.550 3.760 ;
        RECT  1.310 1.280 1.550 3.760 ;
        RECT  0.380 1.280 1.550 1.520 ;
        RECT  0.380 0.910 0.620 1.520 ;
    END
END BUF2CK

MACRO BUF3
    CLASS CORE ;
    FOREIGN BUF3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.570 2.310 2.100 ;
        RECT  3.170 1.490 3.550 2.100 ;
        RECT  2.030 1.820 3.550 2.100 ;
        RECT  3.180 2.800 3.550 3.220 ;
        RECT  3.270 1.270 3.550 3.220 ;
        RECT  1.430 2.940 3.550 3.220 ;
        RECT  1.810 1.570 2.310 1.810 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.150 0.540 2.550 ;
        RECT  0.170 1.740 0.450 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 -0.380 2.780 1.210 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.700 -0.380 1.100 0.900 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 4.010 2.700 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.670 4.100 1.070 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.190 3.520 1.050 3.760 ;
        RECT  0.810 1.260 1.050 3.760 ;
        RECT  0.190 3.120 0.480 3.760 ;
        RECT  0.810 2.280 1.550 2.640 ;
        RECT  0.160 1.260 1.050 1.500 ;
    END
END BUF3

MACRO BUF3CK
    CLASS CORE ;
    FOREIGN BUF3CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.350 1.670 4.170 2.250 ;
        RECT  3.770 0.680 4.170 4.040 ;
        RECT  2.350 0.680 2.710 4.040 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.590 1.070 2.280 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.050 -0.380 3.450 0.950 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  1.610 -0.380 2.010 0.870 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.610 4.260 2.010 5.420 ;
        RECT  3.050 4.260 3.450 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.160 3.810 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.860 3.780 2.110 4.020 ;
        RECT  1.870 1.110 2.110 4.020 ;
        RECT  0.960 1.110 2.110 1.350 ;
        RECT  0.960 0.790 1.200 1.350 ;
    END
END BUF3CK

MACRO BUF4
    CLASS CORE ;
    FOREIGN BUF4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.790 3.520 3.200 ;
        RECT  1.410 1.260 3.550 1.820 ;
        RECT  2.640 1.260 2.940 3.200 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.170 0.480 2.570 ;
        RECT  0.170 2.170 0.450 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.270 -0.380 2.690 0.970 ;
        RECT  3.780 -0.380 4.180 0.840 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.670 -0.380 1.070 1.040 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.440 4.100 2.840 5.420 ;
        RECT  3.780 4.100 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.670 4.030 1.070 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.080 1.050 3.440 ;
        RECT  0.810 1.280 1.050 3.440 ;
        RECT  0.810 2.280 2.240 2.520 ;
        RECT  0.160 1.280 1.050 1.760 ;
    END
END BUF4

MACRO BUF4CK
    CLASS CORE ;
    FOREIGN BUF4CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.350 1.670 4.170 2.250 ;
        RECT  3.770 0.680 4.170 4.040 ;
        RECT  2.350 0.680 2.710 4.040 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.590 1.070 2.280 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.050 -0.380 3.450 0.860 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.610 -0.380 2.010 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.610 4.260 2.010 5.420 ;
        RECT  3.050 4.260 3.450 5.420 ;
        RECT  4.400 4.480 4.800 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.160 3.910 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.520 2.110 3.760 ;
        RECT  1.870 1.110 2.110 3.760 ;
        RECT  0.960 1.110 2.110 1.350 ;
        RECT  0.960 0.790 1.200 1.350 ;
    END
END BUF4CK

MACRO BUF6
    CLASS CORE ;
    FOREIGN BUF6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.180 6.660 3.220 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.070 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.550 -0.380 2.950 0.940 ;
        RECT  3.990 -0.380 4.390 0.940 ;
        RECT  5.430 -0.380 5.860 0.940 ;
        RECT  6.880 -0.380 7.280 0.940 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.960 -0.380 1.360 1.340 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.550 4.100 2.950 5.420 ;
        RECT  3.990 4.100 4.390 5.420 ;
        RECT  5.430 4.100 5.830 5.420 ;
        RECT  6.880 4.100 7.280 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.970 4.080 1.370 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.840 2.980 2.290 3.380 ;
        RECT  2.050 1.580 2.290 3.380 ;
        RECT  0.190 2.860 0.480 3.260 ;
        RECT  0.190 1.180 0.430 3.260 ;
        RECT  2.050 2.400 2.910 2.640 ;
        RECT  2.670 2.030 3.030 2.430 ;
        RECT  0.190 1.580 2.290 1.820 ;
        RECT  1.840 1.180 2.110 1.820 ;
        RECT  0.190 1.180 0.480 1.820 ;
    END
END BUF6

MACRO BUF6CK
    CLASS CORE ;
    FOREIGN BUF6CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.490 0.680 4.890 4.040 ;
        RECT  3.070 1.540 6.330 2.380 ;
        RECT  5.930 0.680 6.330 4.040 ;
        RECT  3.070 0.680 3.430 4.040 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.590 1.690 2.280 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.330 -0.380 2.730 0.780 ;
        RECT  3.770 -0.380 4.170 0.860 ;
        RECT  5.210 -0.380 5.610 0.860 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.880 -0.380 1.280 1.110 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.330 4.260 2.730 5.420 ;
        RECT  3.770 4.260 4.170 5.420 ;
        RECT  5.210 4.260 5.610 5.420 ;
        RECT  6.650 4.260 7.050 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.880 3.910 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.430 2.830 3.670 ;
        RECT  2.590 1.110 2.830 3.670 ;
        RECT  1.680 1.110 2.830 1.350 ;
        RECT  1.680 0.790 1.920 1.350 ;
    END
END BUF6CK

MACRO BUF8
    CLASS CORE ;
    FOREIGN BUF8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.060 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.070 1.540 6.970 3.240 ;
        RECT  2.210 2.800 6.970 3.240 ;
        RECT  2.250 1.540 6.970 1.820 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.240 0.530 2.640 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.400 -0.380 1.800 1.020 ;
        RECT  2.970 -0.380 3.370 1.130 ;
        RECT  4.410 -0.380 4.810 1.130 ;
        RECT  5.850 -0.380 6.250 1.130 ;
        RECT  7.500 -0.380 7.900 1.730 ;
        RECT  0.000 -0.380 8.060 0.380 ;
        RECT  0.160 -0.380 0.560 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.490 4.180 1.890 5.420 ;
        RECT  2.910 4.180 3.310 5.420 ;
        RECT  4.340 4.180 4.740 5.420 ;
        RECT  5.850 4.180 6.250 5.420 ;
        RECT  7.500 3.650 7.900 5.420 ;
        RECT  0.000 4.660 8.060 5.420 ;
        RECT  0.160 4.180 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.810 1.490 1.050 3.190 ;
        RECT  0.810 2.160 2.730 2.560 ;
    END
END BUF8

MACRO BUF8CK
    CLASS CORE ;
    FOREIGN BUF8CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.210 0.680 5.610 4.040 ;
        RECT  6.650 0.680 7.050 4.040 ;
        RECT  3.790 1.540 8.490 2.380 ;
        RECT  8.090 0.680 8.490 4.040 ;
        RECT  3.790 0.680 4.150 4.040 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.590 1.690 2.280 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.050 -0.380 3.450 0.780 ;
        RECT  4.490 -0.380 4.890 0.860 ;
        RECT  5.930 -0.380 6.330 0.860 ;
        RECT  7.370 -0.380 7.770 0.860 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  1.600 -0.380 2.000 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.050 4.260 3.450 5.420 ;
        RECT  4.490 4.260 4.890 5.420 ;
        RECT  5.930 4.260 6.330 5.420 ;
        RECT  7.370 4.260 7.770 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.160 3.640 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.520 3.550 3.760 ;
        RECT  3.310 1.110 3.550 3.760 ;
        RECT  2.400 1.110 3.550 1.350 ;
        RECT  2.400 0.790 2.640 1.350 ;
    END
END BUF8CK

MACRO BUFB1
    CLASS CORE ;
    FOREIGN BUFB1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.430 1.020 2.490 1.260 ;
        RECT  1.430 3.300 2.550 3.540 ;
        RECT  1.430 1.020 1.670 3.540 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.600 2.400 3.550 2.640 ;
        RECT  3.270 1.550 3.550 2.830 ;
        RECT  3.270 1.550 4.240 2.010 ;
        RECT  2.600 2.400 3.000 2.650 ;
        END
    END EB
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.480 2.140 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.470 -0.380 3.870 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.880 -0.380 1.280 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.300 4.260 3.700 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.800 4.260 1.200 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.480 1.070 4.720 4.120 ;
        RECT  2.000 1.500 2.240 2.230 ;
        RECT  2.000 1.500 2.970 1.740 ;
        RECT  2.730 1.070 2.970 1.740 ;
        RECT  2.730 1.070 4.720 1.310 ;
        RECT  0.900 3.780 4.030 4.020 ;
        RECT  3.790 2.330 4.030 4.020 ;
        RECT  0.160 3.560 1.140 3.800 ;
        RECT  0.900 1.260 1.140 4.020 ;
        RECT  0.160 1.260 1.140 1.500 ;
    END
END BUFB1

MACRO BUFB2
    CLASS CORE ;
    FOREIGN BUFB2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.070 1.260 5.470 1.570 ;
        RECT  5.070 1.260 6.030 1.540 ;
        RECT  5.750 1.260 6.030 3.220 ;
        RECT  5.210 2.940 6.030 3.220 ;
        RECT  5.210 2.800 5.450 3.220 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.070 2.840 ;
        RECT  0.770 2.230 1.070 2.630 ;
        END
    END EB
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.200 2.930 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.960 -0.380 2.400 0.700 ;
        RECT  4.400 -0.380 4.800 0.970 ;
        RECT  5.640 -0.380 6.040 0.920 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.910 -0.380 1.290 1.500 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.880 3.150 3.120 3.760 ;
        RECT  2.880 3.520 4.150 3.760 ;
        RECT  3.910 3.520 4.150 5.420 ;
        RECT  3.910 4.100 4.720 5.420 ;
        RECT  5.640 4.100 6.040 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.790 4.010 1.190 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.050 3.150 2.400 3.550 ;
        RECT  2.050 1.200 2.290 3.550 ;
        RECT  5.270 1.830 5.510 2.230 ;
        RECT  4.530 1.840 5.510 2.080 ;
        RECT  4.530 1.280 4.770 2.080 ;
        RECT  3.910 1.280 4.770 1.520 ;
        RECT  1.600 1.060 2.050 1.520 ;
        RECT  1.600 1.200 2.910 1.440 ;
        RECT  2.670 0.720 2.910 1.440 ;
        RECT  3.910 0.720 4.150 1.520 ;
        RECT  2.670 0.720 4.150 0.960 ;
        RECT  3.520 3.040 4.150 3.280 ;
        RECT  3.910 1.820 4.150 3.280 ;
        RECT  3.910 2.330 4.910 2.570 ;
        RECT  3.290 1.820 4.150 2.060 ;
        RECT  3.290 1.210 3.530 2.060 ;
        RECT  3.150 1.210 3.530 1.610 ;
        RECT  3.220 4.080 3.620 4.370 ;
        RECT  1.430 4.080 3.620 4.320 ;
        RECT  1.430 3.530 1.670 4.320 ;
        RECT  0.190 3.530 1.670 3.770 ;
        RECT  0.190 1.080 0.430 3.770 ;
        RECT  0.190 2.830 0.480 3.230 ;
        RECT  0.190 1.080 0.480 1.480 ;
    END
END BUFB2

MACRO BUFB3
    CLASS CORE ;
    FOREIGN BUFB3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.440 1.260 6.650 1.540 ;
        RECT  6.280 1.240 6.650 1.640 ;
        RECT  6.370 1.240 6.650 3.220 ;
        RECT  5.020 2.940 6.660 3.220 ;
        RECT  4.440 1.120 4.790 1.540 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.100 1.130 2.720 ;
        END
    END EB
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.200 2.930 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.810 -0.380 1.050 1.840 ;
        RECT  0.810 1.520 1.280 1.840 ;
        RECT  3.840 -0.380 4.260 0.880 ;
        RECT  5.320 -0.380 5.760 1.000 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  0.390 -0.380 1.050 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.720 3.080 2.960 3.760 ;
        RECT  2.720 3.520 3.530 3.760 ;
        RECT  3.290 3.520 3.530 5.420 ;
        RECT  4.180 4.120 4.580 5.420 ;
        RECT  5.720 4.100 6.120 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  0.660 4.020 1.060 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.550 2.980 2.320 3.220 ;
        RECT  1.550 0.720 1.790 3.220 ;
        RECT  5.000 1.840 5.400 2.100 ;
        RECT  3.910 1.840 5.400 2.080 ;
        RECT  1.550 1.440 2.240 1.840 ;
        RECT  3.910 1.140 4.150 2.080 ;
        RECT  3.290 1.140 4.150 1.380 ;
        RECT  3.290 0.720 3.530 1.380 ;
        RECT  1.290 0.720 3.530 0.960 ;
        RECT  1.290 0.620 1.690 0.960 ;
        RECT  3.290 2.400 3.680 3.250 ;
        RECT  3.290 2.400 4.720 2.640 ;
        RECT  4.320 2.320 4.720 2.640 ;
        RECT  3.290 1.720 3.530 3.250 ;
        RECT  2.620 1.720 3.530 1.960 ;
        RECT  2.620 1.240 2.860 1.960 ;
        RECT  2.050 4.130 2.880 4.370 ;
        RECT  2.050 3.540 2.290 4.370 ;
        RECT  0.190 3.540 2.290 3.780 ;
        RECT  0.190 1.490 0.430 3.780 ;
        RECT  0.190 2.800 0.480 3.200 ;
        RECT  0.190 1.490 0.480 1.890 ;
    END
END BUFB3

MACRO BUFT1
    CLASS CORE ;
    FOREIGN BUFT1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.430 1.020 2.490 1.260 ;
        RECT  1.430 3.300 2.550 3.540 ;
        RECT  1.430 1.020 1.670 3.540 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.480 2.140 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.550 2.310 3.060 ;
        RECT  3.290 1.770 3.530 3.060 ;
        RECT  2.030 2.820 3.530 3.060 ;
        RECT  4.000 1.610 4.240 2.010 ;
        RECT  3.290 1.770 4.240 2.010 ;
        RECT  2.000 1.830 2.310 2.230 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.470 -0.380 3.870 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.880 -0.380 1.280 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.300 4.260 3.700 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.800 4.260 1.200 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.480 1.070 4.720 4.120 ;
        RECT  2.600 2.340 3.000 2.580 ;
        RECT  2.760 1.070 3.000 2.580 ;
        RECT  2.760 1.070 4.720 1.310 ;
        RECT  0.900 3.780 4.030 4.020 ;
        RECT  3.790 2.330 4.030 4.020 ;
        RECT  0.160 3.560 1.140 3.800 ;
        RECT  0.900 1.260 1.140 4.020 ;
        RECT  0.160 1.260 1.140 1.500 ;
    END
END BUFT1

MACRO BUFT2
    CLASS CORE ;
    FOREIGN BUFT2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.000 1.160 5.400 1.540 ;
        RECT  5.000 1.260 6.030 1.540 ;
        RECT  5.750 1.260 6.030 3.220 ;
        RECT  5.080 2.940 6.030 3.220 ;
        RECT  5.080 2.940 5.380 3.340 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.200 2.930 2.840 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.070 2.840 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.750 -0.380 3.150 0.810 ;
        RECT  4.390 -0.380 4.750 0.860 ;
        RECT  5.620 -0.380 6.060 0.860 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.750 -0.380 1.190 0.920 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.150 4.080 2.770 5.420 ;
        RECT  4.370 4.100 4.770 5.420 ;
        RECT  5.630 4.100 6.030 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.780 4.100 1.180 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.170 2.860 3.460 3.260 ;
        RECT  3.170 2.960 4.150 3.200 ;
        RECT  3.910 0.620 4.150 3.200 ;
        RECT  5.270 1.780 5.510 2.180 ;
        RECT  3.910 1.840 5.510 2.080 ;
        RECT  3.540 0.620 4.150 0.960 ;
        RECT  1.550 3.540 4.770 3.780 ;
        RECT  4.530 2.320 4.770 3.780 ;
        RECT  1.430 1.820 1.670 3.760 ;
        RECT  1.430 2.990 1.900 3.760 ;
        RECT  4.490 2.320 4.890 2.640 ;
        RECT  1.430 1.820 2.250 2.060 ;
        RECT  2.010 1.530 2.410 1.910 ;
        RECT  0.190 2.980 0.480 3.380 ;
        RECT  0.190 1.260 0.430 3.380 ;
        RECT  3.290 1.720 3.670 2.200 ;
        RECT  0.190 1.260 0.480 1.890 ;
        RECT  3.290 1.260 3.530 2.200 ;
        RECT  2.670 1.260 3.530 1.500 ;
        RECT  0.190 1.260 1.670 1.500 ;
        RECT  1.430 1.050 2.910 1.290 ;
    END
END BUFT2

MACRO BUFT3
    CLASS CORE ;
    FOREIGN BUFT3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.030 2.940 6.660 3.220 ;
        RECT  4.910 1.260 6.650 1.540 ;
        RECT  6.370 1.260 6.650 3.360 ;
        RECT  6.310 2.940 6.660 3.360 ;
        RECT  5.030 2.940 5.370 3.390 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.600 2.200 2.930 2.780 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.070 2.840 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.780 -0.380 3.180 0.810 ;
        RECT  4.300 -0.380 4.660 0.860 ;
        RECT  5.530 -0.380 5.970 0.860 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  0.770 -0.380 1.190 0.990 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 4.040 2.780 5.420 ;
        RECT  4.350 4.160 4.750 5.420 ;
        RECT  5.660 4.160 6.060 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  0.780 4.100 1.200 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.180 2.880 3.420 3.280 ;
        RECT  3.180 2.960 4.150 3.200 ;
        RECT  3.910 1.280 4.150 3.200 ;
        RECT  5.140 1.840 5.540 2.100 ;
        RECT  3.910 1.840 5.540 2.080 ;
        RECT  3.720 0.620 3.960 1.520 ;
        RECT  3.500 0.620 3.960 0.930 ;
        RECT  1.430 3.540 4.770 3.780 ;
        RECT  4.530 2.320 4.770 3.780 ;
        RECT  1.430 1.820 1.670 3.780 ;
        RECT  4.530 2.320 4.790 2.720 ;
        RECT  1.430 1.820 2.270 2.060 ;
        RECT  2.030 1.530 2.430 1.910 ;
        RECT  0.190 2.980 0.480 3.380 ;
        RECT  0.190 1.250 0.430 3.380 ;
        RECT  3.290 1.780 3.670 2.200 ;
        RECT  3.010 1.720 3.530 1.960 ;
        RECT  0.190 1.250 0.480 1.890 ;
        RECT  3.010 1.050 3.250 1.960 ;
        RECT  0.190 1.250 1.670 1.490 ;
        RECT  1.430 1.050 3.250 1.290 ;
    END
END BUFT3

MACRO BUFT4
    CLASS CORE ;
    FOREIGN BUFT4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.020 2.900 5.390 3.300 ;
        RECT  6.370 1.180 6.650 3.220 ;
        RECT  5.020 2.940 6.650 3.220 ;
        RECT  6.270 2.890 6.670 3.130 ;
        RECT  6.290 1.180 6.690 1.540 ;
        RECT  4.910 1.260 6.690 1.540 ;
        RECT  4.910 1.160 5.310 1.540 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.200 2.310 2.840 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.070 2.840 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.780 -0.380 3.180 0.810 ;
        RECT  4.220 -0.380 4.660 0.810 ;
        RECT  5.530 -0.380 5.970 0.840 ;
        RECT  6.880 -0.380 7.280 0.840 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.300 -0.380 0.700 0.900 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.250 4.040 2.650 5.420 ;
        RECT  4.220 4.100 4.620 5.420 ;
        RECT  5.550 4.100 5.950 5.420 ;
        RECT  6.880 4.100 7.280 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.670 4.100 1.090 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.040 2.960 3.440 3.270 ;
        RECT  3.040 2.960 4.150 3.200 ;
        RECT  3.910 1.050 4.150 3.200 ;
        RECT  5.110 1.820 5.510 2.100 ;
        RECT  3.910 1.820 5.510 2.060 ;
        RECT  3.480 0.730 3.920 1.290 ;
        RECT  1.430 3.490 1.860 3.810 ;
        RECT  1.430 3.520 4.770 3.760 ;
        RECT  4.530 2.320 4.770 3.760 ;
        RECT  1.430 1.580 1.670 3.810 ;
        RECT  4.410 2.320 4.810 2.560 ;
        RECT  1.430 1.580 2.430 1.820 ;
        RECT  2.030 1.570 2.430 1.820 ;
        RECT  0.190 2.980 0.480 3.380 ;
        RECT  0.190 1.260 0.430 3.380 ;
        RECT  3.270 1.840 3.670 2.100 ;
        RECT  2.670 1.840 3.670 2.080 ;
        RECT  0.190 1.260 0.480 1.890 ;
        RECT  2.670 1.050 2.910 2.080 ;
        RECT  0.190 1.260 1.190 1.500 ;
        RECT  0.950 1.050 2.910 1.290 ;
    END
END BUFT4

MACRO CMPE4
    CLASS CORE ;
    FOREIGN CMPE4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 29.140 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  28.480 2.300 28.970 2.740 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  23.110 2.300 23.390 2.740 ;
        RECT  22.870 2.330 23.390 2.730 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 2.330 6.250 2.730 ;
        RECT  5.750 2.300 6.030 2.740 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.300 0.590 2.740 ;
        END
    END B0
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  25.930 2.080 26.490 2.480 ;
        RECT  26.210 1.550 26.490 2.480 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  20.630 2.140 20.910 2.870 ;
        RECT  20.390 2.320 20.910 2.720 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.320 8.750 2.720 ;
        RECT  8.230 2.120 8.510 2.850 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.300 3.160 2.740 ;
        END
    END A0
    PIN OEQ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.120 1.580 17.810 1.860 ;
        RECT  17.530 1.580 17.810 4.020 ;
        RECT  15.900 3.740 17.810 4.020 ;
        RECT  15.900 3.740 16.180 4.240 ;
        END
    END OEQ
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.460 -0.380 2.860 0.560 ;
        RECT  5.610 -0.380 6.010 0.560 ;
        RECT  6.620 -0.380 7.020 0.560 ;
        RECT  12.450 -0.380 12.850 0.560 ;
        RECT  22.200 -0.380 22.600 0.560 ;
        RECT  23.080 -0.380 23.480 0.560 ;
        RECT  26.240 -0.380 26.640 0.560 ;
        RECT  28.580 -0.380 28.980 0.560 ;
        RECT  0.000 -0.380 29.140 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 3.950 2.960 5.420 ;
        RECT  5.750 4.480 6.150 5.420 ;
        RECT  8.150 4.200 8.550 5.420 ;
        RECT  11.240 4.480 11.640 5.420 ;
        RECT  12.750 4.480 13.150 5.420 ;
        RECT  14.130 4.480 14.530 5.420 ;
        RECT  17.350 4.260 17.750 5.420 ;
        RECT  20.540 4.200 20.940 5.420 ;
        RECT  22.940 4.480 23.340 5.420 ;
        RECT  26.130 3.950 26.530 5.420 ;
        RECT  28.580 4.480 28.980 5.420 ;
        RECT  0.000 4.660 29.140 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  27.890 2.910 28.170 3.310 ;
        RECT  27.890 0.970 28.130 3.310 ;
        RECT  26.730 0.970 28.130 1.210 ;
        RECT  25.250 0.910 26.970 1.150 ;
        RECT  23.940 3.470 27.450 3.710 ;
        RECT  27.210 2.910 27.450 3.710 ;
        RECT  23.940 1.450 24.180 3.710 ;
        RECT  23.840 2.910 24.180 3.310 ;
        RECT  27.250 1.450 27.490 3.150 ;
        RECT  27.090 1.450 27.490 1.690 ;
        RECT  23.830 1.450 24.230 1.690 ;
        RECT  25.360 2.990 26.970 3.230 ;
        RECT  26.730 2.190 26.970 3.230 ;
        RECT  25.360 1.450 25.600 3.230 ;
        RECT  26.730 2.190 27.010 2.590 ;
        RECT  25.360 1.450 25.950 1.690 ;
        RECT  24.620 2.990 25.020 3.230 ;
        RECT  24.660 0.970 24.900 3.230 ;
        RECT  13.160 0.620 13.400 2.650 ;
        RECT  24.660 1.370 25.010 1.770 ;
        RECT  22.780 0.970 24.900 1.210 ;
        RECT  21.630 0.800 23.020 1.040 ;
        RECT  13.160 0.620 21.870 0.860 ;
        RECT  22.300 3.160 22.600 3.560 ;
        RECT  22.300 1.280 22.540 3.560 ;
        RECT  21.150 1.280 22.540 1.520 ;
        RECT  19.660 1.100 21.390 1.340 ;
        RECT  18.350 3.720 21.880 3.960 ;
        RECT  21.640 3.160 21.880 3.960 ;
        RECT  18.350 1.640 18.590 3.960 ;
        RECT  18.250 3.160 18.590 3.560 ;
        RECT  21.660 1.760 21.900 3.400 ;
        RECT  21.500 1.760 21.900 2.000 ;
        RECT  18.240 1.640 18.640 1.880 ;
        RECT  19.770 3.240 21.390 3.480 ;
        RECT  21.150 2.440 21.390 3.480 ;
        RECT  19.770 1.760 20.010 3.480 ;
        RECT  21.150 2.440 21.420 2.840 ;
        RECT  19.770 1.760 20.360 2.000 ;
        RECT  19.030 3.240 19.430 3.480 ;
        RECT  19.070 1.100 19.310 3.480 ;
        RECT  14.050 1.100 14.290 2.500 ;
        RECT  19.070 1.560 19.420 1.960 ;
        RECT  14.050 1.100 19.310 1.340 ;
        RECT  12.680 3.470 15.250 3.710 ;
        RECT  15.010 2.450 15.250 3.710 ;
        RECT  12.680 1.560 12.920 3.710 ;
        RECT  11.930 2.990 12.920 3.230 ;
        RECT  15.010 2.660 17.220 2.900 ;
        RECT  16.820 2.450 17.220 2.900 ;
        RECT  15.010 2.450 15.410 2.900 ;
        RECT  12.540 1.560 12.920 1.960 ;
        RECT  13.780 2.990 14.770 3.230 ;
        RECT  14.530 1.640 14.770 3.230 ;
        RECT  15.860 2.100 16.260 2.420 ;
        RECT  15.640 1.840 15.880 2.340 ;
        RECT  14.530 1.840 15.880 2.080 ;
        RECT  14.530 1.640 14.930 2.080 ;
        RECT  4.070 2.990 4.470 3.230 ;
        RECT  4.190 0.800 4.430 3.230 ;
        RECT  11.970 2.250 12.440 2.650 ;
        RECT  11.970 0.620 12.210 2.650 ;
        RECT  4.150 1.370 4.430 1.770 ;
        RECT  4.190 0.800 7.510 1.040 ;
        RECT  7.270 0.620 12.210 0.860 ;
        RECT  9.660 3.240 10.060 3.480 ;
        RECT  9.780 1.100 10.020 3.480 ;
        RECT  11.490 1.100 11.730 2.500 ;
        RECT  9.590 1.680 10.020 1.920 ;
        RECT  9.780 1.100 11.730 1.340 ;
        RECT  7.270 3.720 10.740 3.960 ;
        RECT  10.500 1.580 10.740 3.960 ;
        RECT  7.270 3.160 7.510 3.960 ;
        RECT  10.500 3.160 10.840 3.560 ;
        RECT  7.190 1.760 7.430 3.400 ;
        RECT  7.190 1.760 7.590 2.000 ;
        RECT  10.450 1.680 10.850 1.920 ;
        RECT  6.550 1.280 6.790 3.560 ;
        RECT  6.550 1.280 7.990 1.520 ;
        RECT  7.750 1.100 9.430 1.340 ;
        RECT  7.750 3.240 9.320 3.480 ;
        RECT  9.080 1.760 9.320 3.480 ;
        RECT  7.750 2.440 7.990 3.480 ;
        RECT  7.670 2.440 7.990 2.840 ;
        RECT  8.730 1.760 9.320 2.000 ;
        RECT  1.680 3.470 5.150 3.710 ;
        RECT  4.910 1.370 5.150 3.710 ;
        RECT  1.680 2.910 1.920 3.710 ;
        RECT  4.910 2.910 5.250 3.310 ;
        RECT  1.600 1.450 1.840 3.150 ;
        RECT  4.910 1.370 5.250 1.770 ;
        RECT  1.600 1.450 2.000 1.690 ;
        RECT  0.960 0.800 1.200 3.310 ;
        RECT  0.960 0.800 3.840 1.040 ;
        RECT  2.160 2.990 3.730 3.230 ;
        RECT  3.490 1.370 3.730 3.230 ;
        RECT  2.160 2.200 2.400 3.230 ;
        RECT  2.080 2.190 2.320 2.590 ;
        RECT  3.290 1.370 3.730 1.770 ;
    END
END CMPE4

MACRO CMPE4S
    CLASS CORE ;
    FOREIGN CMPE4S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 29.140 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  28.480 2.300 28.970 2.740 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  23.110 2.300 23.390 2.740 ;
        RECT  22.870 2.330 23.390 2.730 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 2.330 6.250 2.730 ;
        RECT  5.750 2.300 6.030 2.740 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.300 0.590 2.740 ;
        END
    END B0
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  25.930 2.300 26.490 2.740 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  20.630 2.060 20.910 2.860 ;
        RECT  20.390 2.320 20.910 2.720 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.320 8.750 2.720 ;
        RECT  8.230 2.050 8.510 2.820 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.300 3.160 2.740 ;
        END
    END A0
    PIN OEQ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.530 1.580 17.810 3.710 ;
        RECT  15.550 3.430 17.810 3.710 ;
        RECT  16.120 1.580 17.810 1.860 ;
        END
    END OEQ
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.460 -0.380 2.860 0.560 ;
        RECT  5.610 -0.380 6.010 0.560 ;
        RECT  6.630 -0.380 7.030 0.560 ;
        RECT  12.450 -0.380 12.850 0.560 ;
        RECT  22.210 -0.380 22.610 0.560 ;
        RECT  23.080 -0.380 23.480 0.560 ;
        RECT  26.230 -0.380 26.630 0.560 ;
        RECT  28.580 -0.380 28.980 0.560 ;
        RECT  0.000 -0.380 29.140 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 4.200 2.960 5.420 ;
        RECT  5.750 4.480 6.150 5.420 ;
        RECT  8.150 4.200 8.550 5.420 ;
        RECT  11.240 4.480 11.640 5.420 ;
        RECT  12.750 4.480 13.150 5.420 ;
        RECT  14.130 4.480 14.530 5.420 ;
        RECT  17.350 3.950 17.750 5.420 ;
        RECT  20.540 4.200 20.940 5.420 ;
        RECT  22.940 4.480 23.340 5.420 ;
        RECT  26.130 4.200 26.530 5.420 ;
        RECT  28.580 4.480 28.980 5.420 ;
        RECT  0.000 4.660 29.140 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  27.970 0.800 28.210 3.310 ;
        RECT  25.250 0.800 28.210 1.040 ;
        RECT  25.250 0.740 25.650 1.040 ;
        RECT  23.840 4.080 25.890 4.320 ;
        RECT  25.650 3.720 25.890 4.320 ;
        RECT  23.840 1.280 24.080 4.320 ;
        RECT  25.650 3.720 27.490 3.960 ;
        RECT  27.250 1.280 27.490 3.960 ;
        RECT  25.480 3.230 27.010 3.470 ;
        RECT  26.770 1.280 27.010 3.470 ;
        RECT  25.550 1.280 27.010 1.520 ;
        RECT  24.380 3.230 25.020 3.470 ;
        RECT  24.380 0.800 24.620 3.470 ;
        RECT  13.160 0.620 13.400 2.650 ;
        RECT  24.380 1.280 25.020 1.520 ;
        RECT  21.630 0.800 24.620 1.040 ;
        RECT  13.160 0.620 21.870 0.860 ;
        RECT  22.300 3.160 22.600 3.560 ;
        RECT  22.300 1.280 22.540 3.560 ;
        RECT  21.150 1.280 22.540 1.520 ;
        RECT  19.660 1.100 21.390 1.340 ;
        RECT  18.350 3.720 21.880 3.960 ;
        RECT  21.640 3.160 21.880 3.960 ;
        RECT  18.350 1.580 18.590 3.960 ;
        RECT  18.250 3.160 18.590 3.560 ;
        RECT  21.660 1.760 21.900 3.400 ;
        RECT  21.500 1.760 21.900 2.000 ;
        RECT  18.240 1.580 18.640 1.820 ;
        RECT  19.770 3.240 21.390 3.480 ;
        RECT  21.150 2.440 21.390 3.480 ;
        RECT  19.770 1.760 20.010 3.480 ;
        RECT  21.150 2.440 21.420 2.840 ;
        RECT  19.770 1.760 20.360 2.000 ;
        RECT  19.030 3.240 19.430 3.480 ;
        RECT  19.070 1.100 19.310 3.480 ;
        RECT  14.050 1.100 14.290 2.500 ;
        RECT  19.070 1.500 19.420 1.900 ;
        RECT  14.050 1.100 19.310 1.340 ;
        RECT  12.680 3.470 15.310 3.710 ;
        RECT  15.070 2.660 15.310 3.710 ;
        RECT  12.680 1.560 12.920 3.710 ;
        RECT  11.930 2.990 12.920 3.230 ;
        RECT  15.070 2.660 17.220 2.900 ;
        RECT  16.820 2.450 17.220 2.900 ;
        RECT  12.540 1.560 12.920 1.960 ;
        RECT  13.780 2.990 14.770 3.230 ;
        RECT  14.530 1.640 14.770 3.230 ;
        RECT  15.870 2.100 16.270 2.420 ;
        RECT  15.640 1.840 15.880 2.340 ;
        RECT  14.530 1.840 15.880 2.080 ;
        RECT  14.530 1.640 14.930 2.080 ;
        RECT  4.150 0.800 4.390 3.570 ;
        RECT  11.970 2.250 12.440 2.650 ;
        RECT  11.970 0.620 12.210 2.650 ;
        RECT  4.150 0.800 7.510 1.040 ;
        RECT  7.270 0.620 12.210 0.860 ;
        RECT  9.660 3.240 10.060 3.480 ;
        RECT  9.780 1.100 10.020 3.480 ;
        RECT  11.490 1.100 11.730 2.500 ;
        RECT  9.590 1.580 10.020 1.820 ;
        RECT  9.780 1.100 11.730 1.340 ;
        RECT  7.270 3.720 10.740 3.960 ;
        RECT  10.500 1.580 10.740 3.960 ;
        RECT  7.270 3.160 7.510 3.960 ;
        RECT  10.500 3.160 10.840 3.560 ;
        RECT  7.190 1.760 7.430 3.400 ;
        RECT  7.190 1.760 7.590 2.000 ;
        RECT  10.450 1.580 10.850 1.820 ;
        RECT  6.550 1.280 6.790 3.560 ;
        RECT  6.550 1.280 7.990 1.520 ;
        RECT  7.750 1.100 9.430 1.340 ;
        RECT  7.750 3.240 9.320 3.480 ;
        RECT  9.080 1.680 9.320 3.480 ;
        RECT  7.750 2.440 7.990 3.480 ;
        RECT  7.670 2.440 7.990 2.840 ;
        RECT  8.810 1.680 9.320 2.080 ;
        RECT  3.290 4.180 5.250 4.420 ;
        RECT  5.010 1.370 5.250 4.420 ;
        RECT  3.290 3.720 3.530 4.420 ;
        RECT  1.600 3.720 3.530 3.960 ;
        RECT  1.600 1.450 1.840 3.960 ;
        RECT  1.600 1.450 2.000 1.690 ;
        RECT  0.880 2.910 1.200 3.310 ;
        RECT  0.960 0.800 1.200 3.310 ;
        RECT  0.960 0.800 3.910 1.040 ;
        RECT  2.080 3.240 3.730 3.480 ;
        RECT  3.490 1.370 3.730 3.480 ;
        RECT  2.080 2.620 2.320 3.480 ;
        RECT  3.290 1.370 3.730 1.770 ;
    END
END CMPE4S

MACRO DBFRBN
    CLASS CORE ;
    FOREIGN DBFRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.140 8.610 2.540 ;
        RECT  8.230 1.930 8.510 2.650 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 1.300 12.850 3.840 ;
        RECT  12.510 3.440 12.850 3.840 ;
        RECT  12.510 1.300 12.850 1.700 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  2.010 2.230 2.310 2.630 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.140 1.080 2.540 ;
        RECT  0.790 2.120 1.070 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 1.300 11.610 3.400 ;
        RECT  11.280 3.000 11.610 3.400 ;
        RECT  11.280 1.300 11.610 1.700 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  8.250 -0.380 8.650 0.560 ;
        RECT  10.480 -0.380 10.880 0.860 ;
        RECT  11.710 -0.380 12.110 0.860 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  1.100 -0.380 2.790 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.500 4.020 2.900 5.420 ;
        RECT  8.080 4.480 8.480 5.420 ;
        RECT  10.110 4.130 10.510 5.420 ;
        RECT  11.710 4.260 12.110 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.460 4.180 5.900 4.420 ;
        RECT  5.660 3.580 5.900 4.420 ;
        RECT  4.460 0.620 4.700 4.420 ;
        RECT  4.380 3.620 4.700 4.020 ;
        RECT  10.720 3.720 12.260 3.960 ;
        RECT  12.020 2.140 12.260 3.960 ;
        RECT  5.660 3.580 9.000 3.820 ;
        RECT  8.760 2.880 9.000 3.820 ;
        RECT  10.720 1.100 10.960 3.960 ;
        RECT  8.760 2.880 10.960 3.120 ;
        RECT  9.920 1.100 10.960 1.340 ;
        RECT  9.920 0.620 10.160 1.340 ;
        RECT  9.760 0.620 10.160 0.860 ;
        RECT  4.300 0.620 4.700 0.860 ;
        RECT  10.240 1.640 10.480 2.540 ;
        RECT  9.660 1.640 10.480 1.880 ;
        RECT  9.660 1.580 10.060 1.880 ;
        RECT  9.010 4.090 9.530 4.330 ;
        RECT  9.290 3.420 9.530 4.330 ;
        RECT  9.290 3.420 10.460 3.660 ;
        RECT  4.940 3.700 5.420 3.940 ;
        RECT  4.940 1.100 5.180 3.940 ;
        RECT  8.980 2.120 9.830 2.360 ;
        RECT  8.980 1.120 9.220 2.360 ;
        RECT  6.830 1.120 9.220 1.360 ;
        RECT  4.940 1.100 7.070 1.340 ;
        RECT  5.310 0.860 5.710 1.340 ;
        RECT  7.580 0.620 7.980 0.880 ;
        RECT  6.180 0.620 7.980 0.860 ;
        RECT  7.730 1.600 7.970 3.220 ;
        RECT  6.140 2.880 7.970 3.120 ;
        RECT  6.140 1.600 7.970 1.840 ;
        RECT  6.140 1.580 6.540 1.840 ;
        RECT  6.190 4.160 7.820 4.400 ;
        RECT  5.420 2.880 5.820 3.120 ;
        RECT  5.500 1.580 5.740 3.120 ;
        RECT  5.500 2.220 6.820 2.460 ;
        RECT  5.420 1.580 5.820 1.820 ;
        RECT  3.980 1.290 4.220 3.200 ;
        RECT  0.190 2.800 0.480 3.200 ;
        RECT  0.190 0.800 0.430 3.200 ;
        RECT  3.820 0.800 4.060 1.530 ;
        RECT  0.190 0.800 0.480 1.330 ;
        RECT  0.190 0.800 4.060 1.040 ;
        RECT  3.300 3.940 4.080 4.340 ;
        RECT  3.300 3.430 3.540 4.340 ;
        RECT  3.260 1.500 3.500 3.670 ;
        RECT  3.260 2.040 3.690 2.440 ;
        RECT  1.710 3.540 2.800 3.780 ;
        RECT  2.560 1.580 2.800 3.780 ;
        RECT  2.560 2.260 3.010 2.660 ;
        RECT  1.710 1.580 2.800 1.820 ;
    END
END DBFRBN

MACRO DBFRSBN
    CLASS CORE ;
    FOREIGN DBFRSBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.370 3.210 ;
        RECT  9.700 2.140 10.370 2.540 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 1.300 14.710 3.840 ;
        RECT  14.400 3.440 14.710 3.840 ;
        RECT  14.400 1.300 14.710 1.700 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  2.020 2.230 2.310 2.630 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.300 13.470 3.400 ;
        RECT  13.170 3.000 13.470 3.400 ;
        RECT  13.170 1.300 13.470 1.700 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.100 1.620 9.340 2.450 ;
        RECT  7.370 2.210 9.340 2.450 ;
        RECT  10.100 1.100 10.340 1.860 ;
        RECT  9.100 1.620 10.340 1.860 ;
        RECT  10.100 1.100 11.610 1.340 ;
        RECT  11.330 1.100 11.610 2.210 ;
        RECT  7.370 2.140 7.610 2.540 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.360 -0.380 2.760 0.560 ;
        RECT  8.980 -0.380 9.380 0.560 ;
        RECT  12.370 -0.380 12.770 0.860 ;
        RECT  13.600 -0.380 14.000 0.860 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  1.410 -0.380 1.810 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.500 4.030 2.900 5.420 ;
        RECT  9.410 4.480 9.810 5.420 ;
        RECT  12.130 4.130 12.530 5.420 ;
        RECT  13.600 4.260 14.000 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.460 4.180 5.900 4.420 ;
        RECT  5.660 3.580 5.900 4.420 ;
        RECT  4.460 0.620 4.700 4.420 ;
        RECT  4.380 3.620 4.700 4.020 ;
        RECT  12.690 3.690 14.150 3.930 ;
        RECT  13.910 2.140 14.150 3.930 ;
        RECT  8.430 3.580 10.850 3.820 ;
        RECT  10.610 2.940 10.850 3.820 ;
        RECT  5.660 3.580 7.300 3.820 ;
        RECT  12.690 1.100 12.930 3.930 ;
        RECT  7.060 3.360 8.670 3.600 ;
        RECT  10.610 2.940 12.930 3.180 ;
        RECT  11.890 1.100 12.930 1.340 ;
        RECT  11.890 0.620 12.130 1.340 ;
        RECT  11.090 0.620 12.130 0.860 ;
        RECT  4.300 0.620 4.700 0.860 ;
        RECT  10.730 2.450 12.450 2.690 ;
        RECT  12.210 2.140 12.450 2.690 ;
        RECT  10.730 1.580 10.970 2.690 ;
        RECT  10.580 1.580 10.980 1.820 ;
        RECT  10.340 4.090 11.330 4.330 ;
        RECT  11.090 3.480 11.330 4.330 ;
        RECT  11.090 3.480 12.350 3.720 ;
        RECT  4.940 3.700 5.420 3.940 ;
        RECT  4.940 1.100 5.180 3.940 ;
        RECT  6.830 1.120 9.860 1.360 ;
        RECT  9.620 0.620 9.860 1.360 ;
        RECT  4.940 1.100 7.070 1.340 ;
        RECT  5.310 0.860 5.710 1.340 ;
        RECT  9.620 0.620 10.710 0.860 ;
        RECT  9.060 2.820 9.300 3.220 ;
        RECT  6.140 2.880 9.300 3.120 ;
        RECT  6.890 1.600 7.130 3.120 ;
        RECT  6.140 1.600 8.660 1.840 ;
        RECT  6.140 1.580 6.540 1.840 ;
        RECT  6.190 4.160 9.150 4.400 ;
        RECT  7.670 3.840 8.070 4.400 ;
        RECT  8.340 0.620 8.740 0.880 ;
        RECT  6.180 0.620 8.740 0.860 ;
        RECT  5.420 2.880 5.820 3.120 ;
        RECT  5.500 1.580 5.740 3.120 ;
        RECT  6.410 2.140 6.650 2.540 ;
        RECT  5.500 2.220 6.650 2.460 ;
        RECT  5.420 1.580 5.820 1.820 ;
        RECT  3.980 1.290 4.220 3.200 ;
        RECT  0.960 1.010 1.200 3.190 ;
        RECT  3.840 1.010 4.080 1.530 ;
        RECT  0.160 1.010 4.080 1.250 ;
        RECT  3.230 3.950 4.080 4.350 ;
        RECT  3.230 1.500 3.470 4.350 ;
        RECT  3.230 2.040 3.660 2.440 ;
        RECT  1.710 3.930 2.110 4.170 ;
        RECT  1.870 3.540 2.110 4.170 ;
        RECT  1.870 3.540 2.910 3.780 ;
        RECT  2.670 1.580 2.910 3.780 ;
        RECT  2.670 3.100 2.980 3.500 ;
        RECT  1.710 1.580 2.910 1.820 ;
    END
END DBFRSBN

MACRO DBHRBN
    CLASS CORE ;
    FOREIGN DBHRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.300 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.760 2.930 2.700 ;
        RECT  2.500 2.050 2.930 2.450 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.820 2.790 9.130 3.190 ;
        RECT  8.850 1.280 9.130 3.300 ;
        RECT  8.820 1.280 9.130 1.680 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.410 0.480 2.430 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.180 0.450 2.750 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.860 3.550 2.870 ;
        RECT  3.210 2.180 3.550 2.580 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.430 2.790 7.890 3.190 ;
        RECT  7.610 1.280 7.890 3.300 ;
        RECT  7.430 1.280 7.890 1.680 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.310 -0.380 6.710 0.560 ;
        RECT  8.000 -0.380 8.400 0.560 ;
        RECT  0.000 -0.380 9.300 0.380 ;
        RECT  1.260 -0.380 2.330 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 4.480 2.940 5.420 ;
        RECT  6.630 4.480 7.030 5.420 ;
        RECT  8.070 4.180 8.470 5.420 ;
        RECT  0.000 4.660 9.300 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.830 2.760 6.440 3.000 ;
        RECT  5.830 0.800 6.070 3.000 ;
        RECT  8.250 2.150 8.580 2.550 ;
        RECT  8.250 0.800 8.490 2.550 ;
        RECT  5.830 1.460 6.440 1.700 ;
        RECT  5.830 0.800 8.490 1.040 ;
        RECT  4.760 4.180 6.250 4.420 ;
        RECT  6.950 2.020 7.190 4.230 ;
        RECT  6.010 3.990 7.190 4.230 ;
        RECT  4.760 0.620 5.000 4.420 ;
        RECT  1.940 2.870 2.340 3.110 ;
        RECT  2.020 1.310 2.260 3.110 ;
        RECT  2.250 0.800 2.490 1.550 ;
        RECT  2.250 0.800 2.810 1.040 ;
        RECT  4.630 0.620 5.000 1.020 ;
        RECT  2.570 0.620 5.000 0.860 ;
        RECT  5.350 3.700 5.750 3.940 ;
        RECT  5.350 0.620 5.590 3.940 ;
        RECT  4.280 1.750 4.520 4.420 ;
        RECT  1.690 3.360 1.930 3.760 ;
        RECT  1.690 3.430 4.520 3.670 ;
        RECT  3.790 1.210 4.030 3.190 ;
        RECT  1.200 4.000 3.920 4.240 ;
        RECT  1.200 2.790 1.440 4.240 ;
        RECT  1.260 1.350 1.500 3.030 ;
        RECT  0.160 3.910 0.560 4.380 ;
        RECT  0.160 3.910 0.960 4.150 ;
        RECT  0.720 2.050 0.960 4.150 ;
        RECT  0.780 0.670 1.020 2.290 ;
        RECT  0.780 0.870 1.880 1.110 ;
        RECT  0.190 0.670 1.020 0.910 ;
    END
END DBHRBN

MACRO DBHRBS
    CLASS CORE ;
    FOREIGN DBHRBS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.300 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.760 2.930 2.700 ;
        RECT  2.500 2.050 2.930 2.450 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.820 2.790 9.130 3.190 ;
        RECT  8.850 1.280 9.130 3.300 ;
        RECT  8.820 1.280 9.130 1.680 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.410 0.480 2.430 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.180 0.450 2.750 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.860 3.550 2.870 ;
        RECT  3.210 2.180 3.550 2.580 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.430 2.790 7.890 3.190 ;
        RECT  7.610 1.280 7.890 3.300 ;
        RECT  7.430 1.280 7.890 1.680 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.310 -0.380 6.710 0.560 ;
        RECT  7.950 -0.380 8.350 0.560 ;
        RECT  0.000 -0.380 9.300 0.380 ;
        RECT  1.260 -0.380 2.330 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 4.480 2.940 5.420 ;
        RECT  6.630 4.480 7.030 5.420 ;
        RECT  7.950 4.180 8.350 5.420 ;
        RECT  0.000 4.660 9.300 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.830 2.760 6.440 3.000 ;
        RECT  5.830 0.800 6.070 3.000 ;
        RECT  8.250 2.150 8.580 2.550 ;
        RECT  8.250 0.800 8.490 2.550 ;
        RECT  5.830 1.460 6.440 1.700 ;
        RECT  5.830 0.800 8.490 1.040 ;
        RECT  4.760 4.180 6.250 4.420 ;
        RECT  6.950 2.020 7.190 4.230 ;
        RECT  6.010 3.990 7.190 4.230 ;
        RECT  4.760 0.620 5.000 4.420 ;
        RECT  1.940 2.870 2.340 3.110 ;
        RECT  2.020 1.310 2.260 3.110 ;
        RECT  2.250 0.800 2.490 1.550 ;
        RECT  2.250 0.800 2.810 1.040 ;
        RECT  4.630 0.620 5.000 1.020 ;
        RECT  2.570 0.620 5.000 0.860 ;
        RECT  5.350 3.700 5.750 3.940 ;
        RECT  5.350 0.620 5.590 3.940 ;
        RECT  4.280 1.750 4.520 4.420 ;
        RECT  1.690 3.360 1.930 3.760 ;
        RECT  1.690 3.430 4.520 3.670 ;
        RECT  3.790 1.210 4.030 3.190 ;
        RECT  1.200 4.000 3.920 4.240 ;
        RECT  1.200 2.790 1.440 4.240 ;
        RECT  1.260 1.350 1.500 3.030 ;
        RECT  0.160 3.910 0.560 4.380 ;
        RECT  0.160 3.910 0.960 4.150 ;
        RECT  0.720 2.050 0.960 4.150 ;
        RECT  0.780 0.670 1.020 2.290 ;
        RECT  0.780 0.870 1.880 1.110 ;
        RECT  0.190 0.670 1.020 0.910 ;
    END
END DBHRBS

MACRO DBZRBN
    CLASS CORE ;
    FOREIGN DBZRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.470 2.540 ;
        RECT  10.090 1.930 10.370 2.650 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.270 2.310 2.670 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 1.300 14.710 3.840 ;
        RECT  14.370 3.440 14.710 3.840 ;
        RECT  14.370 1.300 14.710 1.700 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.300 13.470 3.400 ;
        RECT  13.140 3.000 13.470 3.400 ;
        RECT  13.140 1.300 13.470 1.700 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.380 4.650 0.560 ;
        RECT  10.110 -0.380 10.510 0.560 ;
        RECT  12.340 -0.380 12.740 0.860 ;
        RECT  13.570 -0.380 13.970 0.860 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 4.030 4.720 5.420 ;
        RECT  9.940 4.480 10.340 5.420 ;
        RECT  11.970 4.130 12.370 5.420 ;
        RECT  13.570 4.260 13.970 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  2.090 4.480 2.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 4.180 7.760 4.420 ;
        RECT  7.520 3.580 7.760 4.420 ;
        RECT  6.320 0.780 6.560 4.420 ;
        RECT  6.240 3.620 6.560 4.020 ;
        RECT  12.580 3.720 14.120 3.960 ;
        RECT  13.880 2.140 14.120 3.960 ;
        RECT  7.520 3.580 10.850 3.820 ;
        RECT  10.610 2.880 10.850 3.820 ;
        RECT  12.580 1.100 12.820 3.960 ;
        RECT  10.610 2.880 12.820 3.120 ;
        RECT  11.770 1.100 12.820 1.340 ;
        RECT  6.240 0.780 6.560 1.180 ;
        RECT  11.770 0.620 12.010 1.340 ;
        RECT  11.620 0.620 12.020 0.860 ;
        RECT  12.100 1.640 12.340 2.540 ;
        RECT  11.520 1.640 12.340 1.880 ;
        RECT  11.520 1.580 11.920 1.880 ;
        RECT  10.870 4.090 11.390 4.330 ;
        RECT  11.150 3.420 11.390 4.330 ;
        RECT  11.150 3.420 12.320 3.660 ;
        RECT  6.800 3.700 7.280 3.940 ;
        RECT  6.800 1.100 7.040 3.940 ;
        RECT  10.830 2.120 11.690 2.360 ;
        RECT  10.830 1.120 11.070 2.360 ;
        RECT  8.680 1.120 11.070 1.360 ;
        RECT  6.800 1.100 8.920 1.340 ;
        RECT  7.170 0.860 7.570 1.340 ;
        RECT  9.440 0.620 9.840 0.880 ;
        RECT  8.040 0.620 9.840 0.860 ;
        RECT  9.590 1.600 9.830 3.220 ;
        RECT  8.000 2.880 9.830 3.120 ;
        RECT  8.000 1.600 9.830 1.840 ;
        RECT  8.000 1.580 8.400 1.840 ;
        RECT  8.050 4.160 9.680 4.400 ;
        RECT  7.280 2.880 7.680 3.120 ;
        RECT  7.360 1.580 7.600 3.120 ;
        RECT  7.360 2.220 8.680 2.460 ;
        RECT  7.280 1.580 7.680 1.820 ;
        RECT  5.840 1.500 6.080 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  5.700 1.020 5.940 1.740 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  2.970 1.100 3.830 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  3.590 1.020 5.940 1.260 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.120 3.950 5.900 4.350 ;
        RECT  5.120 1.500 5.360 4.350 ;
        RECT  5.120 2.040 5.550 2.440 ;
        RECT  3.600 4.030 4.000 4.270 ;
        RECT  3.760 3.540 4.000 4.270 ;
        RECT  3.760 3.540 4.800 3.780 ;
        RECT  4.560 1.580 4.800 3.780 ;
        RECT  4.560 3.070 4.870 3.470 ;
        RECT  3.600 1.580 4.800 1.820 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.280 3.700 ;
        RECT  2.880 3.940 3.280 4.420 ;
        RECT  1.230 3.940 3.280 4.180 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
    END
END DBZRBN

MACRO DBZRSBN
    CLASS CORE ;
    FOREIGN DBZRSBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.740 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.140 12.230 3.210 ;
        RECT  11.560 2.140 12.230 2.540 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.270 2.310 2.670 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 1.300 16.570 3.840 ;
        RECT  16.260 3.440 16.570 3.840 ;
        RECT  16.260 1.300 16.570 1.700 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.050 1.300 15.330 3.400 ;
        RECT  15.030 3.000 15.330 3.400 ;
        RECT  15.030 1.300 15.330 1.700 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.960 1.620 11.200 2.450 ;
        RECT  9.230 2.210 11.200 2.450 ;
        RECT  11.960 1.100 12.200 1.860 ;
        RECT  10.960 1.620 12.200 1.860 ;
        RECT  11.960 1.100 13.470 1.340 ;
        RECT  13.190 1.100 13.470 2.210 ;
        RECT  9.230 2.140 9.470 2.540 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.380 4.650 0.560 ;
        RECT  10.840 -0.380 11.240 0.560 ;
        RECT  14.230 -0.380 14.630 0.860 ;
        RECT  15.460 -0.380 15.860 0.860 ;
        RECT  0.000 -0.380 16.740 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 4.030 4.720 5.420 ;
        RECT  11.270 4.480 11.670 5.420 ;
        RECT  13.990 4.130 14.390 5.420 ;
        RECT  15.460 4.260 15.860 5.420 ;
        RECT  0.000 4.660 16.740 5.420 ;
        RECT  2.090 4.480 2.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 4.180 7.760 4.420 ;
        RECT  7.520 3.580 7.760 4.420 ;
        RECT  6.320 0.620 6.560 4.420 ;
        RECT  6.240 3.620 6.560 4.020 ;
        RECT  14.550 3.690 16.010 3.930 ;
        RECT  15.770 2.140 16.010 3.930 ;
        RECT  10.290 3.580 12.710 3.820 ;
        RECT  12.470 2.940 12.710 3.820 ;
        RECT  7.520 3.580 9.160 3.820 ;
        RECT  14.550 1.100 14.790 3.930 ;
        RECT  8.920 3.360 10.530 3.600 ;
        RECT  12.470 2.940 14.790 3.180 ;
        RECT  13.750 1.100 14.790 1.340 ;
        RECT  13.750 0.620 13.990 1.340 ;
        RECT  12.950 0.620 13.990 0.860 ;
        RECT  6.160 0.620 6.560 0.860 ;
        RECT  12.590 2.450 14.310 2.690 ;
        RECT  14.070 2.140 14.310 2.690 ;
        RECT  12.590 1.580 12.830 2.690 ;
        RECT  12.440 1.580 12.840 1.820 ;
        RECT  12.200 4.090 13.190 4.330 ;
        RECT  12.950 3.480 13.190 4.330 ;
        RECT  12.950 3.480 14.210 3.720 ;
        RECT  6.800 3.700 7.280 3.940 ;
        RECT  6.800 1.100 7.040 3.940 ;
        RECT  8.690 1.120 11.720 1.360 ;
        RECT  11.480 0.620 11.720 1.360 ;
        RECT  6.800 1.100 8.930 1.340 ;
        RECT  7.170 0.860 7.570 1.340 ;
        RECT  11.480 0.620 12.570 0.860 ;
        RECT  10.920 2.820 11.160 3.220 ;
        RECT  8.000 2.880 11.160 3.120 ;
        RECT  8.750 1.600 8.990 3.120 ;
        RECT  8.000 1.600 10.520 1.840 ;
        RECT  8.000 1.580 8.400 1.840 ;
        RECT  8.050 4.160 11.010 4.400 ;
        RECT  9.530 3.840 9.930 4.400 ;
        RECT  10.200 0.620 10.600 0.880 ;
        RECT  8.040 0.620 10.600 0.860 ;
        RECT  7.280 2.880 7.680 3.120 ;
        RECT  7.360 1.580 7.600 3.120 ;
        RECT  8.270 2.140 8.510 2.540 ;
        RECT  7.360 2.220 8.510 2.460 ;
        RECT  7.280 1.580 7.680 1.820 ;
        RECT  5.840 1.290 6.080 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.680 1.020 5.920 1.530 ;
        RECT  2.970 1.100 3.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  3.700 1.020 5.920 1.260 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.120 3.950 5.900 4.350 ;
        RECT  5.120 1.500 5.360 4.350 ;
        RECT  5.120 2.040 5.550 2.440 ;
        RECT  3.600 4.030 4.000 4.270 ;
        RECT  3.760 3.540 4.000 4.270 ;
        RECT  3.760 3.540 4.800 3.780 ;
        RECT  4.560 1.580 4.800 3.780 ;
        RECT  4.560 3.100 4.870 3.500 ;
        RECT  3.600 1.580 4.800 1.820 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.280 3.700 ;
        RECT  2.880 3.940 3.280 4.420 ;
        RECT  1.230 3.940 3.280 4.180 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
    END
END DBZRSBN

MACRO DELA
    CLASS CORE ;
    FOREIGN DELA 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 3.460 4.790 3.860 ;
        RECT  4.510 1.100 4.790 4.020 ;
        RECT  4.480 1.100 4.790 1.500 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.210 0.480 2.610 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 -0.380 4.010 0.570 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.950 -0.380 1.350 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.620 4.260 4.020 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.400 3.670 4.150 3.910 ;
        RECT  3.910 0.850 4.150 3.910 ;
        RECT  2.400 0.850 4.150 1.090 ;
        RECT  2.180 1.490 2.420 3.220 ;
        RECT  2.180 2.240 3.360 2.480 ;
        RECT  0.160 3.720 1.880 3.960 ;
        RECT  1.640 1.150 1.880 3.960 ;
        RECT  0.160 1.150 1.880 1.390 ;
    END
END DELA

MACRO DELB
    CLASS CORE ;
    FOREIGN DELB 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 3.460 4.790 3.860 ;
        RECT  4.510 1.100 4.790 4.020 ;
        RECT  4.480 1.100 4.790 1.500 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.210 0.480 2.610 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 -0.380 4.010 0.570 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.950 -0.380 1.350 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.620 4.260 4.020 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.400 3.670 4.150 3.910 ;
        RECT  3.910 0.850 4.150 3.910 ;
        RECT  2.400 0.850 4.150 1.090 ;
        RECT  2.180 1.490 2.420 3.220 ;
        RECT  2.180 2.240 3.360 2.480 ;
        RECT  0.160 3.720 1.880 3.960 ;
        RECT  1.640 1.150 1.880 3.960 ;
        RECT  0.160 1.150 1.880 1.390 ;
    END
END DELB

MACRO DELC
    CLASS CORE ;
    FOREIGN DELC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 3.460 4.790 3.860 ;
        RECT  4.510 1.100 4.790 4.020 ;
        RECT  4.480 1.100 4.790 1.500 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.210 0.480 2.610 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 -0.380 4.010 0.570 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.950 -0.380 1.350 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.620 4.260 4.020 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.400 3.670 4.150 3.910 ;
        RECT  3.910 0.850 4.150 3.910 ;
        RECT  2.400 0.850 4.150 1.090 ;
        RECT  2.180 1.490 2.420 3.220 ;
        RECT  2.180 2.240 3.360 2.480 ;
        RECT  0.160 3.720 1.880 3.960 ;
        RECT  1.640 1.150 1.880 3.960 ;
        RECT  0.160 1.150 1.880 1.390 ;
    END
END DELC

MACRO DFCLRBN
    CLASS CORE ;
    FOREIGN DFCLRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.800 ;
        RECT  1.870 2.100 2.310 2.500 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 2.120 6.030 2.840 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.590 2.880 15.950 3.280 ;
        RECT  15.670 1.260 15.950 3.370 ;
        RECT  15.590 1.340 15.950 1.740 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.060 3.550 2.710 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.190 0.620 14.470 1.320 ;
        RECT  14.430 1.040 14.710 3.190 ;
        RECT  14.150 2.790 14.710 3.190 ;
        RECT  14.070 0.620 14.470 0.860 ;
        END
    END Q
    PIN LD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.810 1.620 2.790 1.860 ;
        RECT  2.550 1.620 2.790 3.430 ;
        RECT  3.900 2.260 4.140 3.430 ;
        RECT  2.550 3.190 4.140 3.430 ;
        RECT  3.900 2.260 4.200 2.660 ;
        RECT  0.810 1.620 1.050 2.800 ;
        END
    END LD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.000 -0.380 6.400 0.560 ;
        RECT  6.840 -0.380 7.240 0.560 ;
        RECT  10.070 -0.380 10.470 0.860 ;
        RECT  13.070 -0.380 13.470 0.560 ;
        RECT  14.790 -0.380 15.190 0.800 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  1.420 -0.380 1.820 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.290 4.200 2.690 5.420 ;
        RECT  4.960 4.480 5.360 5.420 ;
        RECT  6.110 4.480 6.510 5.420 ;
        RECT  10.160 4.200 10.560 5.420 ;
        RECT  13.220 4.400 13.460 5.420 ;
        RECT  14.790 4.260 15.190 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  0.960 3.040 1.200 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.380 4.180 12.980 4.420 ;
        RECT  12.740 3.720 12.980 4.420 ;
        RECT  7.190 4.180 9.480 4.420 ;
        RECT  9.240 3.720 9.480 4.420 ;
        RECT  4.920 4.000 7.430 4.240 ;
        RECT  11.380 3.720 11.620 4.420 ;
        RECT  8.120 0.620 8.360 4.420 ;
        RECT  4.920 2.250 5.160 4.240 ;
        RECT  12.740 3.720 15.300 3.960 ;
        RECT  15.060 2.160 15.300 3.960 ;
        RECT  9.240 3.720 11.620 3.960 ;
        RECT  7.670 3.700 8.360 3.940 ;
        RECT  13.640 3.530 13.890 3.960 ;
        RECT  13.650 1.320 13.890 3.960 ;
        RECT  13.640 1.320 13.890 1.720 ;
        RECT  7.610 0.620 8.360 0.860 ;
        RECT  12.260 3.200 12.500 3.940 ;
        RECT  12.260 3.200 13.330 3.440 ;
        RECT  13.090 0.890 13.330 3.440 ;
        RECT  13.090 2.160 13.410 2.560 ;
        RECT  12.260 0.890 13.330 1.130 ;
        RECT  12.260 0.730 12.500 1.130 ;
        RECT  8.600 3.700 9.000 3.940 ;
        RECT  8.600 0.620 8.840 3.940 ;
        RECT  11.750 1.100 11.990 3.200 ;
        RECT  11.750 2.210 12.570 2.450 ;
        RECT  9.530 1.100 11.990 1.340 ;
        RECT  9.530 0.620 9.770 1.340 ;
        RECT  8.600 0.620 9.770 0.860 ;
        RECT  9.990 2.880 11.430 3.120 ;
        RECT  11.190 1.580 11.430 3.120 ;
        RECT  9.990 2.260 10.230 3.120 ;
        RECT  10.950 1.580 11.430 1.820 ;
        RECT  9.080 1.500 9.320 3.200 ;
        RECT  10.470 2.170 10.950 2.570 ;
        RECT  10.470 1.730 10.710 2.570 ;
        RECT  9.080 1.730 10.710 1.970 ;
        RECT  1.470 3.720 1.710 4.160 ;
        RECT  1.470 3.720 4.680 3.960 ;
        RECT  4.440 1.100 4.680 3.960 ;
        RECT  7.640 1.100 7.880 3.200 ;
        RECT  3.510 1.100 7.880 1.340 ;
        RECT  6.900 3.520 7.300 3.760 ;
        RECT  6.980 1.580 7.220 3.760 ;
        RECT  6.980 2.240 7.340 2.640 ;
        RECT  6.840 1.580 7.240 1.820 ;
        RECT  5.460 3.520 6.590 3.760 ;
        RECT  6.350 1.580 6.590 3.760 ;
        RECT  6.350 2.900 6.690 3.300 ;
        RECT  6.000 1.580 6.590 1.820 ;
        RECT  2.140 0.620 5.190 0.860 ;
        RECT  0.240 4.020 0.720 4.420 ;
        RECT  0.240 1.100 0.480 4.420 ;
        RECT  3.960 1.580 4.200 1.980 ;
        RECT  3.030 1.580 4.200 1.820 ;
        RECT  3.030 1.100 3.270 1.820 ;
        RECT  0.240 1.100 3.270 1.340 ;
    END
END DFCLRBN

MACRO DFCRBN
    CLASS CORE ;
    FOREIGN DFCRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.690 2.840 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.230 2.550 2.630 ;
        RECT  2.030 2.120 2.310 2.840 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 1.090 12.850 3.280 ;
        RECT  12.490 2.880 12.850 3.280 ;
        RECT  12.490 1.200 12.850 1.600 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.230 0.690 2.630 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.270 1.280 11.670 3.110 ;
        RECT  10.970 2.870 11.670 3.110 ;
        RECT  10.970 1.280 11.670 1.520 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.760 -0.380 3.160 0.560 ;
        RECT  6.810 -0.380 7.210 0.860 ;
        RECT  9.720 -0.380 10.120 0.560 ;
        RECT  11.690 -0.380 12.090 0.800 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  1.830 -0.380 2.230 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.760 4.260 3.160 5.420 ;
        RECT  6.810 4.200 7.210 5.420 ;
        RECT  9.870 4.400 10.110 5.420 ;
        RECT  11.690 4.260 12.090 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.030 4.180 9.630 4.420 ;
        RECT  9.390 3.720 9.630 4.420 ;
        RECT  4.770 4.180 6.130 4.420 ;
        RECT  5.890 3.720 6.130 4.420 ;
        RECT  8.030 3.720 8.270 4.420 ;
        RECT  4.770 0.620 5.010 4.420 ;
        RECT  9.390 3.720 12.240 3.960 ;
        RECT  12.000 2.160 12.240 3.960 ;
        RECT  5.890 3.720 8.270 3.960 ;
        RECT  4.320 3.700 5.010 3.940 ;
        RECT  10.300 3.530 10.570 3.960 ;
        RECT  10.300 1.320 10.540 3.960 ;
        RECT  10.300 1.320 10.570 1.720 ;
        RECT  4.260 0.620 5.010 0.860 ;
        RECT  8.910 3.200 9.150 3.940 ;
        RECT  8.910 3.200 10.060 3.440 ;
        RECT  9.820 0.890 10.060 3.440 ;
        RECT  8.910 0.890 10.060 1.130 ;
        RECT  8.910 0.730 9.150 1.130 ;
        RECT  5.250 3.700 5.650 3.940 ;
        RECT  5.250 0.620 5.490 3.940 ;
        RECT  8.400 1.100 8.640 3.200 ;
        RECT  8.400 2.210 9.220 2.450 ;
        RECT  6.180 1.100 8.640 1.340 ;
        RECT  6.180 0.620 6.420 1.340 ;
        RECT  5.250 0.620 6.420 0.860 ;
        RECT  6.640 2.880 8.160 3.120 ;
        RECT  7.920 1.580 8.160 3.120 ;
        RECT  6.640 2.260 6.880 3.120 ;
        RECT  7.600 1.580 8.160 1.820 ;
        RECT  5.730 1.500 5.970 3.200 ;
        RECT  7.120 2.170 7.600 2.570 ;
        RECT  7.120 1.730 7.360 2.570 ;
        RECT  5.730 1.730 7.360 1.970 ;
        RECT  1.550 4.180 2.000 4.420 ;
        RECT  1.550 3.400 1.790 4.420 ;
        RECT  0.160 3.400 1.790 3.640 ;
        RECT  0.930 0.800 1.170 3.640 ;
        RECT  4.290 1.100 4.530 3.200 ;
        RECT  2.890 1.100 4.530 1.340 ;
        RECT  2.890 0.800 3.130 1.340 ;
        RECT  0.160 0.800 3.130 1.040 ;
        RECT  3.550 3.500 3.950 3.740 ;
        RECT  3.630 1.580 3.870 3.740 ;
        RECT  3.630 2.290 4.000 2.690 ;
        RECT  3.490 1.580 3.890 1.820 ;
        RECT  2.110 3.460 3.240 3.700 ;
        RECT  3.000 1.580 3.240 3.700 ;
        RECT  3.000 2.840 3.340 3.240 ;
        RECT  2.110 1.580 3.240 1.820 ;
    END
END DFCRBN

MACRO DFFN
    CLASS CORE ;
    FOREIGN DFFN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.970 2.230 2.310 2.630 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.710 1.480 10.990 3.200 ;
        RECT  10.680 2.800 10.990 3.200 ;
        RECT  10.680 1.480 10.990 1.880 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.660 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.360 0.620 9.640 1.540 ;
        RECT  9.470 1.260 9.750 3.200 ;
        RECT  9.240 2.800 9.750 3.200 ;
        RECT  9.240 0.620 9.640 1.020 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.310 -0.380 2.710 0.560 ;
        RECT  7.890 -0.380 8.130 0.640 ;
        RECT  9.880 -0.380 10.280 0.940 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.910 -0.380 1.310 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 4.040 2.780 5.420 ;
        RECT  5.970 4.480 6.370 5.420 ;
        RECT  7.680 4.480 8.080 5.420 ;
        RECT  9.880 4.260 10.280 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.190 4.260 0.590 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.650 3.850 9.050 4.090 ;
        RECT  10.180 2.160 10.420 4.020 ;
        RECT  8.730 3.780 10.420 4.020 ;
        RECT  8.730 1.370 8.970 4.090 ;
        RECT  7.890 2.480 8.970 2.720 ;
        RECT  7.360 0.890 8.820 1.130 ;
        RECT  8.420 0.730 8.820 1.130 ;
        RECT  4.800 0.620 5.040 1.020 ;
        RECT  7.360 0.620 7.600 1.130 ;
        RECT  4.800 0.620 7.600 0.860 ;
        RECT  4.720 4.000 8.380 4.240 ;
        RECT  8.140 3.080 8.380 4.240 ;
        RECT  4.000 3.520 4.240 4.160 ;
        RECT  4.000 3.520 7.780 3.760 ;
        RECT  7.410 1.660 7.650 3.760 ;
        RECT  4.320 0.620 4.560 3.760 ;
        RECT  7.350 1.660 7.650 2.060 ;
        RECT  3.810 0.620 4.560 0.860 ;
        RECT  5.790 3.040 7.110 3.280 ;
        RECT  6.870 1.100 7.110 3.280 ;
        RECT  5.790 2.120 6.030 3.280 ;
        RECT  5.630 2.120 6.030 2.360 ;
        RECT  6.560 1.100 7.110 1.340 ;
        RECT  4.800 1.500 5.040 3.200 ;
        RECT  6.290 2.260 6.630 2.660 ;
        RECT  6.290 1.580 6.530 2.660 ;
        RECT  4.800 1.580 6.530 1.820 ;
        RECT  0.940 3.240 1.230 3.640 ;
        RECT  0.940 1.100 1.180 3.640 ;
        RECT  3.840 1.100 4.080 3.200 ;
        RECT  0.190 1.100 4.080 1.340 ;
        RECT  3.180 1.580 3.420 4.360 ;
        RECT  3.040 1.580 3.440 1.820 ;
        RECT  1.660 4.040 2.130 4.280 ;
        RECT  1.890 3.560 2.130 4.280 ;
        RECT  1.890 3.560 2.930 3.800 ;
        RECT  2.550 3.400 2.930 3.800 ;
        RECT  2.550 1.580 2.790 3.800 ;
        RECT  1.660 1.580 2.790 1.820 ;
    END
END DFFN

MACRO DFFP
    CLASS CORE ;
    FOREIGN DFFP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.640 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.230 1.930 2.630 ;
        RECT  1.410 2.120 1.690 2.840 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.140 1.260 13.520 3.220 ;
        RECT  12.320 2.940 13.520 3.220 ;
        RECT  12.320 1.260 13.520 1.540 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.550 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.650 1.280 11.280 1.520 ;
        RECT  10.650 2.960 11.280 3.200 ;
        RECT  10.650 1.280 11.050 3.200 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.040 -0.380 2.440 0.560 ;
        RECT  6.190 -0.380 6.590 0.860 ;
        RECT  9.100 -0.380 9.500 0.560 ;
        RECT  10.160 -0.380 10.560 0.800 ;
        RECT  11.600 -0.380 12.000 0.800 ;
        RECT  13.040 -0.380 13.440 0.800 ;
        RECT  0.000 -0.380 13.640 0.380 ;
        RECT  0.880 -0.380 1.280 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.110 4.180 2.510 5.420 ;
        RECT  6.190 4.200 6.590 5.420 ;
        RECT  9.250 4.400 9.490 5.420 ;
        RECT  10.160 4.260 10.560 5.420 ;
        RECT  11.600 4.260 12.000 5.420 ;
        RECT  13.040 4.260 13.440 5.420 ;
        RECT  0.000 4.660 13.640 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.410 4.180 9.010 4.420 ;
        RECT  8.770 3.720 9.010 4.420 ;
        RECT  4.050 4.180 5.410 4.420 ;
        RECT  5.170 3.720 5.410 4.420 ;
        RECT  7.410 3.720 7.650 4.420 ;
        RECT  4.050 0.620 4.290 4.420 ;
        RECT  8.770 3.720 12.050 3.960 ;
        RECT  11.810 2.240 12.050 3.960 ;
        RECT  5.170 3.720 7.650 3.960 ;
        RECT  3.600 3.700 4.290 3.940 ;
        RECT  9.680 1.320 9.920 3.960 ;
        RECT  9.680 2.810 9.970 3.210 ;
        RECT  11.810 2.240 12.590 2.480 ;
        RECT  9.680 1.320 9.970 1.720 ;
        RECT  3.540 0.620 4.290 0.860 ;
        RECT  8.290 3.200 8.530 3.940 ;
        RECT  8.290 3.200 9.420 3.440 ;
        RECT  9.180 0.800 9.420 3.440 ;
        RECT  9.180 2.160 9.440 2.560 ;
        RECT  8.290 0.720 8.530 1.120 ;
        RECT  8.290 0.800 9.420 1.040 ;
        RECT  4.530 3.700 4.930 3.940 ;
        RECT  4.530 0.620 4.770 3.940 ;
        RECT  7.780 1.100 8.020 3.200 ;
        RECT  7.780 2.210 8.600 2.450 ;
        RECT  5.560 1.100 8.020 1.340 ;
        RECT  5.560 0.620 5.800 1.340 ;
        RECT  4.530 0.620 5.800 0.860 ;
        RECT  5.960 2.880 7.540 3.120 ;
        RECT  7.300 1.580 7.540 3.120 ;
        RECT  5.960 2.260 6.200 3.120 ;
        RECT  6.980 1.580 7.540 1.820 ;
        RECT  5.010 1.500 5.250 3.200 ;
        RECT  6.500 2.170 6.980 2.570 ;
        RECT  6.500 1.730 6.740 2.570 ;
        RECT  5.010 1.730 6.740 1.970 ;
        RECT  0.880 3.380 1.200 3.780 ;
        RECT  0.880 1.100 1.120 3.780 ;
        RECT  3.570 1.100 3.810 3.200 ;
        RECT  0.320 1.100 3.810 1.340 ;
        RECT  0.320 0.640 0.560 1.340 ;
        RECT  0.160 0.640 0.560 0.880 ;
        RECT  2.830 4.180 3.230 4.420 ;
        RECT  2.910 1.580 3.150 4.420 ;
        RECT  2.770 1.580 3.170 1.820 ;
        RECT  1.390 4.180 1.790 4.420 ;
        RECT  1.550 3.700 1.790 4.420 ;
        RECT  1.550 3.700 2.520 3.940 ;
        RECT  2.280 1.580 2.520 3.940 ;
        RECT  2.280 3.220 2.660 3.620 ;
        RECT  1.390 1.580 2.520 1.820 ;
    END
END DFFP

MACRO DFFRBN
    CLASS CORE ;
    FOREIGN DFFRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.140 8.610 2.540 ;
        RECT  8.230 1.930 8.510 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 1.300 12.850 3.840 ;
        RECT  12.510 3.440 12.850 3.840 ;
        RECT  12.510 1.300 12.850 1.700 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.140 1.080 2.540 ;
        RECT  0.790 2.120 1.070 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 1.300 11.610 3.400 ;
        RECT  11.280 3.000 11.610 3.400 ;
        RECT  11.280 1.300 11.610 1.700 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  8.250 -0.380 8.650 0.560 ;
        RECT  10.480 -0.380 10.880 0.860 ;
        RECT  11.710 -0.380 12.110 0.860 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  1.100 -0.380 2.790 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.670 4.020 3.070 5.420 ;
        RECT  8.080 4.480 8.480 5.420 ;
        RECT  10.110 4.130 10.510 5.420 ;
        RECT  11.710 4.260 12.110 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.460 4.180 5.900 4.420 ;
        RECT  5.660 3.580 5.900 4.420 ;
        RECT  4.460 0.620 4.700 4.420 ;
        RECT  4.380 3.620 4.700 4.020 ;
        RECT  10.720 3.720 12.260 3.960 ;
        RECT  12.020 2.140 12.260 3.960 ;
        RECT  5.660 3.580 9.000 3.820 ;
        RECT  8.760 2.880 9.000 3.820 ;
        RECT  10.720 1.100 10.960 3.960 ;
        RECT  8.760 2.880 10.960 3.120 ;
        RECT  9.920 1.100 10.960 1.340 ;
        RECT  9.920 0.620 10.160 1.340 ;
        RECT  9.760 0.620 10.160 0.860 ;
        RECT  4.300 0.620 4.700 0.860 ;
        RECT  10.240 1.640 10.480 2.540 ;
        RECT  9.660 1.640 10.480 1.880 ;
        RECT  9.660 1.580 10.060 1.880 ;
        RECT  9.010 4.090 9.530 4.330 ;
        RECT  9.290 3.540 9.530 4.330 ;
        RECT  9.290 3.540 10.460 3.780 ;
        RECT  4.940 3.700 5.420 3.940 ;
        RECT  4.940 1.100 5.180 3.940 ;
        RECT  8.980 2.120 9.830 2.360 ;
        RECT  8.980 1.120 9.220 2.360 ;
        RECT  6.830 1.120 9.220 1.360 ;
        RECT  4.940 1.100 7.070 1.340 ;
        RECT  5.310 0.860 5.710 1.340 ;
        RECT  7.580 0.620 7.980 0.880 ;
        RECT  6.180 0.620 7.980 0.860 ;
        RECT  7.730 1.600 7.970 3.220 ;
        RECT  6.140 2.880 7.970 3.120 ;
        RECT  6.140 1.600 7.970 1.840 ;
        RECT  6.140 1.580 6.540 1.840 ;
        RECT  6.190 4.160 7.820 4.400 ;
        RECT  5.420 2.880 5.820 3.120 ;
        RECT  5.500 1.580 5.740 3.120 ;
        RECT  5.500 2.220 6.820 2.460 ;
        RECT  5.420 1.580 5.820 1.820 ;
        RECT  3.980 1.290 4.220 3.200 ;
        RECT  0.190 2.800 0.480 3.200 ;
        RECT  0.190 1.010 0.430 3.200 ;
        RECT  3.840 1.010 4.080 1.530 ;
        RECT  0.160 1.010 4.080 1.250 ;
        RECT  3.390 4.020 3.790 4.260 ;
        RECT  3.390 3.430 3.630 4.260 ;
        RECT  3.260 1.580 3.500 3.670 ;
        RECT  3.260 2.260 3.690 2.660 ;
        RECT  3.180 1.580 3.580 1.820 ;
        RECT  1.740 3.540 2.940 3.780 ;
        RECT  2.700 1.580 2.940 3.780 ;
        RECT  2.700 2.260 3.010 2.660 ;
        RECT  1.740 1.580 2.940 1.820 ;
    END
END DFFRBN

MACRO DFFRBP
    CLASS CORE ;
    FOREIGN DFFRBP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.930 8.510 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.230 2.310 2.630 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.280 13.470 3.260 ;
        RECT  12.950 2.860 13.470 3.260 ;
        RECT  12.950 1.280 13.470 1.680 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.120 1.070 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 1.260 12.230 3.220 ;
        RECT  11.430 2.940 12.230 3.220 ;
        RECT  11.430 1.260 12.230 1.540 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  8.070 -0.380 8.470 0.560 ;
        RECT  10.710 -0.380 11.110 0.860 ;
        RECT  12.150 -0.380 12.550 0.860 ;
        RECT  13.590 -0.380 13.990 0.860 ;
        RECT  0.000 -0.380 14.260 0.380 ;
        RECT  1.090 -0.380 2.680 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 4.020 2.820 5.420 ;
        RECT  7.970 4.480 8.370 5.420 ;
        RECT  9.690 4.480 10.090 5.420 ;
        RECT  10.500 4.480 10.900 5.420 ;
        RECT  12.150 4.260 12.550 5.420 ;
        RECT  13.590 4.260 13.990 5.420 ;
        RECT  0.000 4.660 14.260 5.420 ;
        RECT  0.880 3.740 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.350 4.180 5.790 4.420 ;
        RECT  5.550 3.580 5.790 4.420 ;
        RECT  4.350 0.620 4.590 4.420 ;
        RECT  4.270 3.620 4.590 4.020 ;
        RECT  5.550 3.580 12.710 3.820 ;
        RECT  12.470 2.140 12.710 3.820 ;
        RECT  10.950 1.100 11.190 3.820 ;
        RECT  12.470 2.140 12.780 2.540 ;
        RECT  10.150 1.100 11.190 1.340 ;
        RECT  10.150 0.620 10.390 1.340 ;
        RECT  9.990 0.620 10.390 0.860 ;
        RECT  4.190 0.620 4.590 0.860 ;
        RECT  8.900 3.100 10.710 3.340 ;
        RECT  10.470 1.640 10.710 3.340 ;
        RECT  9.480 1.640 10.710 1.880 ;
        RECT  9.480 1.570 9.880 1.880 ;
        RECT  4.830 3.700 5.310 3.940 ;
        RECT  4.830 1.100 5.070 3.940 ;
        RECT  8.870 2.220 9.720 2.460 ;
        RECT  8.870 1.120 9.110 2.460 ;
        RECT  6.720 1.120 9.110 1.360 ;
        RECT  4.830 1.100 6.960 1.340 ;
        RECT  5.200 0.860 5.600 1.340 ;
        RECT  7.620 1.600 7.860 3.220 ;
        RECT  6.030 2.880 7.860 3.120 ;
        RECT  6.030 1.600 7.860 1.840 ;
        RECT  6.030 1.580 6.430 1.840 ;
        RECT  7.400 0.620 7.800 0.880 ;
        RECT  6.070 0.620 7.800 0.860 ;
        RECT  6.080 4.160 7.710 4.400 ;
        RECT  5.310 2.880 5.710 3.120 ;
        RECT  5.390 1.580 5.630 3.120 ;
        RECT  5.390 2.220 6.710 2.460 ;
        RECT  5.310 1.580 5.710 1.820 ;
        RECT  0.140 2.890 0.480 3.290 ;
        RECT  3.870 1.290 4.110 3.200 ;
        RECT  0.140 1.090 0.380 3.290 ;
        RECT  3.730 1.290 4.110 1.530 ;
        RECT  0.140 1.090 3.970 1.330 ;
        RECT  0.160 1.010 0.560 1.330 ;
        RECT  3.150 3.940 3.460 4.340 ;
        RECT  3.150 1.570 3.390 4.340 ;
        RECT  3.150 2.260 3.580 2.660 ;
        RECT  3.070 1.570 3.470 1.810 ;
        RECT  1.630 3.930 2.030 4.170 ;
        RECT  1.790 3.540 2.030 4.170 ;
        RECT  1.790 3.540 2.830 3.780 ;
        RECT  2.590 1.570 2.830 3.780 ;
        RECT  2.590 2.260 2.900 2.660 ;
        RECT  1.630 1.570 2.830 1.810 ;
    END
END DFFRBP

MACRO DFFRBS
    CLASS CORE ;
    FOREIGN DFFRBS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.140 8.610 2.540 ;
        RECT  8.230 1.930 8.510 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 0.650 12.850 4.100 ;
        RECT  12.510 3.700 12.850 4.100 ;
        RECT  12.510 0.650 12.850 1.050 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.140 1.080 2.540 ;
        RECT  0.790 2.120 1.070 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 1.400 11.610 3.190 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  8.250 -0.380 8.650 0.560 ;
        RECT  10.480 -0.380 10.880 0.860 ;
        RECT  11.710 -0.380 12.110 0.860 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  1.100 -0.380 2.790 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.670 4.020 3.070 5.420 ;
        RECT  8.080 4.480 8.480 5.420 ;
        RECT  10.110 4.130 10.510 5.420 ;
        RECT  11.710 4.260 12.110 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.460 4.180 5.900 4.420 ;
        RECT  5.660 3.580 5.900 4.420 ;
        RECT  4.460 0.620 4.700 4.420 ;
        RECT  4.380 3.620 4.700 4.020 ;
        RECT  10.720 3.720 12.260 3.960 ;
        RECT  12.020 2.140 12.260 3.960 ;
        RECT  5.660 3.580 9.000 3.820 ;
        RECT  8.760 2.880 9.000 3.820 ;
        RECT  10.720 1.100 10.960 3.960 ;
        RECT  8.760 2.880 10.960 3.120 ;
        RECT  9.920 1.100 10.960 1.340 ;
        RECT  9.920 0.620 10.160 1.340 ;
        RECT  9.760 0.620 10.160 0.860 ;
        RECT  4.300 0.620 4.700 0.860 ;
        RECT  10.240 1.640 10.480 2.540 ;
        RECT  9.660 1.640 10.480 1.880 ;
        RECT  9.660 1.580 10.060 1.880 ;
        RECT  9.010 4.090 9.530 4.330 ;
        RECT  9.290 3.580 9.530 4.330 ;
        RECT  9.290 3.580 10.460 3.820 ;
        RECT  4.940 3.700 5.420 3.940 ;
        RECT  4.940 1.100 5.180 3.940 ;
        RECT  8.980 2.120 9.830 2.360 ;
        RECT  8.980 1.120 9.220 2.360 ;
        RECT  6.830 1.120 9.220 1.360 ;
        RECT  4.940 1.100 7.070 1.340 ;
        RECT  5.310 0.860 5.710 1.340 ;
        RECT  7.580 0.620 7.980 0.880 ;
        RECT  6.180 0.620 7.980 0.860 ;
        RECT  7.730 1.600 7.970 3.220 ;
        RECT  6.140 2.880 7.970 3.120 ;
        RECT  6.140 1.600 7.970 1.840 ;
        RECT  6.140 1.580 6.540 1.840 ;
        RECT  6.190 4.160 7.820 4.400 ;
        RECT  5.420 2.880 5.820 3.120 ;
        RECT  5.500 1.580 5.740 3.120 ;
        RECT  5.500 2.220 6.820 2.460 ;
        RECT  5.420 1.580 5.820 1.820 ;
        RECT  3.980 1.290 4.220 3.200 ;
        RECT  0.190 2.800 0.480 3.200 ;
        RECT  0.190 1.010 0.430 3.200 ;
        RECT  3.840 1.010 4.080 1.530 ;
        RECT  0.160 1.010 4.080 1.250 ;
        RECT  3.390 4.020 3.790 4.260 ;
        RECT  3.390 3.430 3.630 4.260 ;
        RECT  3.260 1.580 3.500 3.670 ;
        RECT  3.260 2.260 3.690 2.660 ;
        RECT  3.180 1.580 3.580 1.820 ;
        RECT  1.740 3.540 2.940 3.780 ;
        RECT  2.700 1.580 2.940 3.780 ;
        RECT  2.700 2.260 3.010 2.660 ;
        RECT  1.740 1.580 2.940 1.820 ;
    END
END DFFRBS

MACRO DFFRBT
    CLASS CORE ;
    FOREIGN DFFRBT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.930 8.510 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.910 2.230 2.310 2.630 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.370 1.200 14.650 3.710 ;
        RECT  14.140 3.310 14.650 3.710 ;
        RECT  15.580 1.200 15.950 1.600 ;
        RECT  14.370 2.320 15.950 2.720 ;
        RECT  15.670 1.200 15.950 3.710 ;
        RECT  15.580 3.310 15.950 3.710 ;
        RECT  14.140 1.200 14.650 1.600 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.470 2.820 11.710 3.220 ;
        RECT  11.470 1.260 13.230 1.540 ;
        RECT  12.510 1.260 12.910 3.220 ;
        RECT  12.510 1.260 13.230 1.580 ;
        RECT  11.470 2.940 13.230 3.220 ;
        RECT  11.470 1.260 11.710 1.660 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.250 -0.380 2.650 0.560 ;
        RECT  8.090 -0.380 8.490 0.560 ;
        RECT  10.670 -0.380 11.070 0.860 ;
        RECT  12.110 -0.380 12.510 0.860 ;
        RECT  13.340 -0.380 13.740 0.860 ;
        RECT  14.780 -0.380 15.180 0.860 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  1.200 -0.380 1.600 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.020 2.720 5.420 ;
        RECT  8.070 4.480 8.470 5.420 ;
        RECT  9.650 4.480 10.050 5.420 ;
        RECT  10.470 4.480 10.870 5.420 ;
        RECT  12.110 4.260 12.510 5.420 ;
        RECT  13.340 4.260 13.740 5.420 ;
        RECT  14.780 4.260 15.180 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.320 4.180 5.760 4.420 ;
        RECT  5.520 3.580 5.760 4.420 ;
        RECT  4.320 0.620 4.560 4.420 ;
        RECT  4.240 3.620 4.560 4.020 ;
        RECT  5.520 3.580 13.890 3.820 ;
        RECT  13.650 2.140 13.890 3.820 ;
        RECT  10.990 1.100 11.230 3.820 ;
        RECT  10.110 1.100 11.230 1.340 ;
        RECT  10.110 0.620 10.350 1.340 ;
        RECT  9.950 0.620 10.350 0.860 ;
        RECT  4.160 0.620 4.560 0.860 ;
        RECT  8.860 3.100 10.750 3.340 ;
        RECT  10.510 1.640 10.750 3.340 ;
        RECT  9.440 1.640 10.750 1.880 ;
        RECT  9.440 1.570 9.840 1.880 ;
        RECT  4.800 3.700 5.280 3.940 ;
        RECT  4.800 1.100 5.040 3.940 ;
        RECT  8.840 2.220 9.690 2.460 ;
        RECT  8.840 1.120 9.080 2.460 ;
        RECT  6.690 1.120 9.080 1.360 ;
        RECT  4.800 1.100 6.930 1.340 ;
        RECT  5.170 0.860 5.570 1.340 ;
        RECT  7.590 2.820 7.830 3.220 ;
        RECT  6.000 2.880 7.830 3.120 ;
        RECT  7.510 1.600 7.750 3.120 ;
        RECT  6.000 1.600 7.750 1.840 ;
        RECT  6.000 1.580 6.400 1.840 ;
        RECT  7.350 0.620 7.750 0.880 ;
        RECT  6.040 0.620 7.750 0.860 ;
        RECT  6.050 4.160 7.680 4.400 ;
        RECT  5.280 2.880 5.680 3.120 ;
        RECT  5.360 1.580 5.600 3.120 ;
        RECT  5.360 2.220 6.680 2.460 ;
        RECT  5.280 1.580 5.680 1.820 ;
        RECT  3.840 1.290 4.080 3.200 ;
        RECT  0.960 1.020 1.200 3.190 ;
        RECT  3.700 1.020 3.940 1.530 ;
        RECT  0.160 1.020 3.940 1.260 ;
        RECT  3.120 1.580 3.360 4.340 ;
        RECT  3.120 2.260 3.550 2.660 ;
        RECT  3.040 1.580 3.440 1.820 ;
        RECT  1.530 3.930 1.930 4.170 ;
        RECT  1.690 3.540 1.930 4.170 ;
        RECT  1.690 3.540 2.800 3.780 ;
        RECT  2.560 1.580 2.800 3.780 ;
        RECT  2.560 2.260 2.870 2.660 ;
        RECT  1.600 1.580 2.800 1.820 ;
    END
END DFFRBT

MACRO DFFRSBN
    CLASS CORE ;
    FOREIGN DFFRSBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 2.140 9.750 3.210 ;
        RECT  9.080 2.140 9.750 2.540 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.690 2.840 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 1.300 14.090 3.840 ;
        RECT  13.780 3.440 14.090 3.840 ;
        RECT  13.780 1.300 14.090 1.700 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 1.300 12.850 3.400 ;
        RECT  12.550 3.000 12.850 3.400 ;
        RECT  12.550 1.300 12.850 1.700 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.480 1.620 8.720 2.450 ;
        RECT  6.780 2.210 8.720 2.450 ;
        RECT  9.480 1.100 9.720 1.860 ;
        RECT  8.480 1.620 9.720 1.860 ;
        RECT  9.480 1.100 10.990 1.340 ;
        RECT  10.710 1.100 10.990 2.210 ;
        RECT  6.780 2.140 7.020 2.540 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  8.360 -0.380 8.760 0.560 ;
        RECT  11.750 -0.380 12.150 0.860 ;
        RECT  12.980 -0.380 13.380 0.860 ;
        RECT  0.000 -0.380 14.260 0.380 ;
        RECT  1.040 -0.380 2.990 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.720 4.480 2.120 5.420 ;
        RECT  2.870 4.480 3.270 5.420 ;
        RECT  8.790 4.480 9.190 5.420 ;
        RECT  11.510 4.130 11.910 5.420 ;
        RECT  12.980 4.260 13.380 5.420 ;
        RECT  0.000 4.660 14.260 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.870 4.180 5.310 4.420 ;
        RECT  5.070 3.580 5.310 4.420 ;
        RECT  3.870 0.620 4.110 4.420 ;
        RECT  3.790 3.620 4.110 4.020 ;
        RECT  12.070 3.690 13.530 3.930 ;
        RECT  13.290 2.140 13.530 3.930 ;
        RECT  7.810 3.580 10.230 3.820 ;
        RECT  9.990 2.940 10.230 3.820 ;
        RECT  5.070 3.580 6.680 3.820 ;
        RECT  12.070 1.100 12.310 3.930 ;
        RECT  6.440 3.360 8.050 3.600 ;
        RECT  9.990 2.940 12.310 3.180 ;
        RECT  11.270 1.100 12.310 1.340 ;
        RECT  11.270 0.620 11.510 1.340 ;
        RECT  10.470 0.620 11.510 0.860 ;
        RECT  3.710 0.620 4.110 0.860 ;
        RECT  10.110 2.450 11.830 2.690 ;
        RECT  11.590 2.140 11.830 2.690 ;
        RECT  10.110 1.580 10.350 2.690 ;
        RECT  9.960 1.580 10.360 1.820 ;
        RECT  9.720 4.090 10.710 4.330 ;
        RECT  10.470 3.540 10.710 4.330 ;
        RECT  10.470 3.540 11.730 3.780 ;
        RECT  4.350 3.700 4.830 3.940 ;
        RECT  4.350 1.100 4.590 3.940 ;
        RECT  6.240 1.120 9.240 1.360 ;
        RECT  9.000 0.620 9.240 1.360 ;
        RECT  4.350 1.100 6.480 1.340 ;
        RECT  4.720 0.860 5.120 1.340 ;
        RECT  9.000 0.620 10.090 0.860 ;
        RECT  8.440 2.820 8.680 3.220 ;
        RECT  5.550 2.880 8.680 3.120 ;
        RECT  6.300 1.600 6.540 3.120 ;
        RECT  5.550 1.600 8.040 1.840 ;
        RECT  5.550 1.580 5.950 1.840 ;
        RECT  5.600 4.160 8.530 4.400 ;
        RECT  7.050 3.840 7.450 4.400 ;
        RECT  7.720 0.620 8.120 0.880 ;
        RECT  5.590 0.620 8.120 0.860 ;
        RECT  4.830 2.880 5.230 3.120 ;
        RECT  4.910 1.580 5.150 3.120 ;
        RECT  5.820 2.140 6.060 2.540 ;
        RECT  4.910 2.220 6.060 2.460 ;
        RECT  4.830 1.580 5.230 1.820 ;
        RECT  0.930 3.440 1.200 3.840 ;
        RECT  0.930 1.010 1.170 3.840 ;
        RECT  3.390 1.290 3.630 3.200 ;
        RECT  3.250 1.010 3.490 1.530 ;
        RECT  0.160 1.010 3.490 1.250 ;
        RECT  2.670 3.620 3.190 4.040 ;
        RECT  2.670 1.580 2.910 4.040 ;
        RECT  2.670 2.260 3.100 2.660 ;
        RECT  2.590 1.580 2.990 1.820 ;
        RECT  1.720 3.540 2.320 3.780 ;
        RECT  2.080 1.580 2.320 3.780 ;
        RECT  2.080 2.260 2.390 2.660 ;
        RECT  1.720 1.580 2.320 1.820 ;
    END
END DFFRSBN

MACRO DFFS
    CLASS CORE ;
    FOREIGN DFFS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.970 2.230 2.310 2.630 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.710 0.830 10.990 3.200 ;
        RECT  10.680 2.800 10.990 3.200 ;
        RECT  10.680 0.830 10.990 1.230 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.660 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.360 0.620 9.640 1.540 ;
        RECT  9.470 1.260 9.750 3.200 ;
        RECT  9.240 2.800 9.750 3.200 ;
        RECT  9.240 0.620 9.640 1.020 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.310 -0.380 2.710 0.560 ;
        RECT  7.890 -0.380 8.130 0.640 ;
        RECT  9.880 -0.380 10.280 0.940 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.910 -0.380 1.310 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 4.040 2.780 5.420 ;
        RECT  5.970 4.480 6.370 5.420 ;
        RECT  7.680 4.480 8.080 5.420 ;
        RECT  9.950 4.130 10.350 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.190 4.260 0.590 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.650 4.100 9.050 4.340 ;
        RECT  8.730 1.370 8.970 4.340 ;
        RECT  8.730 3.440 10.420 3.680 ;
        RECT  10.180 2.160 10.420 3.680 ;
        RECT  7.890 2.480 8.970 2.720 ;
        RECT  7.360 0.890 8.820 1.130 ;
        RECT  8.420 0.730 8.820 1.130 ;
        RECT  4.800 0.620 5.040 1.020 ;
        RECT  7.360 0.620 7.600 1.130 ;
        RECT  4.800 0.620 7.600 0.860 ;
        RECT  4.720 4.000 8.380 4.240 ;
        RECT  8.140 3.080 8.380 4.240 ;
        RECT  4.000 3.520 4.240 4.160 ;
        RECT  4.000 3.520 7.780 3.760 ;
        RECT  7.410 1.660 7.650 3.760 ;
        RECT  4.320 0.620 4.560 3.760 ;
        RECT  7.350 1.660 7.650 2.060 ;
        RECT  3.810 0.620 4.560 0.860 ;
        RECT  5.790 3.040 7.110 3.280 ;
        RECT  6.870 1.100 7.110 3.280 ;
        RECT  5.790 2.120 6.030 3.280 ;
        RECT  5.630 2.120 6.030 2.360 ;
        RECT  6.560 1.100 7.110 1.340 ;
        RECT  4.800 1.500 5.040 3.200 ;
        RECT  6.290 2.260 6.630 2.660 ;
        RECT  6.290 1.580 6.530 2.660 ;
        RECT  4.800 1.580 6.530 1.820 ;
        RECT  0.940 3.240 1.230 3.640 ;
        RECT  0.940 1.100 1.180 3.640 ;
        RECT  3.840 1.100 4.080 3.200 ;
        RECT  0.190 1.100 4.080 1.340 ;
        RECT  3.180 1.580 3.420 4.360 ;
        RECT  3.040 1.580 3.440 1.820 ;
        RECT  1.660 4.040 2.130 4.280 ;
        RECT  1.890 3.560 2.130 4.280 ;
        RECT  1.890 3.560 2.930 3.800 ;
        RECT  2.550 3.400 2.930 3.800 ;
        RECT  2.550 1.580 2.790 3.800 ;
        RECT  1.660 1.580 2.790 1.820 ;
    END
END DFFS

MACRO DFFSBN
    CLASS CORE ;
    FOREIGN DFFSBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.690 2.840 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 1.490 12.850 3.190 ;
        RECT  12.540 2.790 12.850 3.190 ;
        RECT  12.540 1.490 12.850 1.890 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.100 1.490 11.640 1.890 ;
        RECT  11.100 2.790 11.640 3.190 ;
        RECT  11.330 1.490 11.610 3.190 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.230 8.610 2.630 ;
        RECT  8.230 2.120 8.510 2.840 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  8.440 -0.380 8.840 0.560 ;
        RECT  9.620 -0.380 10.020 0.560 ;
        RECT  11.740 -0.380 12.140 0.950 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  1.040 -0.380 2.990 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.720 4.480 2.120 5.420 ;
        RECT  2.870 4.480 3.270 5.420 ;
        RECT  6.730 4.480 7.130 5.420 ;
        RECT  8.240 3.840 8.640 5.420 ;
        RECT  9.600 4.480 10.000 5.420 ;
        RECT  11.740 4.260 12.140 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.870 4.180 5.310 4.420 ;
        RECT  5.070 3.360 5.310 4.420 ;
        RECT  9.830 4.000 11.380 4.240 ;
        RECT  3.870 0.620 4.110 4.420 ;
        RECT  12.040 2.230 12.280 4.020 ;
        RECT  3.790 3.620 4.110 4.020 ;
        RECT  11.140 3.780 12.280 4.020 ;
        RECT  9.830 3.360 10.070 4.240 ;
        RECT  5.070 3.360 10.070 3.600 ;
        RECT  8.940 1.650 9.180 3.600 ;
        RECT  8.940 1.650 9.810 1.890 ;
        RECT  9.570 1.490 9.810 1.890 ;
        RECT  3.710 0.620 4.110 0.860 ;
        RECT  10.390 3.520 10.790 3.760 ;
        RECT  10.480 2.190 10.720 3.760 ;
        RECT  9.450 2.190 11.040 2.430 ;
        RECT  10.590 0.680 10.830 2.430 ;
        RECT  4.350 3.700 4.830 3.940 ;
        RECT  4.350 1.100 4.590 3.940 ;
        RECT  10.050 1.410 10.350 1.810 ;
        RECT  6.420 1.380 8.070 1.620 ;
        RECT  7.830 0.800 8.070 1.620 ;
        RECT  10.050 0.800 10.290 1.810 ;
        RECT  6.420 1.100 6.660 1.620 ;
        RECT  4.350 1.100 6.660 1.340 ;
        RECT  4.530 0.760 4.930 1.340 ;
        RECT  7.830 0.800 10.290 1.040 ;
        RECT  5.550 3.840 5.790 4.420 ;
        RECT  6.130 3.840 6.530 4.240 ;
        RECT  5.550 3.840 7.920 4.080 ;
        RECT  5.760 2.880 7.730 3.120 ;
        RECT  7.490 1.860 7.730 3.120 ;
        RECT  5.870 1.860 7.730 2.100 ;
        RECT  5.870 1.580 6.110 2.100 ;
        RECT  5.550 1.580 6.110 1.820 ;
        RECT  7.080 0.900 7.590 1.140 ;
        RECT  7.080 0.620 7.320 1.140 ;
        RECT  5.330 0.620 7.320 0.860 ;
        RECT  4.830 2.880 5.230 3.120 ;
        RECT  4.910 1.580 5.150 3.120 ;
        RECT  4.910 2.340 7.250 2.580 ;
        RECT  4.830 1.580 5.230 1.820 ;
        RECT  0.930 3.440 1.200 3.840 ;
        RECT  0.930 1.010 1.170 3.840 ;
        RECT  3.390 1.290 3.630 3.200 ;
        RECT  3.250 1.010 3.490 1.530 ;
        RECT  0.160 1.010 3.490 1.250 ;
        RECT  2.670 3.620 3.190 4.040 ;
        RECT  2.670 1.580 2.910 4.040 ;
        RECT  2.670 2.260 3.100 2.660 ;
        RECT  2.590 1.580 2.990 1.820 ;
        RECT  1.720 3.540 2.320 3.780 ;
        RECT  2.080 1.580 2.320 3.780 ;
        RECT  2.080 2.260 2.390 2.660 ;
        RECT  1.720 1.580 2.320 1.820 ;
    END
END DFFSBN

MACRO DFTRBN
    CLASS CORE ;
    FOREIGN DFTRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN QZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.520 2.790 14.090 3.190 ;
        RECT  13.810 1.320 14.090 3.430 ;
        RECT  13.520 1.320 14.090 1.720 ;
        END
    END QZ
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.880 2.280 8.120 2.680 ;
        RECT  7.610 1.930 7.890 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.230 1.800 2.630 ;
        RECT  1.410 2.120 1.690 2.840 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.670 1.890 15.950 2.750 ;
        RECT  15.540 2.020 15.950 2.420 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.140 1.080 2.540 ;
        RECT  0.790 2.120 1.070 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.770 1.510 11.610 1.820 ;
        RECT  11.330 1.510 11.610 3.400 ;
        RECT  10.850 3.000 11.610 3.400 ;
        RECT  10.770 1.480 11.170 1.820 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  7.760 -0.380 8.160 0.560 ;
        RECT  9.980 -0.380 10.380 0.860 ;
        RECT  12.000 -0.380 12.400 0.780 ;
        RECT  15.560 -0.380 15.960 1.480 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  1.100 -0.380 3.090 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.890 4.480 2.290 5.420 ;
        RECT  2.980 4.480 3.380 5.420 ;
        RECT  7.590 4.480 7.990 5.420 ;
        RECT  9.620 4.130 10.020 5.420 ;
        RECT  12.000 4.260 12.400 5.420 ;
        RECT  15.560 3.690 15.960 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  0.880 4.100 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  14.920 1.160 15.160 3.450 ;
        RECT  14.730 2.510 15.160 2.910 ;
        RECT  11.440 1.030 13.120 1.270 ;
        RECT  14.160 0.650 14.560 1.080 ;
        RECT  12.880 0.840 14.560 1.080 ;
        RECT  11.440 0.620 11.680 1.270 ;
        RECT  11.280 0.620 11.680 0.860 ;
        RECT  11.280 4.180 11.680 4.420 ;
        RECT  11.440 3.780 11.680 4.420 ;
        RECT  11.440 3.780 14.560 4.020 ;
        RECT  3.970 4.180 5.460 4.420 ;
        RECT  5.220 3.580 5.460 4.420 ;
        RECT  3.970 0.620 4.210 4.420 ;
        RECT  3.890 3.620 4.210 4.020 ;
        RECT  5.220 3.580 8.510 3.820 ;
        RECT  8.270 2.880 8.510 3.820 ;
        RECT  8.270 2.880 10.470 3.120 ;
        RECT  10.230 1.100 10.470 3.120 ;
        RECT  9.420 1.100 10.470 1.340 ;
        RECT  9.420 0.620 9.660 1.340 ;
        RECT  9.260 0.620 9.660 0.860 ;
        RECT  3.810 0.620 4.210 0.860 ;
        RECT  9.750 1.640 9.990 2.540 ;
        RECT  9.170 1.640 9.990 1.880 ;
        RECT  9.170 1.580 9.570 1.880 ;
        RECT  8.520 4.090 9.040 4.330 ;
        RECT  8.800 3.420 9.040 4.330 ;
        RECT  8.800 3.420 9.970 3.660 ;
        RECT  4.450 3.700 4.980 3.940 ;
        RECT  4.450 1.100 4.690 3.940 ;
        RECT  8.490 2.120 9.340 2.360 ;
        RECT  8.490 1.120 8.730 2.360 ;
        RECT  6.340 1.120 8.730 1.360 ;
        RECT  4.450 1.100 6.580 1.340 ;
        RECT  4.700 0.860 5.100 1.340 ;
        RECT  5.650 2.980 7.560 3.220 ;
        RECT  7.130 1.600 7.370 3.220 ;
        RECT  5.650 2.880 6.050 3.220 ;
        RECT  5.650 1.600 7.370 1.840 ;
        RECT  5.650 1.580 6.050 1.840 ;
        RECT  7.090 0.620 7.490 0.880 ;
        RECT  5.690 0.620 7.490 0.860 ;
        RECT  5.700 4.160 7.330 4.400 ;
        RECT  4.930 2.880 5.330 3.120 ;
        RECT  5.010 1.580 5.250 3.120 ;
        RECT  5.010 2.220 6.330 2.460 ;
        RECT  4.930 1.580 5.330 1.820 ;
        RECT  3.490 1.100 3.730 3.200 ;
        RECT  0.190 2.800 0.480 3.200 ;
        RECT  0.190 1.010 0.430 3.200 ;
        RECT  3.060 1.100 3.730 1.340 ;
        RECT  0.160 1.010 3.300 1.250 ;
        RECT  2.770 3.540 3.300 3.940 ;
        RECT  2.770 1.580 3.010 3.940 ;
        RECT  2.770 2.480 3.190 2.880 ;
        RECT  2.690 1.580 3.090 1.820 ;
        RECT  1.780 3.620 2.450 3.860 ;
        RECT  2.210 1.580 2.450 3.860 ;
        RECT  2.210 2.970 2.510 3.370 ;
        RECT  1.910 1.580 2.450 1.820 ;
    END
END DFTRBN

MACRO DFTRBS
    CLASS CORE ;
    FOREIGN DFTRBS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN QZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 0.620 12.780 1.020 ;
        RECT  11.950 4.020 12.790 4.420 ;
        RECT  11.950 0.620 12.230 4.420 ;
        END
    END QZ
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.880 2.280 8.120 2.680 ;
        RECT  7.610 1.930 7.890 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.230 1.800 2.630 ;
        RECT  1.410 2.120 1.690 2.840 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 1.880 14.090 2.750 ;
        RECT  13.680 1.880 14.090 2.280 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.140 1.080 2.540 ;
        RECT  0.790 2.120 1.070 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 1.300 11.610 3.400 ;
        RECT  10.850 3.000 11.610 3.400 ;
        RECT  10.850 1.300 11.610 1.700 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  7.760 -0.380 8.160 0.560 ;
        RECT  9.980 -0.380 10.380 0.860 ;
        RECT  11.280 -0.380 11.680 0.780 ;
        RECT  13.700 -0.380 14.100 1.500 ;
        RECT  0.000 -0.380 14.260 0.380 ;
        RECT  1.100 -0.380 3.090 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.890 4.480 2.290 5.420 ;
        RECT  2.980 4.480 3.380 5.420 ;
        RECT  7.590 4.480 7.990 5.420 ;
        RECT  9.620 4.130 10.020 5.420 ;
        RECT  11.280 4.260 11.680 5.420 ;
        RECT  13.700 3.690 14.100 5.420 ;
        RECT  0.000 4.660 14.260 5.420 ;
        RECT  0.880 4.100 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.060 1.340 13.300 3.450 ;
        RECT  12.870 2.510 13.300 2.910 ;
        RECT  3.970 4.180 5.460 4.420 ;
        RECT  5.220 3.580 5.460 4.420 ;
        RECT  3.970 0.620 4.210 4.420 ;
        RECT  3.890 3.620 4.210 4.020 ;
        RECT  5.220 3.580 8.510 3.820 ;
        RECT  8.270 2.880 8.510 3.820 ;
        RECT  8.270 2.880 10.470 3.120 ;
        RECT  10.230 1.100 10.470 3.120 ;
        RECT  9.420 1.100 10.470 1.340 ;
        RECT  9.420 0.620 9.660 1.340 ;
        RECT  9.260 0.620 9.660 0.860 ;
        RECT  3.810 0.620 4.210 0.860 ;
        RECT  9.750 1.640 9.990 2.540 ;
        RECT  9.170 1.640 9.990 1.880 ;
        RECT  9.170 1.580 9.570 1.880 ;
        RECT  8.520 4.090 9.040 4.330 ;
        RECT  8.800 3.420 9.040 4.330 ;
        RECT  8.800 3.420 9.970 3.660 ;
        RECT  4.450 3.700 4.980 3.940 ;
        RECT  4.450 1.100 4.690 3.940 ;
        RECT  8.490 2.120 9.340 2.360 ;
        RECT  8.490 1.120 8.730 2.360 ;
        RECT  6.340 1.120 8.730 1.360 ;
        RECT  4.450 1.100 6.580 1.340 ;
        RECT  4.700 0.860 5.100 1.340 ;
        RECT  5.650 2.980 7.560 3.220 ;
        RECT  7.130 1.600 7.370 3.220 ;
        RECT  5.650 2.880 6.050 3.220 ;
        RECT  5.650 1.600 7.370 1.840 ;
        RECT  5.650 1.580 6.050 1.840 ;
        RECT  7.090 0.620 7.490 0.880 ;
        RECT  5.690 0.620 7.490 0.860 ;
        RECT  5.700 4.160 7.330 4.400 ;
        RECT  4.930 2.880 5.330 3.120 ;
        RECT  5.010 1.580 5.250 3.120 ;
        RECT  5.010 2.220 6.330 2.460 ;
        RECT  4.930 1.580 5.330 1.820 ;
        RECT  3.490 1.100 3.730 3.200 ;
        RECT  0.190 2.800 0.480 3.200 ;
        RECT  0.190 1.010 0.430 3.200 ;
        RECT  3.060 1.100 3.730 1.340 ;
        RECT  0.160 1.010 3.300 1.250 ;
        RECT  2.770 3.540 3.300 3.940 ;
        RECT  2.770 1.580 3.010 3.940 ;
        RECT  2.770 2.480 3.190 2.880 ;
        RECT  2.690 1.580 3.090 1.820 ;
        RECT  1.780 3.620 2.450 3.860 ;
        RECT  2.210 1.580 2.450 3.860 ;
        RECT  2.210 2.970 2.510 3.370 ;
        RECT  1.910 1.580 2.450 1.820 ;
    END
END DFTRBS

MACRO DFZCLRBN
    CLASS CORE ;
    FOREIGN DFZCLRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.940 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.330 2.500 ;
        RECT  2.030 2.100 2.310 3.160 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.230 11.850 2.630 ;
        RECT  11.330 2.120 11.610 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 1.590 10.370 2.550 ;
        RECT  9.970 1.860 10.370 2.260 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  22.490 1.260 22.770 3.220 ;
        RECT  22.280 2.940 22.770 3.220 ;
        RECT  22.280 1.260 22.770 1.540 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.060 3.690 2.460 ;
        RECT  3.270 2.060 3.550 2.710 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  20.570 1.280 20.970 3.200 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.030 3.520 10.970 3.760 ;
        RECT  10.730 2.030 11.070 2.430 ;
        RECT  10.730 2.030 10.970 3.760 ;
        END
    END SEL
    PIN LD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.430 1.620 1.670 2.630 ;
        RECT  1.430 1.620 3.010 1.860 ;
        RECT  2.770 1.620 3.010 3.430 ;
        RECT  4.190 2.280 4.430 3.430 ;
        RECT  2.770 3.190 4.430 3.430 ;
        RECT  1.410 2.140 1.670 2.540 ;
        END
    END LD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.780 ;
        RECT  6.500 -0.380 6.900 0.780 ;
        RECT  9.360 -0.380 9.760 0.780 ;
        RECT  11.960 -0.380 12.360 0.560 ;
        RECT  16.110 -0.380 16.510 0.860 ;
        RECT  19.020 -0.380 19.420 0.560 ;
        RECT  21.290 -0.380 21.960 0.800 ;
        RECT  0.000 -0.380 22.940 0.380 ;
        RECT  0.290 -0.380 0.530 1.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.470 4.200 2.870 5.420 ;
        RECT  5.060 4.260 5.460 5.420 ;
        RECT  6.560 4.480 7.600 5.420 ;
        RECT  10.260 4.480 10.660 5.420 ;
        RECT  11.960 4.480 12.360 5.420 ;
        RECT  16.110 4.200 16.510 5.420 ;
        RECT  19.170 4.400 19.410 5.420 ;
        RECT  21.560 4.260 21.960 5.420 ;
        RECT  0.000 4.660 22.940 5.420 ;
        RECT  0.290 2.790 0.530 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  17.330 4.180 18.930 4.420 ;
        RECT  18.690 3.720 18.930 4.420 ;
        RECT  13.040 4.180 15.330 4.420 ;
        RECT  15.090 3.720 15.330 4.420 ;
        RECT  5.700 4.000 13.280 4.240 ;
        RECT  17.330 3.720 17.570 4.420 ;
        RECT  13.970 0.620 14.210 4.420 ;
        RECT  5.700 3.700 5.940 4.240 ;
        RECT  18.690 3.720 21.840 3.960 ;
        RECT  21.600 2.160 21.840 3.960 ;
        RECT  15.090 3.720 17.570 3.960 ;
        RECT  13.520 3.700 14.210 3.940 ;
        RECT  5.170 3.700 5.940 3.940 ;
        RECT  19.600 1.320 19.840 3.960 ;
        RECT  5.170 2.250 5.410 3.940 ;
        RECT  19.600 2.980 19.890 3.380 ;
        RECT  19.600 1.320 19.890 1.720 ;
        RECT  13.460 0.620 14.210 0.860 ;
        RECT  18.210 3.200 18.450 3.940 ;
        RECT  18.210 3.200 19.340 3.440 ;
        RECT  19.100 0.890 19.340 3.440 ;
        RECT  19.100 2.160 19.360 2.560 ;
        RECT  18.210 0.890 19.340 1.130 ;
        RECT  18.210 0.730 18.450 1.130 ;
        RECT  14.450 3.700 14.850 3.940 ;
        RECT  14.450 0.620 14.690 3.940 ;
        RECT  17.700 1.100 17.940 3.200 ;
        RECT  17.700 2.210 18.520 2.450 ;
        RECT  15.480 1.100 17.940 1.340 ;
        RECT  15.480 0.620 15.720 1.340 ;
        RECT  14.450 0.620 15.720 0.860 ;
        RECT  15.880 2.880 17.460 3.120 ;
        RECT  17.220 1.580 17.460 3.120 ;
        RECT  15.880 2.260 16.120 3.120 ;
        RECT  16.900 1.580 17.460 1.820 ;
        RECT  14.930 1.500 15.170 3.200 ;
        RECT  16.420 2.170 16.900 2.570 ;
        RECT  16.420 1.730 16.660 2.570 ;
        RECT  14.930 1.730 16.660 1.970 ;
        RECT  8.700 3.030 9.730 3.270 ;
        RECT  9.490 1.100 9.730 3.270 ;
        RECT  13.490 1.100 13.730 3.200 ;
        RECT  8.880 1.100 13.730 1.340 ;
        RECT  10.800 0.860 11.200 1.340 ;
        RECT  8.880 0.620 9.120 1.340 ;
        RECT  8.120 0.620 9.120 0.860 ;
        RECT  12.750 3.520 13.150 3.760 ;
        RECT  12.830 1.580 13.070 3.760 ;
        RECT  12.830 2.300 13.190 2.700 ;
        RECT  12.690 1.580 13.090 1.820 ;
        RECT  11.310 3.520 12.440 3.760 ;
        RECT  12.200 1.580 12.440 3.760 ;
        RECT  12.200 2.900 12.540 3.300 ;
        RECT  11.310 1.580 12.440 1.820 ;
        RECT  6.880 2.440 7.120 3.190 ;
        RECT  6.880 2.440 9.250 2.680 ;
        RECT  9.010 2.240 9.250 2.680 ;
        RECT  7.150 1.570 7.550 2.680 ;
        RECT  5.650 2.790 5.890 3.190 ;
        RECT  5.650 2.790 6.640 3.030 ;
        RECT  6.400 1.090 6.640 3.030 ;
        RECT  7.790 1.940 8.630 2.180 ;
        RECT  7.790 1.090 8.030 2.180 ;
        RECT  5.860 1.090 8.030 1.330 ;
        RECT  5.860 0.930 6.100 1.330 ;
        RECT  1.590 3.720 1.990 4.080 ;
        RECT  1.590 3.720 4.930 3.960 ;
        RECT  4.690 1.100 4.930 3.960 ;
        RECT  5.920 1.770 6.160 2.260 ;
        RECT  5.310 1.770 6.160 2.010 ;
        RECT  5.310 1.100 5.550 2.010 ;
        RECT  3.800 1.100 5.550 1.340 ;
        RECT  2.320 0.620 5.460 0.860 ;
        RECT  0.810 3.730 1.150 4.130 ;
        RECT  0.810 1.140 1.050 4.130 ;
        RECT  0.810 2.790 1.250 3.190 ;
        RECT  4.190 1.580 4.430 1.980 ;
        RECT  3.320 1.580 4.430 1.820 ;
        RECT  3.320 1.140 3.560 1.820 ;
        RECT  0.810 1.140 3.560 1.380 ;
    END
END DFZCLRBN

MACRO DFZCRBN
    CLASS CORE ;
    FOREIGN DFZCRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.580 4.170 2.560 ;
        RECT  3.750 1.860 4.170 2.260 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 2.230 5.490 2.630 ;
        RECT  5.130 2.120 5.410 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.460 2.410 2.860 ;
        RECT  2.030 2.360 2.310 3.230 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.020 2.880 15.330 3.280 ;
        RECT  15.050 1.250 15.330 3.400 ;
        RECT  15.020 1.350 15.330 1.750 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.580 4.790 2.560 ;
        RECT  4.460 1.860 4.790 2.260 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 1.260 14.090 3.190 ;
        RECT  13.580 2.790 14.090 3.190 ;
        RECT  13.580 0.770 13.860 1.540 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.410 0.480 2.810 ;
        RECT  0.170 2.210 0.450 2.950 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.490 -0.380 2.890 0.840 ;
        RECT  5.440 -0.380 5.840 0.560 ;
        RECT  6.220 -0.380 6.620 0.600 ;
        RECT  9.560 -0.380 9.960 0.860 ;
        RECT  12.370 -0.380 12.770 0.560 ;
        RECT  14.300 -0.380 14.620 1.030 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.440 -0.380 0.840 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.270 4.200 2.670 5.420 ;
        RECT  5.810 4.180 6.210 5.420 ;
        RECT  9.560 4.200 9.960 5.420 ;
        RECT  12.620 4.400 12.860 5.420 ;
        RECT  14.220 4.260 14.620 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.440 4.210 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.780 4.180 12.380 4.420 ;
        RECT  12.140 3.720 12.380 4.420 ;
        RECT  7.520 4.180 8.880 4.420 ;
        RECT  8.640 3.720 8.880 4.420 ;
        RECT  10.780 3.720 11.020 4.420 ;
        RECT  7.520 0.620 7.760 4.420 ;
        RECT  12.140 3.720 14.730 3.960 ;
        RECT  14.490 2.160 14.730 3.960 ;
        RECT  8.640 3.720 11.020 3.960 ;
        RECT  7.280 3.700 7.760 3.940 ;
        RECT  13.050 3.530 13.310 3.960 ;
        RECT  13.050 1.490 13.290 3.960 ;
        RECT  13.050 1.490 13.310 1.890 ;
        RECT  7.010 0.620 7.760 0.860 ;
        RECT  11.660 3.200 11.900 3.940 ;
        RECT  11.660 3.200 12.810 3.440 ;
        RECT  12.570 0.890 12.810 3.440 ;
        RECT  11.660 0.890 12.810 1.130 ;
        RECT  11.660 0.730 11.900 1.130 ;
        RECT  8.000 3.700 8.400 3.940 ;
        RECT  8.000 0.620 8.240 3.940 ;
        RECT  11.150 1.100 11.390 3.200 ;
        RECT  11.150 2.210 11.970 2.450 ;
        RECT  9.030 1.100 11.390 1.340 ;
        RECT  9.030 0.620 9.270 1.340 ;
        RECT  8.000 0.620 9.270 0.860 ;
        RECT  9.390 2.880 10.910 3.120 ;
        RECT  10.670 1.580 10.910 3.120 ;
        RECT  9.390 2.260 9.630 3.120 ;
        RECT  10.350 1.580 10.910 1.820 ;
        RECT  8.480 1.500 8.720 3.200 ;
        RECT  9.870 2.170 10.350 2.570 ;
        RECT  9.870 1.730 10.110 2.570 ;
        RECT  8.480 1.730 10.110 1.970 ;
        RECT  1.280 3.700 1.680 4.080 ;
        RECT  1.280 3.700 4.260 3.940 ;
        RECT  3.270 0.800 3.510 3.940 ;
        RECT  7.040 1.100 7.280 3.200 ;
        RECT  1.210 1.080 1.610 1.640 ;
        RECT  5.620 1.100 7.280 1.340 ;
        RECT  1.210 1.080 3.510 1.320 ;
        RECT  5.620 0.800 5.860 1.340 ;
        RECT  3.270 0.800 5.860 1.040 ;
        RECT  6.530 4.180 6.930 4.420 ;
        RECT  6.560 1.580 6.800 4.420 ;
        RECT  6.500 2.460 6.800 2.860 ;
        RECT  6.220 1.580 6.800 1.820 ;
        RECT  5.090 4.180 5.490 4.420 ;
        RECT  5.250 3.700 5.490 4.420 ;
        RECT  5.250 3.700 6.320 3.940 ;
        RECT  5.730 3.420 6.320 3.940 ;
        RECT  5.730 1.580 5.970 3.940 ;
        RECT  5.440 1.580 5.970 1.820 ;
        RECT  3.090 4.180 4.850 4.420 ;
        RECT  4.610 2.960 4.850 4.420 ;
        RECT  4.610 2.960 4.900 3.360 ;
        RECT  0.520 3.190 0.960 3.590 ;
        RECT  0.720 1.320 0.960 3.590 ;
        RECT  0.720 2.260 1.670 2.660 ;
        RECT  1.430 1.880 1.670 2.660 ;
        RECT  2.790 1.860 3.030 2.260 ;
        RECT  1.430 1.880 3.030 2.120 ;
        RECT  0.520 1.320 0.960 1.720 ;
    END
END DFZCRBN

MACRO DFZN
    CLASS CORE ;
    FOREIGN DFZN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        RECT  3.830 2.230 4.170 2.630 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.220 2.310 2.620 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 1.480 12.850 3.200 ;
        RECT  12.540 2.800 12.850 3.200 ;
        RECT  12.540 1.480 12.850 1.880 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.220 0.620 11.500 1.540 ;
        RECT  11.330 1.260 11.610 3.200 ;
        RECT  11.100 2.800 11.610 3.200 ;
        RECT  11.100 0.620 11.500 1.020 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.170 -0.380 4.570 0.560 ;
        RECT  9.750 -0.380 9.990 0.640 ;
        RECT  11.740 -0.380 12.140 0.940 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.240 4.040 4.640 5.420 ;
        RECT  7.830 4.480 8.230 5.420 ;
        RECT  9.540 4.480 9.940 5.420 ;
        RECT  11.740 4.260 12.140 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  2.010 4.480 2.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.510 3.850 10.910 4.090 ;
        RECT  12.040 2.160 12.280 4.020 ;
        RECT  10.590 3.780 12.280 4.020 ;
        RECT  10.590 1.370 10.830 4.090 ;
        RECT  9.750 2.480 10.830 2.720 ;
        RECT  9.220 0.890 10.680 1.130 ;
        RECT  10.280 0.730 10.680 1.130 ;
        RECT  6.660 0.620 6.900 1.020 ;
        RECT  9.220 0.620 9.460 1.130 ;
        RECT  6.660 0.620 9.460 0.860 ;
        RECT  6.580 4.000 10.240 4.240 ;
        RECT  10.000 3.080 10.240 4.240 ;
        RECT  5.860 3.520 6.100 4.160 ;
        RECT  5.860 3.520 9.640 3.760 ;
        RECT  9.270 1.660 9.510 3.760 ;
        RECT  6.180 0.620 6.420 3.760 ;
        RECT  9.210 1.660 9.510 2.060 ;
        RECT  5.670 0.620 6.420 0.860 ;
        RECT  7.650 3.040 8.970 3.280 ;
        RECT  8.730 1.100 8.970 3.280 ;
        RECT  7.650 2.120 7.890 3.280 ;
        RECT  7.490 2.120 7.890 2.360 ;
        RECT  8.420 1.100 8.970 1.340 ;
        RECT  6.660 1.500 6.900 3.200 ;
        RECT  8.150 2.260 8.490 2.660 ;
        RECT  8.150 1.580 8.390 2.660 ;
        RECT  6.660 1.580 8.390 1.820 ;
        RECT  5.700 1.100 5.940 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.040 1.580 5.280 4.360 ;
        RECT  4.900 1.580 5.300 1.820 ;
        RECT  3.520 4.040 3.990 4.280 ;
        RECT  3.750 3.560 3.990 4.280 ;
        RECT  3.750 3.560 4.790 3.800 ;
        RECT  4.410 3.400 4.790 3.800 ;
        RECT  4.410 1.580 4.650 3.800 ;
        RECT  3.520 1.580 4.650 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.180 0.990 4.420 ;
        RECT  0.750 3.460 0.990 4.420 ;
        RECT  0.750 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END DFZN

MACRO DFZP
    CLASS CORE ;
    FOREIGN DFZP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        RECT  3.830 2.230 4.170 2.630 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.220 2.310 2.620 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.050 1.240 15.330 3.220 ;
        RECT  14.220 2.940 15.330 3.220 ;
        RECT  14.220 1.240 15.330 1.520 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.510 1.260 13.180 1.500 ;
        RECT  12.510 2.960 13.180 3.200 ;
        RECT  12.510 1.260 12.910 3.200 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.170 -0.380 4.570 0.560 ;
        RECT  8.220 -0.380 8.620 0.860 ;
        RECT  12.060 -0.380 12.460 0.780 ;
        RECT  13.500 -0.380 13.900 0.780 ;
        RECT  14.940 -0.380 15.340 0.780 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.240 4.020 4.640 5.420 ;
        RECT  8.220 4.200 8.620 5.420 ;
        RECT  12.060 4.260 12.460 5.420 ;
        RECT  13.500 4.260 13.900 5.420 ;
        RECT  14.940 4.260 15.340 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  2.010 4.480 2.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.440 4.180 11.040 4.420 ;
        RECT  10.800 3.720 11.040 4.420 ;
        RECT  6.180 4.180 7.540 4.420 ;
        RECT  7.300 3.720 7.540 4.420 ;
        RECT  9.440 3.720 9.680 4.420 ;
        RECT  6.180 0.620 6.420 4.420 ;
        RECT  10.800 3.720 13.950 3.960 ;
        RECT  13.710 2.240 13.950 3.960 ;
        RECT  7.300 3.720 9.680 3.960 ;
        RECT  5.730 3.700 6.420 3.940 ;
        RECT  11.710 1.320 11.950 3.960 ;
        RECT  11.630 2.810 11.950 3.210 ;
        RECT  13.710 2.240 14.490 2.480 ;
        RECT  11.630 1.320 11.950 1.720 ;
        RECT  5.670 0.620 6.420 0.860 ;
        RECT  10.320 3.200 10.560 3.940 ;
        RECT  10.320 3.200 11.340 3.440 ;
        RECT  11.100 0.800 11.340 3.440 ;
        RECT  11.100 2.160 11.470 2.560 ;
        RECT  10.320 0.720 10.560 1.120 ;
        RECT  10.320 0.800 11.340 1.040 ;
        RECT  6.660 3.700 7.060 3.940 ;
        RECT  6.660 0.620 6.900 3.940 ;
        RECT  9.810 1.100 10.050 3.200 ;
        RECT  9.810 2.210 10.630 2.450 ;
        RECT  7.690 1.100 10.050 1.340 ;
        RECT  7.690 0.620 7.930 1.340 ;
        RECT  6.660 0.620 7.930 0.860 ;
        RECT  8.050 2.880 9.570 3.120 ;
        RECT  9.330 1.580 9.570 3.120 ;
        RECT  8.050 2.260 8.290 3.120 ;
        RECT  9.010 1.580 9.570 1.820 ;
        RECT  7.140 1.500 7.380 3.200 ;
        RECT  8.530 2.170 9.010 2.570 ;
        RECT  8.530 1.730 8.770 2.570 ;
        RECT  7.140 1.730 8.770 1.970 ;
        RECT  5.700 1.100 5.940 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.040 1.580 5.280 4.340 ;
        RECT  4.900 1.580 5.300 1.820 ;
        RECT  3.520 4.020 3.920 4.260 ;
        RECT  3.680 3.540 3.920 4.260 ;
        RECT  3.680 3.540 4.650 3.780 ;
        RECT  4.410 1.580 4.650 3.780 ;
        RECT  4.410 3.220 4.790 3.620 ;
        RECT  3.520 1.580 4.650 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.160 0.990 4.400 ;
        RECT  0.750 3.460 0.990 4.400 ;
        RECT  0.750 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END DFZP

MACRO DFZRBN
    CLASS CORE ;
    FOREIGN DFZRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.470 2.540 ;
        RECT  10.090 1.930 10.370 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.270 2.310 2.670 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 1.300 14.710 3.840 ;
        RECT  14.370 3.440 14.710 3.840 ;
        RECT  14.370 1.300 14.710 1.700 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.300 13.470 3.400 ;
        RECT  13.140 3.000 13.470 3.400 ;
        RECT  13.140 1.300 13.470 1.700 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.380 4.650 0.560 ;
        RECT  10.110 -0.380 10.510 0.560 ;
        RECT  12.340 -0.380 12.740 0.860 ;
        RECT  13.570 -0.380 13.970 0.860 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 4.030 4.720 5.420 ;
        RECT  9.940 4.480 10.340 5.420 ;
        RECT  11.970 4.130 12.370 5.420 ;
        RECT  13.570 4.260 13.970 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  2.090 4.480 2.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 4.180 7.760 4.420 ;
        RECT  7.520 3.580 7.760 4.420 ;
        RECT  6.320 0.620 6.560 4.420 ;
        RECT  6.240 3.620 6.560 4.020 ;
        RECT  12.580 3.720 14.120 3.960 ;
        RECT  13.880 2.140 14.120 3.960 ;
        RECT  7.520 3.580 10.860 3.820 ;
        RECT  10.620 2.880 10.860 3.820 ;
        RECT  12.580 1.100 12.820 3.960 ;
        RECT  10.620 2.880 12.820 3.120 ;
        RECT  11.780 1.100 12.820 1.340 ;
        RECT  11.780 0.620 12.020 1.340 ;
        RECT  11.620 0.620 12.020 0.860 ;
        RECT  6.160 0.620 6.560 0.860 ;
        RECT  12.100 1.640 12.340 2.540 ;
        RECT  11.520 1.640 12.340 1.880 ;
        RECT  11.520 1.580 11.920 1.880 ;
        RECT  10.870 4.090 11.390 4.330 ;
        RECT  11.150 3.540 11.390 4.330 ;
        RECT  11.150 3.540 12.320 3.780 ;
        RECT  6.800 3.700 7.280 3.940 ;
        RECT  6.800 1.100 7.040 3.940 ;
        RECT  10.840 2.120 11.690 2.360 ;
        RECT  10.840 1.120 11.080 2.360 ;
        RECT  8.690 1.120 11.080 1.360 ;
        RECT  6.800 1.100 8.930 1.340 ;
        RECT  7.170 0.860 7.570 1.340 ;
        RECT  9.440 0.620 9.840 0.880 ;
        RECT  8.040 0.620 9.840 0.860 ;
        RECT  9.590 1.600 9.830 3.220 ;
        RECT  8.000 2.880 9.830 3.120 ;
        RECT  8.000 1.600 9.830 1.840 ;
        RECT  8.000 1.580 8.400 1.840 ;
        RECT  8.050 4.160 9.680 4.400 ;
        RECT  7.280 2.880 7.680 3.120 ;
        RECT  7.360 1.580 7.600 3.120 ;
        RECT  7.360 2.220 8.680 2.460 ;
        RECT  7.280 1.580 7.680 1.820 ;
        RECT  5.840 1.290 6.080 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.700 1.290 6.080 1.530 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.120 1.580 5.360 4.350 ;
        RECT  5.120 2.260 5.550 2.660 ;
        RECT  5.040 1.580 5.440 1.820 ;
        RECT  3.600 4.030 4.000 4.270 ;
        RECT  3.760 3.540 4.000 4.270 ;
        RECT  3.760 3.540 4.800 3.780 ;
        RECT  4.560 1.580 4.800 3.780 ;
        RECT  4.560 2.260 4.870 2.660 ;
        RECT  3.600 1.580 4.800 1.820 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.280 3.700 ;
        RECT  2.880 3.940 3.280 4.420 ;
        RECT  1.230 3.940 3.280 4.180 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
    END
END DFZRBN

MACRO DFZRBP
    CLASS CORE ;
    FOREIGN DFZRBP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.470 2.540 ;
        RECT  10.090 1.930 10.370 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.270 2.310 2.670 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.050 1.280 15.330 3.260 ;
        RECT  14.920 2.860 15.330 3.260 ;
        RECT  14.920 1.280 15.330 1.680 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 1.260 14.090 3.220 ;
        RECT  13.400 2.940 14.090 3.220 ;
        RECT  13.400 1.260 14.090 1.540 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.380 4.650 0.560 ;
        RECT  10.040 -0.380 10.440 0.560 ;
        RECT  12.680 -0.380 13.080 0.860 ;
        RECT  14.120 -0.380 14.520 0.860 ;
        RECT  15.560 -0.380 15.960 0.860 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 4.020 4.720 5.420 ;
        RECT  9.940 4.480 10.340 5.420 ;
        RECT  11.660 4.480 12.060 5.420 ;
        RECT  12.470 4.480 12.870 5.420 ;
        RECT  14.120 4.260 14.520 5.420 ;
        RECT  15.560 4.260 15.960 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  2.090 4.480 2.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 4.180 7.760 4.420 ;
        RECT  7.520 3.580 7.760 4.420 ;
        RECT  6.320 0.620 6.560 4.420 ;
        RECT  6.240 3.620 6.560 4.020 ;
        RECT  7.520 3.580 14.590 3.820 ;
        RECT  14.350 2.140 14.590 3.820 ;
        RECT  12.920 1.100 13.160 3.820 ;
        RECT  14.350 2.140 14.750 2.540 ;
        RECT  12.120 1.100 13.160 1.340 ;
        RECT  12.120 0.620 12.360 1.340 ;
        RECT  11.960 0.620 12.360 0.860 ;
        RECT  6.160 0.620 6.560 0.860 ;
        RECT  10.870 3.100 12.680 3.340 ;
        RECT  12.440 1.640 12.680 3.340 ;
        RECT  11.450 1.640 12.680 1.880 ;
        RECT  11.450 1.570 11.850 1.880 ;
        RECT  6.800 3.700 7.280 3.940 ;
        RECT  6.800 1.100 7.040 3.940 ;
        RECT  10.840 2.220 11.690 2.460 ;
        RECT  10.840 1.120 11.080 2.460 ;
        RECT  8.690 1.120 11.080 1.360 ;
        RECT  6.800 1.100 8.930 1.340 ;
        RECT  7.170 0.860 7.570 1.340 ;
        RECT  9.590 1.600 9.830 3.220 ;
        RECT  8.000 2.880 9.830 3.120 ;
        RECT  8.000 1.600 9.830 1.840 ;
        RECT  8.000 1.580 8.400 1.840 ;
        RECT  9.370 0.620 9.770 0.880 ;
        RECT  8.040 0.620 9.770 0.860 ;
        RECT  8.050 4.160 9.680 4.400 ;
        RECT  7.280 2.880 7.680 3.120 ;
        RECT  7.360 1.580 7.600 3.120 ;
        RECT  7.360 2.220 8.680 2.460 ;
        RECT  7.280 1.580 7.680 1.820 ;
        RECT  5.840 1.290 6.080 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.700 1.290 6.080 1.530 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.120 1.580 5.360 4.340 ;
        RECT  5.120 2.260 5.550 2.660 ;
        RECT  5.040 1.580 5.440 1.820 ;
        RECT  3.600 4.020 4.000 4.260 ;
        RECT  3.760 3.540 4.000 4.260 ;
        RECT  3.760 3.540 4.800 3.780 ;
        RECT  4.560 1.580 4.800 3.780 ;
        RECT  4.560 2.260 4.870 2.660 ;
        RECT  3.600 1.580 4.800 1.820 ;
        RECT  0.160 4.140 0.990 4.380 ;
        RECT  0.750 3.460 0.990 4.380 ;
        RECT  0.750 3.460 3.280 3.700 ;
        RECT  2.880 3.940 3.280 4.420 ;
        RECT  1.230 3.940 3.280 4.180 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
    END
END DFZRBP

MACRO DFZRBS
    CLASS CORE ;
    FOREIGN DFZRBS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.470 2.540 ;
        RECT  10.090 1.930 10.370 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.270 2.310 2.670 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 0.650 14.710 4.100 ;
        RECT  14.370 3.700 14.710 4.100 ;
        RECT  14.370 0.650 14.710 1.050 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.150 2.790 13.470 3.190 ;
        RECT  13.190 1.400 13.470 3.190 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.380 4.650 0.560 ;
        RECT  10.110 -0.380 10.510 0.560 ;
        RECT  12.340 -0.380 12.740 0.860 ;
        RECT  13.570 -0.380 13.970 0.860 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 4.030 4.720 5.420 ;
        RECT  9.940 4.480 10.340 5.420 ;
        RECT  11.970 4.130 12.370 5.420 ;
        RECT  13.570 4.260 13.970 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  2.090 4.480 2.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 4.180 7.760 4.420 ;
        RECT  7.520 3.580 7.760 4.420 ;
        RECT  6.320 0.620 6.560 4.420 ;
        RECT  6.240 3.620 6.560 4.020 ;
        RECT  12.580 3.720 14.120 3.960 ;
        RECT  13.880 2.140 14.120 3.960 ;
        RECT  7.520 3.580 10.860 3.820 ;
        RECT  10.620 2.880 10.860 3.820 ;
        RECT  12.580 1.100 12.820 3.960 ;
        RECT  10.620 2.880 12.820 3.120 ;
        RECT  11.780 1.100 12.820 1.340 ;
        RECT  11.780 0.620 12.020 1.340 ;
        RECT  11.620 0.620 12.020 0.860 ;
        RECT  6.160 0.620 6.560 0.860 ;
        RECT  12.100 1.640 12.340 2.540 ;
        RECT  11.520 1.640 12.340 1.880 ;
        RECT  11.520 1.580 11.920 1.880 ;
        RECT  10.870 4.090 11.390 4.330 ;
        RECT  11.150 3.580 11.390 4.330 ;
        RECT  11.150 3.580 12.320 3.820 ;
        RECT  6.800 3.700 7.280 3.940 ;
        RECT  6.800 1.100 7.040 3.940 ;
        RECT  10.840 2.120 11.690 2.360 ;
        RECT  10.840 1.120 11.080 2.360 ;
        RECT  8.690 1.120 11.080 1.360 ;
        RECT  6.800 1.100 8.930 1.340 ;
        RECT  7.170 0.860 7.570 1.340 ;
        RECT  9.440 0.620 9.840 0.880 ;
        RECT  8.040 0.620 9.840 0.860 ;
        RECT  9.590 1.600 9.830 3.220 ;
        RECT  8.000 2.880 9.830 3.120 ;
        RECT  8.000 1.600 9.830 1.840 ;
        RECT  8.000 1.580 8.400 1.840 ;
        RECT  8.050 4.160 9.680 4.400 ;
        RECT  7.280 2.880 7.680 3.120 ;
        RECT  7.360 1.580 7.600 3.120 ;
        RECT  7.360 2.220 8.680 2.460 ;
        RECT  7.280 1.580 7.680 1.820 ;
        RECT  5.840 1.290 6.080 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.700 1.290 6.080 1.530 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.120 1.580 5.360 4.350 ;
        RECT  5.120 2.260 5.550 2.660 ;
        RECT  5.040 1.580 5.440 1.820 ;
        RECT  3.600 4.030 4.000 4.270 ;
        RECT  3.760 3.540 4.000 4.270 ;
        RECT  3.760 3.540 4.800 3.780 ;
        RECT  4.560 1.580 4.800 3.780 ;
        RECT  4.560 2.260 4.870 2.660 ;
        RECT  3.600 1.580 4.800 1.820 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.280 3.700 ;
        RECT  2.880 3.940 3.280 4.420 ;
        RECT  1.230 3.940 3.280 4.180 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
    END
END DFZRBS

MACRO DFZRBT
    CLASS CORE ;
    FOREIGN DFZRBT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.980 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.390 2.540 ;
        RECT  10.090 1.930 10.370 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        RECT  3.830 2.230 4.170 2.630 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.250 2.310 2.650 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 1.200 16.570 3.710 ;
        RECT  16.060 3.310 16.570 3.710 ;
        RECT  17.500 1.200 17.810 1.600 ;
        RECT  16.290 2.320 17.810 2.720 ;
        RECT  17.530 1.200 17.810 3.710 ;
        RECT  17.500 3.310 17.810 3.710 ;
        RECT  16.060 1.200 16.570 1.600 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.390 2.820 13.630 3.220 ;
        RECT  13.390 1.260 15.150 1.540 ;
        RECT  14.370 1.260 14.770 3.220 ;
        RECT  14.370 1.260 15.150 1.580 ;
        RECT  13.390 2.940 15.150 3.220 ;
        RECT  13.390 1.260 13.630 1.660 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.170 -0.380 4.570 0.560 ;
        RECT  10.010 -0.380 10.410 0.560 ;
        RECT  12.590 -0.380 12.990 0.860 ;
        RECT  14.030 -0.380 14.430 0.860 ;
        RECT  15.260 -0.380 15.660 0.860 ;
        RECT  16.700 -0.380 17.100 0.860 ;
        RECT  0.000 -0.380 17.980 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.240 4.020 4.640 5.420 ;
        RECT  9.990 4.480 10.390 5.420 ;
        RECT  11.570 4.480 11.970 5.420 ;
        RECT  12.390 4.480 12.790 5.420 ;
        RECT  14.030 4.260 14.430 5.420 ;
        RECT  15.260 4.260 15.660 5.420 ;
        RECT  16.700 4.260 17.100 5.420 ;
        RECT  0.000 4.660 17.980 5.420 ;
        RECT  2.010 4.480 2.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.240 4.180 7.680 4.420 ;
        RECT  7.440 3.580 7.680 4.420 ;
        RECT  6.240 0.620 6.480 4.420 ;
        RECT  6.160 3.620 6.480 4.020 ;
        RECT  7.440 3.580 15.810 3.820 ;
        RECT  15.570 2.140 15.810 3.820 ;
        RECT  12.910 1.100 13.150 3.820 ;
        RECT  12.030 1.100 13.150 1.340 ;
        RECT  12.030 0.620 12.270 1.340 ;
        RECT  11.870 0.620 12.270 0.860 ;
        RECT  6.080 0.620 6.480 0.860 ;
        RECT  10.780 3.100 12.670 3.340 ;
        RECT  12.430 1.640 12.670 3.340 ;
        RECT  11.360 1.640 12.670 1.880 ;
        RECT  11.360 1.570 11.760 1.880 ;
        RECT  6.720 3.700 7.200 3.940 ;
        RECT  6.720 1.100 6.960 3.940 ;
        RECT  10.760 2.220 11.610 2.460 ;
        RECT  10.760 1.120 11.000 2.460 ;
        RECT  8.610 1.120 11.000 1.360 ;
        RECT  6.720 1.100 8.850 1.340 ;
        RECT  7.090 0.860 7.490 1.340 ;
        RECT  9.510 2.820 9.750 3.220 ;
        RECT  7.920 2.880 9.750 3.120 ;
        RECT  9.430 1.600 9.670 3.120 ;
        RECT  7.920 1.600 9.670 1.840 ;
        RECT  7.920 1.580 8.320 1.840 ;
        RECT  9.270 0.620 9.670 0.880 ;
        RECT  7.960 0.620 9.670 0.860 ;
        RECT  7.970 4.160 9.600 4.400 ;
        RECT  7.200 2.880 7.600 3.120 ;
        RECT  7.280 1.580 7.520 3.120 ;
        RECT  7.280 2.220 8.600 2.460 ;
        RECT  7.200 1.580 7.600 1.820 ;
        RECT  5.760 1.290 6.000 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.620 1.290 6.000 1.530 ;
        RECT  2.970 1.100 5.860 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.040 1.580 5.280 4.340 ;
        RECT  5.040 2.260 5.470 2.660 ;
        RECT  4.960 1.580 5.360 1.820 ;
        RECT  3.520 4.020 3.920 4.260 ;
        RECT  3.680 3.540 3.920 4.260 ;
        RECT  3.680 3.540 4.720 3.780 ;
        RECT  4.480 1.580 4.720 3.780 ;
        RECT  4.480 2.260 4.790 2.660 ;
        RECT  3.520 1.580 4.720 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END DFZRBT

MACRO DFZRSBN
    CLASS CORE ;
    FOREIGN DFZRSBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.010 2.140 11.680 2.540 ;
        RECT  11.330 2.140 11.610 3.210 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.170 3.590 2.570 ;
        RECT  3.270 2.120 3.550 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.250 2.310 2.650 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.670 0.650 15.950 4.100 ;
        RECT  15.640 3.700 15.950 4.100 ;
        RECT  15.640 0.650 15.950 1.050 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 1.400 14.710 3.190 ;
        RECT  14.410 2.790 14.710 3.190 ;
        RECT  14.410 1.400 14.710 1.800 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.410 1.620 10.650 2.450 ;
        RECT  8.680 2.210 10.650 2.450 ;
        RECT  11.410 1.100 11.650 1.860 ;
        RECT  10.410 1.620 11.650 1.860 ;
        RECT  11.410 1.100 12.850 1.340 ;
        RECT  12.570 1.100 12.850 2.210 ;
        RECT  12.570 1.540 12.900 1.940 ;
        RECT  8.680 2.140 8.920 2.540 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.640 -0.380 4.040 0.560 ;
        RECT  4.480 -0.380 4.880 0.560 ;
        RECT  10.290 -0.380 10.690 0.560 ;
        RECT  13.610 -0.380 14.010 0.860 ;
        RECT  14.840 -0.380 15.240 0.950 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.640 4.480 4.040 5.420 ;
        RECT  4.760 4.480 5.160 5.420 ;
        RECT  10.720 4.480 11.120 5.420 ;
        RECT  13.100 4.130 13.500 5.420 ;
        RECT  14.840 4.260 15.240 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  2.010 4.480 2.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.770 4.180 7.210 4.420 ;
        RECT  6.970 3.580 7.210 4.420 ;
        RECT  5.770 0.620 6.010 4.420 ;
        RECT  5.690 3.620 6.010 4.020 ;
        RECT  9.740 3.580 12.160 3.820 ;
        RECT  11.920 2.940 12.160 3.820 ;
        RECT  6.970 3.580 8.610 3.820 ;
        RECT  13.930 3.430 15.260 3.670 ;
        RECT  15.020 2.140 15.260 3.670 ;
        RECT  8.370 3.360 9.980 3.600 ;
        RECT  13.930 1.100 14.170 3.670 ;
        RECT  11.920 2.940 14.170 3.180 ;
        RECT  15.020 2.140 15.430 2.540 ;
        RECT  13.090 1.100 14.170 1.340 ;
        RECT  13.090 0.620 13.330 1.340 ;
        RECT  12.400 0.620 13.330 0.860 ;
        RECT  5.610 0.620 6.010 0.860 ;
        RECT  12.040 2.450 13.690 2.690 ;
        RECT  13.450 2.140 13.690 2.690 ;
        RECT  12.040 1.580 12.280 2.690 ;
        RECT  11.890 1.580 12.290 1.820 ;
        RECT  11.650 4.090 12.640 4.330 ;
        RECT  12.400 3.540 12.640 4.330 ;
        RECT  12.400 3.540 13.660 3.780 ;
        RECT  6.250 3.700 6.730 3.940 ;
        RECT  6.250 1.100 6.490 3.940 ;
        RECT  8.140 1.120 11.170 1.360 ;
        RECT  10.930 0.620 11.170 1.360 ;
        RECT  6.250 1.100 8.380 1.340 ;
        RECT  6.620 0.860 7.020 1.340 ;
        RECT  10.930 0.620 12.020 0.860 ;
        RECT  10.370 2.820 10.610 3.220 ;
        RECT  7.450 2.880 10.610 3.120 ;
        RECT  8.200 1.600 8.440 3.120 ;
        RECT  7.450 1.600 9.970 1.840 ;
        RECT  7.450 1.580 7.850 1.840 ;
        RECT  7.500 4.160 10.460 4.400 ;
        RECT  8.980 3.840 9.380 4.400 ;
        RECT  9.650 0.620 10.050 0.880 ;
        RECT  7.490 0.620 10.050 0.860 ;
        RECT  6.730 2.880 7.130 3.120 ;
        RECT  6.810 1.580 7.050 3.120 ;
        RECT  7.720 2.140 7.960 2.540 ;
        RECT  6.810 2.220 7.960 2.460 ;
        RECT  6.730 1.580 7.130 1.820 ;
        RECT  5.230 2.800 5.530 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  5.230 1.290 5.470 3.200 ;
        RECT  5.230 1.500 5.530 1.900 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.120 1.100 5.360 1.530 ;
        RECT  2.970 1.100 5.360 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  4.560 3.620 5.080 4.040 ;
        RECT  4.560 1.580 4.800 4.040 ;
        RECT  4.560 2.260 4.990 2.660 ;
        RECT  4.480 1.580 4.880 1.820 ;
        RECT  3.640 3.350 4.240 3.590 ;
        RECT  4.000 1.580 4.240 3.590 ;
        RECT  4.000 2.260 4.310 2.660 ;
        RECT  3.640 1.580 4.240 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.150 0.980 4.390 ;
        RECT  0.740 3.460 0.980 4.390 ;
        RECT  0.740 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END DFZRSBN

MACRO DFZS
    CLASS CORE ;
    FOREIGN DFZS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        RECT  3.830 2.230 4.170 2.630 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.220 2.310 2.620 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 0.830 12.850 3.200 ;
        RECT  12.540 2.800 12.850 3.200 ;
        RECT  12.540 0.830 12.850 1.230 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.220 0.620 11.500 1.540 ;
        RECT  11.330 1.260 11.610 3.200 ;
        RECT  11.100 2.800 11.610 3.200 ;
        RECT  11.100 0.620 11.500 1.020 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.170 -0.380 4.570 0.560 ;
        RECT  9.720 -0.380 10.120 0.560 ;
        RECT  11.740 -0.380 12.140 0.940 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.240 4.040 4.640 5.420 ;
        RECT  7.830 4.480 8.230 5.420 ;
        RECT  9.540 4.480 9.940 5.420 ;
        RECT  11.670 4.130 12.070 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  2.010 4.480 2.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.510 4.180 10.910 4.420 ;
        RECT  10.590 1.410 10.830 4.420 ;
        RECT  10.590 3.440 12.280 3.680 ;
        RECT  12.040 2.160 12.280 3.680 ;
        RECT  9.750 2.480 10.830 2.720 ;
        RECT  10.510 1.420 10.910 1.660 ;
        RECT  9.220 0.930 10.680 1.170 ;
        RECT  10.280 0.830 10.680 1.170 ;
        RECT  6.660 0.620 6.900 1.020 ;
        RECT  9.220 0.620 9.460 1.170 ;
        RECT  6.660 0.620 9.460 0.860 ;
        RECT  6.580 4.000 10.240 4.240 ;
        RECT  10.000 3.080 10.240 4.240 ;
        RECT  5.860 3.520 6.100 4.160 ;
        RECT  5.860 3.520 9.640 3.760 ;
        RECT  9.270 1.660 9.510 3.760 ;
        RECT  6.180 0.620 6.420 3.760 ;
        RECT  9.210 1.660 9.510 2.060 ;
        RECT  5.670 0.620 6.420 0.860 ;
        RECT  7.650 3.040 8.970 3.280 ;
        RECT  8.730 1.100 8.970 3.280 ;
        RECT  7.650 2.120 7.890 3.280 ;
        RECT  7.490 2.120 7.890 2.360 ;
        RECT  8.420 1.100 8.970 1.340 ;
        RECT  6.660 1.500 6.900 3.200 ;
        RECT  8.150 2.260 8.490 2.660 ;
        RECT  8.150 1.580 8.390 2.660 ;
        RECT  6.660 1.580 8.390 1.820 ;
        RECT  5.700 1.100 5.940 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.040 1.580 5.280 4.360 ;
        RECT  4.900 1.580 5.300 1.820 ;
        RECT  3.520 4.040 3.990 4.280 ;
        RECT  3.750 3.560 3.990 4.280 ;
        RECT  3.750 3.560 4.790 3.800 ;
        RECT  4.410 3.400 4.790 3.800 ;
        RECT  4.410 1.580 4.650 3.800 ;
        RECT  3.520 1.580 4.650 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.180 0.990 4.420 ;
        RECT  0.750 3.460 0.990 4.420 ;
        RECT  0.750 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END DFZS

MACRO DFZSBN
    CLASS CORE ;
    FOREIGN DFZSBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.170 3.590 2.570 ;
        RECT  3.270 2.120 3.550 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.250 2.310 2.650 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 1.490 14.710 3.190 ;
        RECT  14.400 2.790 14.710 3.190 ;
        RECT  14.400 1.490 14.710 1.890 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.490 13.470 3.190 ;
        RECT  12.960 2.790 13.470 3.190 ;
        RECT  12.960 1.490 13.470 1.890 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.230 10.470 2.630 ;
        RECT  10.090 2.120 10.370 2.840 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.640 -0.380 4.040 0.560 ;
        RECT  4.480 -0.380 4.880 0.560 ;
        RECT  10.300 -0.380 10.700 0.560 ;
        RECT  11.480 -0.380 11.880 0.560 ;
        RECT  13.600 -0.380 14.000 0.950 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.640 4.480 4.040 5.420 ;
        RECT  4.760 4.480 5.160 5.420 ;
        RECT  8.590 4.480 8.990 5.420 ;
        RECT  10.100 3.840 10.500 5.420 ;
        RECT  11.460 4.480 11.860 5.420 ;
        RECT  13.600 4.260 14.000 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  2.010 4.480 2.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.760 4.180 7.200 4.420 ;
        RECT  6.960 3.360 7.200 4.420 ;
        RECT  11.770 4.000 13.240 4.240 ;
        RECT  5.760 0.620 6.000 4.420 ;
        RECT  13.890 2.230 14.130 4.020 ;
        RECT  5.680 3.620 6.000 4.020 ;
        RECT  13.000 3.780 14.130 4.020 ;
        RECT  11.770 3.360 12.010 4.240 ;
        RECT  6.960 3.360 12.010 3.600 ;
        RECT  10.800 1.650 11.040 3.600 ;
        RECT  10.800 1.650 11.670 1.890 ;
        RECT  11.430 1.490 11.670 1.890 ;
        RECT  5.600 0.620 6.000 0.860 ;
        RECT  12.250 3.520 12.650 3.760 ;
        RECT  12.340 2.190 12.580 3.760 ;
        RECT  11.310 2.190 12.860 2.430 ;
        RECT  12.450 0.680 12.690 2.430 ;
        RECT  6.240 3.700 6.720 3.940 ;
        RECT  6.240 1.100 6.480 3.940 ;
        RECT  11.910 1.410 12.210 1.810 ;
        RECT  8.280 1.380 9.930 1.620 ;
        RECT  9.690 0.800 9.930 1.620 ;
        RECT  11.910 0.800 12.150 1.810 ;
        RECT  8.280 1.100 8.520 1.620 ;
        RECT  6.240 1.100 8.520 1.340 ;
        RECT  6.420 0.760 6.820 1.340 ;
        RECT  9.690 0.800 12.150 1.040 ;
        RECT  7.440 3.840 7.680 4.420 ;
        RECT  7.990 3.840 8.390 4.240 ;
        RECT  7.440 3.840 9.780 4.080 ;
        RECT  7.650 2.880 9.590 3.120 ;
        RECT  9.350 1.860 9.590 3.120 ;
        RECT  7.730 1.860 9.590 2.100 ;
        RECT  7.730 1.580 7.970 2.100 ;
        RECT  7.440 1.580 7.970 1.820 ;
        RECT  8.940 0.900 9.450 1.140 ;
        RECT  8.940 0.620 9.180 1.140 ;
        RECT  7.220 0.620 9.180 0.860 ;
        RECT  6.720 2.880 7.120 3.120 ;
        RECT  6.800 1.580 7.040 3.120 ;
        RECT  6.800 2.340 9.110 2.580 ;
        RECT  6.720 1.580 7.120 1.820 ;
        RECT  5.230 2.800 5.520 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  5.230 1.290 5.470 3.200 ;
        RECT  5.230 1.500 5.520 1.900 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.120 1.100 5.360 1.530 ;
        RECT  2.970 1.100 5.360 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  4.560 3.620 5.080 4.040 ;
        RECT  4.560 1.580 4.800 4.040 ;
        RECT  4.560 2.260 4.990 2.660 ;
        RECT  4.480 1.580 4.880 1.820 ;
        RECT  3.640 3.350 4.240 3.590 ;
        RECT  4.000 1.580 4.240 3.590 ;
        RECT  4.000 2.260 4.310 2.660 ;
        RECT  3.640 1.580 4.240 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.150 0.980 4.390 ;
        RECT  0.740 3.460 0.980 4.390 ;
        RECT  0.740 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END DFZSBN

MACRO DFZTRBN
    CLASS CORE ;
    FOREIGN DFZTRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.980 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN QZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.670 1.320 15.950 3.190 ;
        RECT  15.380 2.790 15.950 3.190 ;
        RECT  15.380 1.320 15.950 1.720 ;
        END
    END QZ
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.740 2.280 9.980 2.680 ;
        RECT  9.470 1.930 9.750 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.230 3.660 2.630 ;
        RECT  3.270 2.120 3.550 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.230 2.310 2.630 ;
        END
    END TD
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.530 1.890 17.810 2.750 ;
        RECT  17.400 2.020 17.810 2.420 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.510 13.470 3.400 ;
        RECT  12.710 3.000 13.470 3.400 ;
        RECT  12.630 1.510 13.470 1.750 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.770 -0.380 4.170 0.560 ;
        RECT  4.550 -0.380 4.950 0.560 ;
        RECT  9.620 -0.380 10.020 0.560 ;
        RECT  11.840 -0.380 12.240 0.860 ;
        RECT  13.860 -0.380 14.260 0.780 ;
        RECT  17.420 -0.380 17.820 1.480 ;
        RECT  0.000 -0.380 17.980 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.640 4.480 4.040 5.420 ;
        RECT  4.840 4.480 5.240 5.420 ;
        RECT  9.450 4.480 9.850 5.420 ;
        RECT  11.480 4.260 11.880 5.420 ;
        RECT  13.860 4.260 14.260 5.420 ;
        RECT  17.420 3.690 17.820 5.420 ;
        RECT  0.000 4.660 17.980 5.420 ;
        RECT  1.930 4.480 2.330 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  16.780 1.160 17.020 3.450 ;
        RECT  16.590 2.510 17.020 2.910 ;
        RECT  14.580 1.020 14.980 1.270 ;
        RECT  14.740 0.620 14.980 1.270 ;
        RECT  13.300 1.020 14.980 1.260 ;
        RECT  13.300 0.620 13.540 1.260 ;
        RECT  14.740 0.620 16.420 0.860 ;
        RECT  13.140 0.620 13.540 0.860 ;
        RECT  15.500 4.180 16.420 4.420 ;
        RECT  13.140 4.180 13.540 4.420 ;
        RECT  13.300 3.780 13.540 4.420 ;
        RECT  15.500 3.780 15.740 4.420 ;
        RECT  13.300 3.780 15.740 4.020 ;
        RECT  5.830 4.180 7.270 4.420 ;
        RECT  7.030 3.580 7.270 4.420 ;
        RECT  5.830 0.620 6.070 4.420 ;
        RECT  5.750 3.620 6.070 4.020 ;
        RECT  7.030 3.580 10.370 3.820 ;
        RECT  10.130 2.880 10.370 3.820 ;
        RECT  10.130 2.880 12.330 3.120 ;
        RECT  12.090 1.100 12.330 3.120 ;
        RECT  11.280 1.100 12.330 1.340 ;
        RECT  11.280 0.620 11.520 1.340 ;
        RECT  11.120 0.620 11.520 0.860 ;
        RECT  5.670 0.620 6.070 0.860 ;
        RECT  11.610 1.640 11.850 2.540 ;
        RECT  11.030 1.640 11.850 1.880 ;
        RECT  11.030 1.580 11.430 1.880 ;
        RECT  10.380 4.090 10.900 4.330 ;
        RECT  10.660 3.420 10.900 4.330 ;
        RECT  10.660 3.420 11.830 3.660 ;
        RECT  6.310 3.700 6.790 3.940 ;
        RECT  6.310 1.100 6.550 3.940 ;
        RECT  10.350 2.120 11.200 2.360 ;
        RECT  10.350 1.120 10.590 2.360 ;
        RECT  8.200 1.120 10.590 1.360 ;
        RECT  6.310 1.100 8.440 1.340 ;
        RECT  6.560 0.860 6.960 1.340 ;
        RECT  7.510 2.980 9.420 3.220 ;
        RECT  8.990 1.600 9.230 3.220 ;
        RECT  7.510 2.880 7.910 3.220 ;
        RECT  7.510 1.600 9.230 1.840 ;
        RECT  7.510 1.580 7.910 1.840 ;
        RECT  8.950 0.620 9.350 0.880 ;
        RECT  7.550 0.620 9.350 0.860 ;
        RECT  7.560 4.160 9.190 4.400 ;
        RECT  6.790 2.880 7.190 3.120 ;
        RECT  6.870 1.580 7.110 3.120 ;
        RECT  6.870 2.220 8.190 2.460 ;
        RECT  6.790 1.580 7.190 1.820 ;
        RECT  5.350 1.290 5.590 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.210 1.290 5.590 1.530 ;
        RECT  2.970 1.100 5.450 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  4.630 3.540 5.160 3.940 ;
        RECT  4.630 1.580 4.870 3.940 ;
        RECT  4.630 2.480 5.050 2.880 ;
        RECT  4.550 1.580 4.950 1.820 ;
        RECT  3.640 3.620 4.310 3.860 ;
        RECT  4.070 1.580 4.310 3.860 ;
        RECT  4.070 2.970 4.370 3.370 ;
        RECT  3.770 1.580 4.310 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END DFZTRBN

MACRO DFZTRBS
    CLASS CORE ;
    FOREIGN DFZTRBS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN QZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 0.620 14.640 1.020 ;
        RECT  13.810 4.020 14.650 4.420 ;
        RECT  13.810 0.620 14.090 4.420 ;
        END
    END QZ
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.740 2.280 9.980 2.680 ;
        RECT  9.470 1.930 9.750 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.230 3.660 2.630 ;
        RECT  3.270 2.120 3.550 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.230 2.310 2.630 ;
        END
    END TD
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.670 1.880 15.950 2.750 ;
        RECT  15.540 1.880 15.950 2.280 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.300 13.470 3.400 ;
        RECT  12.710 3.000 13.470 3.400 ;
        RECT  12.710 1.300 13.470 1.700 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.770 -0.380 4.170 0.560 ;
        RECT  4.550 -0.380 4.950 0.560 ;
        RECT  9.620 -0.380 10.020 0.560 ;
        RECT  11.840 -0.380 12.240 0.860 ;
        RECT  13.140 -0.380 13.540 0.780 ;
        RECT  15.560 -0.380 15.960 1.500 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.640 4.480 4.040 5.420 ;
        RECT  4.840 4.480 5.240 5.420 ;
        RECT  9.450 4.480 9.850 5.420 ;
        RECT  11.480 4.130 11.880 5.420 ;
        RECT  13.140 4.260 13.540 5.420 ;
        RECT  15.560 3.690 15.960 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  1.930 4.480 2.330 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  14.920 1.340 15.160 3.450 ;
        RECT  14.730 2.510 15.160 2.910 ;
        RECT  5.830 4.180 7.270 4.420 ;
        RECT  7.030 3.580 7.270 4.420 ;
        RECT  5.830 0.620 6.070 4.420 ;
        RECT  5.750 3.620 6.070 4.020 ;
        RECT  7.030 3.580 10.370 3.820 ;
        RECT  10.130 2.880 10.370 3.820 ;
        RECT  10.130 2.880 12.330 3.120 ;
        RECT  12.090 1.100 12.330 3.120 ;
        RECT  11.280 1.100 12.330 1.340 ;
        RECT  11.280 0.620 11.520 1.340 ;
        RECT  11.120 0.620 11.520 0.860 ;
        RECT  5.670 0.620 6.070 0.860 ;
        RECT  11.610 1.640 11.850 2.540 ;
        RECT  11.030 1.640 11.850 1.880 ;
        RECT  11.030 1.580 11.430 1.880 ;
        RECT  10.380 4.090 10.900 4.330 ;
        RECT  10.660 3.420 10.900 4.330 ;
        RECT  10.660 3.420 11.830 3.660 ;
        RECT  6.310 3.700 6.790 3.940 ;
        RECT  6.310 1.100 6.550 3.940 ;
        RECT  10.350 2.120 11.200 2.360 ;
        RECT  10.350 1.120 10.590 2.360 ;
        RECT  8.200 1.120 10.590 1.360 ;
        RECT  6.310 1.100 8.440 1.340 ;
        RECT  6.560 0.860 6.960 1.340 ;
        RECT  7.510 2.980 9.420 3.220 ;
        RECT  8.990 1.600 9.230 3.220 ;
        RECT  7.510 2.880 7.910 3.220 ;
        RECT  7.510 1.600 9.230 1.840 ;
        RECT  7.510 1.580 7.910 1.840 ;
        RECT  8.950 0.620 9.350 0.880 ;
        RECT  7.550 0.620 9.350 0.860 ;
        RECT  7.560 4.160 9.190 4.400 ;
        RECT  6.790 2.880 7.190 3.120 ;
        RECT  6.870 1.580 7.110 3.120 ;
        RECT  6.870 2.220 8.190 2.460 ;
        RECT  6.790 1.580 7.190 1.820 ;
        RECT  5.350 1.290 5.590 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.210 1.290 5.590 1.530 ;
        RECT  2.970 1.100 5.450 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  4.630 3.540 5.160 3.940 ;
        RECT  4.630 1.580 4.870 3.940 ;
        RECT  4.630 2.480 5.050 2.880 ;
        RECT  4.550 1.580 4.950 1.820 ;
        RECT  3.640 3.620 4.310 3.860 ;
        RECT  4.070 1.580 4.310 3.860 ;
        RECT  4.070 2.970 4.370 3.370 ;
        RECT  3.770 1.580 4.310 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END DFZTRBS

MACRO DLHN
    CLASS CORE ;
    FOREIGN DLHN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.230 1.800 2.630 ;
        RECT  1.410 1.820 1.690 2.770 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.230 8.510 3.200 ;
        RECT  8.200 2.800 8.510 3.200 ;
        RECT  8.200 1.230 8.510 1.630 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.680 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.880 0.620 7.160 1.540 ;
        RECT  6.990 1.260 7.270 3.190 ;
        RECT  6.760 2.790 7.270 3.190 ;
        RECT  6.760 0.620 7.160 1.020 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.580 -0.380 2.980 0.560 ;
        RECT  5.960 -0.380 6.360 0.560 ;
        RECT  7.400 -0.380 7.800 0.940 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  1.040 -0.380 1.440 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.110 3.910 2.510 5.420 ;
        RECT  5.380 4.480 5.780 5.420 ;
        RECT  7.400 4.260 7.800 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.160 3.240 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.280 3.780 7.940 4.020 ;
        RECT  7.700 2.160 7.940 4.020 ;
        RECT  6.170 3.590 6.570 3.830 ;
        RECT  6.280 1.420 6.520 4.020 ;
        RECT  5.440 2.420 6.520 2.660 ;
        RECT  5.440 2.260 5.680 2.660 ;
        RECT  6.170 1.420 6.570 1.660 ;
        RECT  4.010 3.680 4.320 4.080 ;
        RECT  4.080 0.790 4.320 4.080 ;
        RECT  4.050 2.860 4.320 3.260 ;
        RECT  4.080 1.560 4.390 1.960 ;
        RECT  5.940 0.800 6.340 1.100 ;
        RECT  4.000 0.800 6.340 1.040 ;
        RECT  4.000 0.790 4.400 1.040 ;
        RECT  4.830 2.860 5.110 3.260 ;
        RECT  4.830 1.570 5.070 3.260 ;
        RECT  4.790 1.570 5.190 1.810 ;
        RECT  0.920 3.060 1.200 3.460 ;
        RECT  3.330 2.860 3.580 3.260 ;
        RECT  3.340 0.800 3.580 3.260 ;
        RECT  0.920 0.800 1.160 3.460 ;
        RECT  3.340 1.560 3.670 1.960 ;
        RECT  0.240 0.800 0.480 1.730 ;
        RECT  0.240 0.800 3.580 1.040 ;
        RECT  2.850 3.830 3.150 4.230 ;
        RECT  2.850 1.520 3.090 4.230 ;
        RECT  2.850 2.190 3.100 2.590 ;
        RECT  2.660 1.520 3.090 1.920 ;
        RECT  1.380 3.910 1.780 4.150 ;
        RECT  1.540 3.270 1.780 4.150 ;
        RECT  1.540 3.270 2.610 3.510 ;
        RECT  2.060 3.110 2.610 3.510 ;
        RECT  2.060 1.340 2.300 3.510 ;
        RECT  1.660 1.340 2.300 1.580 ;
    END
END DLHN

MACRO DLHP
    CLASS CORE ;
    FOREIGN DLHP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.300 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.410 0.450 2.500 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.490 8.510 3.190 ;
        RECT  8.100 2.790 8.510 3.190 ;
        RECT  8.100 1.490 8.510 1.890 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.010 2.200 2.540 2.600 ;
        RECT  2.010 1.840 2.290 2.870 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.440 1.570 7.270 1.810 ;
        RECT  6.520 2.790 7.270 3.190 ;
        RECT  6.970 1.570 7.250 3.190 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.040 -0.380 2.440 0.560 ;
        RECT  5.260 -0.380 5.660 0.560 ;
        RECT  7.230 -0.380 7.630 0.850 ;
        RECT  8.740 -0.380 9.140 1.030 ;
        RECT  0.000 -0.380 9.300 0.380 ;
        RECT  1.380 -0.380 1.780 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.110 4.470 2.510 5.420 ;
        RECT  5.520 4.480 5.920 5.420 ;
        RECT  7.300 4.250 7.700 5.420 ;
        RECT  8.740 4.250 9.140 5.420 ;
        RECT  0.000 4.660 9.300 5.420 ;
        RECT  0.950 4.470 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.220 1.090 5.460 3.480 ;
        RECT  7.610 1.090 7.850 2.500 ;
        RECT  5.030 2.100 5.460 2.500 ;
        RECT  5.220 1.090 7.850 1.330 ;
        RECT  3.530 4.180 5.270 4.420 ;
        RECT  5.970 2.100 6.210 4.230 ;
        RECT  5.030 3.990 6.210 4.230 ;
        RECT  3.530 1.390 3.770 4.420 ;
        RECT  5.970 2.100 6.330 2.500 ;
        RECT  4.300 3.700 4.790 3.940 ;
        RECT  4.550 0.620 4.790 3.940 ;
        RECT  4.070 0.800 4.310 3.190 ;
        RECT  1.320 0.800 1.560 3.190 ;
        RECT  1.320 0.800 4.310 1.040 ;
        RECT  2.960 0.710 3.360 1.040 ;
        RECT  0.160 3.990 3.290 4.230 ;
        RECT  0.780 0.670 1.020 4.230 ;
        RECT  0.780 3.430 1.800 3.670 ;
        RECT  0.300 0.670 1.020 0.910 ;
        RECT  2.810 1.390 3.050 3.190 ;
    END
END DLHP

MACRO DLHRBN
    CLASS CORE ;
    FOREIGN DLHRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.300 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.760 2.930 2.700 ;
        RECT  2.500 2.050 2.930 2.450 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.410 0.480 2.430 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.180 0.450 2.750 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.820 2.790 9.130 3.190 ;
        RECT  8.850 1.280 9.130 3.300 ;
        RECT  8.820 1.280 9.130 1.680 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.860 3.550 2.870 ;
        RECT  3.210 2.180 3.550 2.580 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.430 2.790 7.890 3.190 ;
        RECT  7.610 1.280 7.890 3.300 ;
        RECT  7.430 1.280 7.890 1.680 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.310 -0.380 6.710 0.560 ;
        RECT  8.000 -0.380 8.400 0.560 ;
        RECT  0.000 -0.380 9.300 0.380 ;
        RECT  1.260 -0.380 2.330 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 4.480 2.940 5.420 ;
        RECT  6.630 4.480 7.030 5.420 ;
        RECT  8.070 4.180 8.470 5.420 ;
        RECT  0.000 4.660 9.300 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.830 2.760 6.440 3.000 ;
        RECT  5.830 0.800 6.070 3.000 ;
        RECT  8.250 2.150 8.580 2.550 ;
        RECT  8.250 0.800 8.490 2.550 ;
        RECT  5.830 1.460 6.440 1.700 ;
        RECT  5.830 0.800 8.490 1.040 ;
        RECT  4.760 4.180 6.250 4.420 ;
        RECT  6.950 2.020 7.190 4.230 ;
        RECT  6.010 3.990 7.190 4.230 ;
        RECT  4.760 0.620 5.000 4.420 ;
        RECT  2.020 0.800 2.260 3.190 ;
        RECT  2.020 0.800 2.810 1.040 ;
        RECT  4.630 0.620 5.000 1.020 ;
        RECT  2.570 0.620 5.000 0.860 ;
        RECT  5.350 3.700 5.750 3.940 ;
        RECT  5.350 0.620 5.590 3.940 ;
        RECT  4.280 1.750 4.520 4.420 ;
        RECT  1.200 3.430 4.520 3.670 ;
        RECT  1.200 2.790 1.440 3.670 ;
        RECT  1.260 1.310 1.500 3.030 ;
        RECT  3.790 1.210 4.030 3.190 ;
        RECT  0.160 3.910 0.560 4.380 ;
        RECT  0.160 3.910 3.920 4.150 ;
        RECT  0.720 2.050 0.960 4.150 ;
        RECT  0.780 0.670 1.020 2.290 ;
        RECT  0.190 0.670 1.020 0.910 ;
    END
END DLHRBN

MACRO DLHRBP
    CLASS CORE ;
    FOREIGN DLHRBP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.540 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.760 2.930 2.700 ;
        RECT  2.500 2.050 2.930 2.450 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.410 0.480 2.430 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.180 0.450 2.750 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.370 1.260 10.370 1.540 ;
        RECT  10.090 1.260 10.370 3.220 ;
        RECT  9.380 2.940 10.370 3.220 ;
        RECT  9.370 1.250 9.770 1.540 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.860 3.550 2.870 ;
        RECT  3.210 2.180 3.550 2.580 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.450 8.510 3.300 ;
        RECT  8.200 2.900 8.510 3.300 ;
        RECT  7.770 1.450 8.510 1.730 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.060 -0.380 6.460 0.940 ;
        RECT  6.990 -0.380 7.390 0.560 ;
        RECT  8.570 -0.380 8.970 0.560 ;
        RECT  9.980 -0.380 10.380 0.780 ;
        RECT  0.000 -0.380 10.540 0.380 ;
        RECT  1.260 -0.380 2.330 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 4.480 2.940 5.420 ;
        RECT  6.630 4.480 7.030 5.420 ;
        RECT  7.500 4.260 7.900 5.420 ;
        RECT  8.740 4.260 9.140 5.420 ;
        RECT  9.980 4.260 10.380 5.420 ;
        RECT  0.000 4.660 10.540 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.910 2.920 7.190 3.160 ;
        RECT  5.910 1.460 6.150 3.160 ;
        RECT  8.870 2.060 9.760 2.300 ;
        RECT  8.870 0.970 9.110 2.300 ;
        RECT  5.910 1.460 7.250 1.700 ;
        RECT  7.010 0.970 7.250 1.700 ;
        RECT  7.010 0.970 9.110 1.210 ;
        RECT  4.760 4.180 6.250 4.420 ;
        RECT  6.010 3.700 6.250 4.420 ;
        RECT  4.760 0.620 5.000 4.420 ;
        RECT  6.010 3.700 7.670 3.940 ;
        RECT  7.430 2.020 7.670 3.940 ;
        RECT  2.020 0.800 2.260 3.190 ;
        RECT  2.020 0.800 2.810 1.040 ;
        RECT  4.630 0.620 5.000 1.020 ;
        RECT  2.570 0.620 5.000 0.860 ;
        RECT  5.350 3.700 5.750 3.940 ;
        RECT  5.350 0.620 5.590 3.940 ;
        RECT  4.280 1.750 4.520 4.420 ;
        RECT  1.200 3.430 4.520 3.670 ;
        RECT  1.200 2.790 1.440 3.670 ;
        RECT  1.260 1.310 1.500 3.030 ;
        RECT  3.790 1.210 4.030 3.190 ;
        RECT  3.180 4.170 3.920 4.410 ;
        RECT  0.160 3.910 0.560 4.380 ;
        RECT  3.180 3.910 3.420 4.410 ;
        RECT  0.160 3.910 3.420 4.150 ;
        RECT  0.720 2.050 0.960 4.150 ;
        RECT  0.780 0.670 1.020 2.290 ;
        RECT  0.190 0.670 1.020 0.910 ;
    END
END DLHRBP

MACRO DLHRBS
    CLASS CORE ;
    FOREIGN DLHRBS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.300 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.760 2.930 2.700 ;
        RECT  2.500 2.050 2.930 2.450 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.410 0.480 2.430 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.180 0.450 2.750 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.820 2.790 9.130 3.190 ;
        RECT  8.850 1.280 9.130 3.300 ;
        RECT  8.820 1.280 9.130 1.680 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.860 3.550 2.870 ;
        RECT  3.210 2.180 3.550 2.580 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.430 2.790 7.890 3.190 ;
        RECT  7.610 1.280 7.890 3.300 ;
        RECT  7.430 1.280 7.890 1.680 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.310 -0.380 6.710 0.560 ;
        RECT  8.140 -0.380 8.540 0.560 ;
        RECT  0.000 -0.380 9.300 0.380 ;
        RECT  1.260 -0.380 2.330 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 4.480 2.940 5.420 ;
        RECT  6.630 4.480 7.030 5.420 ;
        RECT  8.070 4.480 8.470 5.420 ;
        RECT  0.000 4.660 9.300 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.830 2.870 6.440 3.110 ;
        RECT  5.830 0.800 6.070 3.110 ;
        RECT  8.250 2.150 8.580 2.550 ;
        RECT  8.250 0.800 8.490 2.550 ;
        RECT  5.830 1.460 6.440 1.700 ;
        RECT  5.830 0.800 8.490 1.040 ;
        RECT  4.760 4.180 6.250 4.420 ;
        RECT  6.950 2.020 7.190 4.230 ;
        RECT  6.010 3.990 7.190 4.230 ;
        RECT  4.760 0.620 5.000 4.420 ;
        RECT  2.020 0.800 2.260 3.190 ;
        RECT  2.020 0.800 2.810 1.040 ;
        RECT  4.630 0.620 5.000 1.020 ;
        RECT  2.570 0.620 5.000 0.860 ;
        RECT  5.350 3.700 5.750 3.940 ;
        RECT  5.350 0.620 5.590 3.940 ;
        RECT  4.280 1.750 4.520 4.420 ;
        RECT  1.200 3.430 4.520 3.670 ;
        RECT  1.200 2.790 1.440 3.670 ;
        RECT  1.260 1.310 1.500 3.030 ;
        RECT  3.790 1.210 4.030 3.190 ;
        RECT  0.160 3.910 0.560 4.380 ;
        RECT  0.160 3.910 3.920 4.150 ;
        RECT  0.720 2.050 0.960 4.150 ;
        RECT  0.780 0.670 1.020 2.290 ;
        RECT  0.190 0.670 1.020 0.910 ;
    END
END DLHRBS

MACRO DLHS
    CLASS CORE ;
    FOREIGN DLHS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.230 1.800 2.630 ;
        RECT  1.410 1.820 1.690 2.770 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 0.920 8.510 3.200 ;
        RECT  8.200 2.800 8.510 3.200 ;
        RECT  8.200 0.920 8.510 1.320 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.680 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.880 0.760 7.160 1.830 ;
        RECT  6.990 1.550 7.270 3.190 ;
        RECT  6.760 2.790 7.270 3.190 ;
        RECT  6.760 0.760 7.160 1.160 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.580 -0.380 2.980 0.560 ;
        RECT  5.960 -0.380 6.360 0.560 ;
        RECT  7.400 -0.380 7.800 1.080 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  1.040 -0.380 1.440 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.110 3.910 2.510 5.420 ;
        RECT  5.380 4.480 5.780 5.420 ;
        RECT  7.400 4.260 7.800 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.160 3.140 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.280 3.780 7.940 4.020 ;
        RECT  7.700 2.160 7.940 4.020 ;
        RECT  6.170 3.590 6.570 3.830 ;
        RECT  6.280 1.570 6.520 4.020 ;
        RECT  5.340 2.420 6.520 2.660 ;
        RECT  5.340 2.260 5.580 2.660 ;
        RECT  6.170 1.570 6.570 1.810 ;
        RECT  4.010 3.680 4.320 4.080 ;
        RECT  4.080 0.790 4.320 4.080 ;
        RECT  4.050 2.860 4.320 3.260 ;
        RECT  4.080 1.560 4.390 1.960 ;
        RECT  5.940 0.800 6.340 1.100 ;
        RECT  4.000 0.800 6.340 1.040 ;
        RECT  4.000 0.790 4.400 1.040 ;
        RECT  4.830 2.860 5.110 3.260 ;
        RECT  4.830 1.570 5.070 3.260 ;
        RECT  4.790 1.570 5.190 1.810 ;
        RECT  0.920 3.060 1.200 3.460 ;
        RECT  3.330 2.860 3.580 3.260 ;
        RECT  3.340 0.800 3.580 3.260 ;
        RECT  0.920 0.800 1.160 3.460 ;
        RECT  3.340 1.560 3.670 1.960 ;
        RECT  0.240 0.800 0.480 1.730 ;
        RECT  0.240 0.800 3.580 1.040 ;
        RECT  2.850 3.830 3.150 4.230 ;
        RECT  2.850 1.520 3.090 4.230 ;
        RECT  2.850 2.190 3.100 2.590 ;
        RECT  2.660 1.520 3.090 1.920 ;
        RECT  1.380 3.910 1.780 4.150 ;
        RECT  1.540 3.270 1.780 4.150 ;
        RECT  1.540 3.270 2.610 3.510 ;
        RECT  2.060 3.110 2.610 3.510 ;
        RECT  2.060 1.340 2.300 3.510 ;
        RECT  1.660 1.340 2.300 1.580 ;
    END
END DLHS

MACRO FA1
    CLASS CORE ;
    FOREIGN FA1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.050 0.620 15.330 3.190 ;
        RECT  15.020 2.790 15.330 3.190 ;
        RECT  15.020 1.240 15.330 1.640 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.390 4.000 5.290 4.240 ;
        RECT  5.050 4.180 9.730 4.420 ;
        RECT  8.850 3.980 12.210 4.220 ;
        RECT  13.790 2.460 14.710 2.740 ;
        RECT  14.430 2.460 14.710 4.320 ;
        RECT  11.970 4.080 14.710 4.320 ;
        RECT  1.390 4.080 2.630 4.320 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.240 0.480 1.640 ;
        RECT  0.170 2.790 0.480 3.190 ;
        RECT  0.170 0.620 0.450 3.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.630 12.230 2.870 ;
        RECT  10.090 2.300 10.370 3.300 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.290 0.620 9.750 0.860 ;
        RECT  9.470 0.620 9.750 1.230 ;
        RECT  9.470 0.950 10.990 1.230 ;
        RECT  10.710 0.950 10.990 2.100 ;
        RECT  10.710 1.820 12.850 2.100 ;
        RECT  12.570 1.820 12.850 2.740 ;
        RECT  12.570 2.210 13.070 2.610 ;
        RECT  6.170 0.850 6.530 1.250 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.480 -0.380 4.880 0.560 ;
        RECT  5.650 -0.380 6.050 0.560 ;
        RECT  10.490 -0.380 10.890 0.560 ;
        RECT  11.940 -0.380 12.340 0.560 ;
        RECT  14.410 -0.380 14.810 0.860 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.940 -0.380 1.340 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.410 4.480 4.810 5.420 ;
        RECT  10.330 4.480 11.730 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.700 4.260 1.100 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  12.980 3.020 13.550 3.260 ;
        RECT  13.310 1.300 13.550 3.260 ;
        RECT  13.310 1.940 14.790 2.180 ;
        RECT  14.390 1.860 14.790 2.180 ;
        RECT  13.070 1.300 13.550 1.700 ;
        RECT  13.790 0.820 14.030 1.700 ;
        RECT  11.230 0.820 11.470 1.500 ;
        RECT  11.230 0.820 14.030 1.060 ;
        RECT  10.920 3.500 14.030 3.740 ;
        RECT  13.790 3.030 14.030 3.740 ;
        RECT  10.920 3.280 11.320 3.740 ;
        RECT  9.550 1.580 9.790 3.530 ;
        RECT  9.300 2.150 9.790 2.550 ;
        RECT  9.550 1.580 10.150 1.820 ;
        RECT  8.820 3.130 9.070 3.530 ;
        RECT  5.800 1.500 6.040 3.200 ;
        RECT  8.820 1.100 9.060 3.530 ;
        RECT  6.770 2.100 7.090 2.500 ;
        RECT  5.800 2.190 7.090 2.430 ;
        RECT  6.770 1.100 7.010 2.500 ;
        RECT  8.820 1.500 9.210 1.900 ;
        RECT  5.800 1.500 6.110 1.900 ;
        RECT  6.770 1.100 9.060 1.340 ;
        RECT  5.570 3.700 8.210 3.940 ;
        RECT  7.970 1.580 8.210 3.940 ;
        RECT  7.970 1.580 8.570 1.820 ;
        RECT  7.100 3.110 7.570 3.350 ;
        RECT  7.330 1.580 7.570 3.350 ;
        RECT  7.310 1.580 7.710 1.820 ;
        RECT  2.420 3.520 5.320 3.760 ;
        RECT  5.080 1.420 5.320 3.760 ;
        RECT  2.420 1.550 2.660 3.760 ;
        RECT  2.260 2.960 2.660 3.360 ;
        RECT  4.240 1.990 4.480 2.390 ;
        RECT  4.240 2.070 5.320 2.310 ;
        RECT  5.080 1.420 5.390 1.820 ;
        RECT  2.330 1.420 2.570 1.820 ;
        RECT  3.620 3.040 4.020 3.280 ;
        RECT  3.700 1.420 3.940 3.280 ;
        RECT  3.700 1.420 4.010 1.820 ;
        RECT  2.900 3.040 3.300 3.280 ;
        RECT  2.980 0.800 3.220 3.280 ;
        RECT  0.690 2.130 1.050 2.530 ;
        RECT  0.810 0.800 1.050 2.530 ;
        RECT  2.980 1.420 3.290 1.820 ;
        RECT  0.810 0.800 3.220 1.040 ;
        RECT  1.540 3.010 1.780 3.410 ;
        RECT  1.550 1.310 1.790 3.300 ;
        RECT  1.550 2.130 2.030 2.530 ;
        RECT  1.530 1.310 1.930 1.550 ;
    END
END FA1

MACRO FA1P
    CLASS CORE ;
    FOREIGN FA1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.740 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 1.260 16.570 3.130 ;
        RECT  15.460 2.850 16.570 3.130 ;
        RECT  15.050 1.260 16.570 1.540 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.940 1.070 3.220 ;
        RECT  0.170 1.260 1.090 1.540 ;
        RECT  0.170 1.260 0.450 3.220 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.650 2.630 12.740 2.870 ;
        RECT  10.710 2.300 10.990 3.300 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 4.000 5.850 4.240 ;
        RECT  5.610 4.180 10.350 4.420 ;
        RECT  9.360 3.980 12.720 4.220 ;
        RECT  14.300 2.480 15.220 2.720 ;
        RECT  14.980 2.480 15.220 4.320 ;
        RECT  14.980 3.520 15.310 4.320 ;
        RECT  12.480 4.080 15.310 4.320 ;
        RECT  2.030 4.000 2.930 4.320 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.760 0.620 10.370 0.860 ;
        RECT  10.090 0.620 10.370 1.230 ;
        RECT  10.090 0.950 11.470 1.230 ;
        RECT  11.190 0.950 11.470 2.100 ;
        RECT  11.190 1.820 12.850 2.100 ;
        RECT  12.570 1.860 13.470 2.140 ;
        RECT  13.190 1.860 13.470 2.740 ;
        RECT  13.190 2.210 13.580 2.610 ;
        RECT  6.680 0.850 7.000 1.250 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.680 -0.380 2.080 0.560 ;
        RECT  4.940 -0.380 5.340 0.560 ;
        RECT  6.060 -0.380 6.460 0.560 ;
        RECT  11.000 -0.380 11.400 0.560 ;
        RECT  12.450 -0.380 12.850 0.560 ;
        RECT  14.920 -0.380 15.340 0.780 ;
        RECT  16.180 -0.380 16.580 0.780 ;
        RECT  0.000 -0.380 16.740 0.380 ;
        RECT  0.170 -0.380 0.570 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 4.180 1.720 5.420 ;
        RECT  4.920 4.480 5.320 5.420 ;
        RECT  10.840 4.480 12.240 5.420 ;
        RECT  16.180 4.260 16.580 5.420 ;
        RECT  0.000 4.660 16.740 5.420 ;
        RECT  0.160 4.120 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.490 3.020 14.060 3.260 ;
        RECT  13.820 1.380 14.060 3.260 ;
        RECT  13.820 2.000 15.300 2.240 ;
        RECT  14.900 1.860 15.300 2.240 ;
        RECT  13.500 1.380 14.060 1.620 ;
        RECT  14.300 0.900 14.540 1.700 ;
        RECT  11.740 0.900 11.980 1.500 ;
        RECT  11.740 0.900 14.540 1.140 ;
        RECT  11.430 3.500 14.540 3.740 ;
        RECT  14.300 3.030 14.540 3.740 ;
        RECT  11.430 3.280 11.830 3.740 ;
        RECT  10.070 1.580 10.310 3.530 ;
        RECT  9.820 2.170 10.310 2.570 ;
        RECT  10.070 1.580 10.660 1.820 ;
        RECT  9.340 1.100 9.580 3.530 ;
        RECT  6.310 2.800 6.560 3.200 ;
        RECT  6.310 1.500 6.550 3.200 ;
        RECT  7.340 2.100 7.600 2.500 ;
        RECT  6.310 2.190 7.600 2.430 ;
        RECT  7.340 1.100 7.580 2.500 ;
        RECT  6.310 1.500 6.620 1.900 ;
        RECT  7.340 1.100 9.580 1.340 ;
        RECT  6.090 3.700 8.730 3.940 ;
        RECT  8.490 1.580 8.730 3.940 ;
        RECT  8.490 1.580 8.940 1.820 ;
        RECT  7.620 3.110 8.080 3.350 ;
        RECT  7.840 1.580 8.080 3.350 ;
        RECT  7.820 1.580 8.220 1.820 ;
        RECT  2.840 3.520 5.840 3.760 ;
        RECT  5.600 1.420 5.840 3.760 ;
        RECT  2.840 1.420 3.080 3.760 ;
        RECT  2.780 2.960 3.080 3.360 ;
        RECT  4.750 1.990 4.990 2.390 ;
        RECT  4.750 2.070 5.840 2.310 ;
        RECT  5.600 1.420 5.900 1.820 ;
        RECT  4.140 3.040 4.540 3.280 ;
        RECT  4.210 1.420 4.450 3.280 ;
        RECT  4.210 1.420 4.520 1.820 ;
        RECT  3.420 3.040 3.820 3.280 ;
        RECT  3.560 0.800 3.800 3.280 ;
        RECT  1.200 2.030 1.570 2.430 ;
        RECT  1.330 0.800 1.570 2.430 ;
        RECT  1.330 0.800 3.800 1.040 ;
        RECT  2.060 3.010 2.310 3.410 ;
        RECT  2.070 1.360 2.310 3.410 ;
        RECT  2.070 2.130 2.550 2.530 ;
        RECT  2.040 1.360 2.440 1.600 ;
    END
END FA1P

MACRO FA1S
    CLASS CORE ;
    FOREIGN FA1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.570 4.790 3.110 ;
        RECT  4.500 2.870 4.900 3.110 ;
        RECT  4.380 1.570 4.790 1.810 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 3.890 6.630 4.420 ;
        RECT  7.400 3.830 9.130 4.130 ;
        RECT  3.320 3.890 10.370 4.130 ;
        RECT  10.090 2.560 10.370 4.130 ;
        RECT  1.960 4.080 3.560 4.320 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 0.620 11.610 3.190 ;
        RECT  11.300 2.790 11.610 3.190 ;
        RECT  11.300 1.490 11.610 1.890 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.300 3.350 6.700 3.650 ;
        RECT  2.840 3.350 9.750 3.590 ;
        RECT  2.680 3.450 9.750 3.590 ;
        RECT  9.470 2.330 9.750 3.590 ;
        RECT  9.400 2.330 9.800 2.570 ;
        RECT  0.390 3.520 3.080 3.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.240 1.390 2.640 ;
        RECT  0.790 0.700 2.310 0.980 ;
        RECT  2.030 0.700 2.310 1.310 ;
        RECT  3.890 0.700 4.170 1.310 ;
        RECT  2.030 1.030 4.170 1.310 ;
        RECT  3.890 0.700 4.790 0.980 ;
        RECT  4.510 0.700 4.790 1.330 ;
        RECT  5.400 1.090 5.640 2.530 ;
        RECT  5.400 2.130 5.880 2.530 ;
        RECT  7.610 0.700 7.890 1.330 ;
        RECT  4.510 1.090 7.890 1.330 ;
        RECT  7.610 0.700 9.750 0.980 ;
        RECT  9.470 0.800 10.370 1.270 ;
        RECT  0.790 0.700 1.070 2.740 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.800 -0.380 3.200 0.560 ;
        RECT  5.220 -0.380 7.070 0.850 ;
        RECT  10.360 -0.380 10.760 0.560 ;
        RECT  0.000 -0.380 11.780 0.380 ;
        RECT  0.140 -0.380 0.550 0.920 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.800 4.480 4.200 5.420 ;
        RECT  5.110 4.480 5.510 5.420 ;
        RECT  6.890 4.480 7.290 5.420 ;
        RECT  0.000 4.660 11.780 5.420 ;
        RECT  0.970 4.480 1.370 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.430 2.870 8.830 3.110 ;
        RECT  8.510 1.490 8.750 3.110 ;
        RECT  10.650 2.070 11.050 2.460 ;
        RECT  10.110 2.070 11.050 2.310 ;
        RECT  8.510 1.840 10.350 2.080 ;
        RECT  8.460 1.490 8.750 1.890 ;
        RECT  6.070 2.870 8.030 3.110 ;
        RECT  5.900 1.570 7.920 1.810 ;
        RECT  2.450 2.870 2.850 3.110 ;
        RECT  2.530 2.140 2.770 3.110 ;
        RECT  3.960 2.080 4.200 2.480 ;
        RECT  1.630 2.140 4.200 2.380 ;
        RECT  1.630 1.490 1.870 2.380 ;
        RECT  1.360 1.490 1.870 1.890 ;
        RECT  2.140 1.570 4.060 1.810 ;
        RECT  0.160 2.980 2.120 3.220 ;
        RECT  1.720 2.870 2.120 3.220 ;
        RECT  0.160 2.870 0.560 3.220 ;
    END
END FA1S

MACRO FA1T
    CLASS CORE ;
    FOREIGN FA1T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.980 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.780 1.260 17.820 1.540 ;
        RECT  16.180 2.940 17.820 3.220 ;
        RECT  16.910 1.260 17.190 3.220 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 2.940 1.800 3.220 ;
        RECT  0.160 1.260 1.820 1.540 ;
        RECT  0.790 1.260 1.070 3.220 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.630 13.470 2.870 ;
        RECT  11.330 2.300 11.610 3.300 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.760 4.000 6.580 4.240 ;
        RECT  9.980 3.980 10.730 4.420 ;
        RECT  6.340 4.180 12.100 4.420 ;
        RECT  11.860 3.980 14.070 4.220 ;
        RECT  15.030 2.470 15.940 2.730 ;
        RECT  15.680 2.470 15.940 4.320 ;
        RECT  13.830 4.080 15.950 4.320 ;
        RECT  15.680 3.520 16.740 3.760 ;
        RECT  2.760 4.000 3.660 4.320 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.490 0.620 11.100 0.860 ;
        RECT  10.820 0.620 11.100 1.230 ;
        RECT  10.820 0.950 12.200 1.230 ;
        RECT  11.920 0.950 12.200 2.100 ;
        RECT  11.920 1.820 13.580 2.100 ;
        RECT  13.300 1.860 14.090 2.140 ;
        RECT  13.810 1.860 14.090 2.740 ;
        RECT  13.810 2.210 14.310 2.610 ;
        RECT  7.410 0.850 7.730 1.250 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.410 -0.380 2.810 0.560 ;
        RECT  5.670 -0.380 6.070 0.560 ;
        RECT  6.790 -0.380 7.190 0.560 ;
        RECT  11.730 -0.380 12.130 0.560 ;
        RECT  13.180 -0.380 13.580 0.560 ;
        RECT  15.640 -0.380 16.060 0.780 ;
        RECT  16.910 -0.380 17.310 0.780 ;
        RECT  0.000 -0.380 17.980 0.380 ;
        RECT  0.850 -0.380 1.250 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.110 4.180 2.450 5.420 ;
        RECT  5.650 4.480 6.050 5.420 ;
        RECT  12.340 4.480 13.240 5.420 ;
        RECT  16.900 4.120 17.300 5.420 ;
        RECT  0.000 4.660 17.980 5.420 ;
        RECT  0.890 4.120 1.290 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  14.220 3.020 14.790 3.260 ;
        RECT  14.550 1.380 14.790 3.260 ;
        RECT  14.550 1.970 16.030 2.210 ;
        RECT  15.630 1.860 16.030 2.210 ;
        RECT  14.230 1.380 14.790 1.620 ;
        RECT  15.030 0.900 15.270 1.700 ;
        RECT  12.470 0.900 12.710 1.500 ;
        RECT  12.470 0.900 15.270 1.140 ;
        RECT  12.160 3.500 15.270 3.740 ;
        RECT  15.030 3.030 15.270 3.740 ;
        RECT  12.160 3.280 12.560 3.740 ;
        RECT  10.800 3.130 11.070 3.530 ;
        RECT  10.830 1.580 11.070 3.530 ;
        RECT  10.550 2.150 11.070 2.550 ;
        RECT  10.830 1.580 11.390 1.820 ;
        RECT  10.070 1.100 10.310 3.530 ;
        RECT  7.040 2.800 7.290 3.200 ;
        RECT  7.040 1.500 7.280 3.200 ;
        RECT  8.010 2.100 8.330 2.500 ;
        RECT  7.040 2.190 8.330 2.430 ;
        RECT  8.010 1.100 8.250 2.500 ;
        RECT  7.040 1.500 7.350 1.900 ;
        RECT  8.010 1.100 10.310 1.340 ;
        RECT  6.820 3.700 9.460 3.940 ;
        RECT  9.220 1.580 9.460 3.940 ;
        RECT  9.220 1.580 9.670 1.820 ;
        RECT  8.350 3.110 8.810 3.350 ;
        RECT  8.570 1.580 8.810 3.350 ;
        RECT  8.550 1.580 8.950 1.820 ;
        RECT  3.660 3.520 6.570 3.760 ;
        RECT  6.330 1.420 6.570 3.760 ;
        RECT  3.660 1.420 3.900 3.760 ;
        RECT  3.510 2.960 3.900 3.360 ;
        RECT  5.480 1.990 5.720 2.390 ;
        RECT  5.480 2.070 6.570 2.310 ;
        RECT  6.330 1.420 6.630 1.820 ;
        RECT  3.570 1.420 3.900 1.820 ;
        RECT  4.870 3.040 5.270 3.280 ;
        RECT  4.940 1.420 5.180 3.280 ;
        RECT  4.940 1.420 5.250 1.820 ;
        RECT  4.150 3.040 4.550 3.280 ;
        RECT  4.220 0.800 4.460 3.280 ;
        RECT  1.430 2.030 2.300 2.430 ;
        RECT  2.060 0.800 2.300 2.430 ;
        RECT  4.220 1.420 4.530 1.820 ;
        RECT  2.060 0.800 4.460 1.040 ;
        RECT  2.790 3.010 3.040 3.410 ;
        RECT  2.800 1.360 3.040 3.410 ;
        RECT  2.800 2.130 3.280 2.530 ;
        RECT  2.770 1.360 3.170 1.600 ;
    END
END FA1T

MACRO FA2
    CLASS CORE ;
    FOREIGN FA2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.600 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.830 1.360 7.670 1.600 ;
        RECT  6.040 2.960 7.670 3.200 ;
        RECT  7.430 1.360 7.670 4.240 ;
        RECT  12.590 3.520 12.830 4.240 ;
        RECT  7.430 4.000 12.830 4.240 ;
        RECT  16.090 1.280 16.330 3.760 ;
        RECT  12.590 3.520 16.330 3.760 ;
        RECT  16.090 1.280 16.550 1.520 ;
        RECT  6.040 2.870 6.280 3.270 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.500 3.910 4.150 4.340 ;
        RECT  3.910 3.520 4.150 4.340 ;
        RECT  2.290 4.060 4.150 4.340 ;
        RECT  3.910 3.520 5.410 3.760 ;
        RECT  5.130 2.940 5.410 4.310 ;
        RECT  5.470 2.390 5.750 3.220 ;
        RECT  5.130 2.940 5.750 3.220 ;
        RECT  5.470 2.390 5.870 2.630 ;
        RECT  3.510 3.890 4.150 4.340 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.240 0.480 1.640 ;
        RECT  0.170 2.790 0.480 3.190 ;
        RECT  0.170 0.620 0.450 3.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 0.800 14.710 2.200 ;
        RECT  14.430 1.800 14.930 2.200 ;
        RECT  12.930 0.800 17.440 1.040 ;
        RECT  17.200 0.800 17.440 2.300 ;
        RECT  17.200 2.060 17.750 2.300 ;
        RECT  11.740 0.620 13.170 0.860 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.530 3.150 17.810 4.240 ;
        RECT  13.430 4.000 18.210 4.240 ;
        RECT  17.620 4.060 18.290 4.340 ;
        RECT  13.330 4.080 14.070 4.320 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.520 -0.380 4.920 0.560 ;
        RECT  7.180 -0.380 7.580 0.560 ;
        RECT  7.970 -0.380 8.370 0.560 ;
        RECT  10.970 -0.380 11.370 0.700 ;
        RECT  13.420 -0.380 13.820 0.560 ;
        RECT  16.800 -0.380 17.200 0.560 ;
        RECT  17.760 -0.380 18.160 0.560 ;
        RECT  0.000 -0.380 18.600 0.380 ;
        RECT  1.030 -0.380 1.970 0.720 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.570 4.080 1.970 5.420 ;
        RECT  4.370 4.480 4.770 5.420 ;
        RECT  4.370 4.560 6.100 5.420 ;
        RECT  7.140 4.480 7.540 5.420 ;
        RECT  7.970 4.480 8.370 5.420 ;
        RECT  10.970 4.480 11.370 5.420 ;
        RECT  12.700 4.480 13.100 5.420 ;
        RECT  14.310 4.480 15.790 5.420 ;
        RECT  16.990 4.480 17.390 5.420 ;
        RECT  0.000 4.660 18.600 5.420 ;
        RECT  0.740 4.170 1.140 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  18.120 3.060 18.410 3.460 ;
        RECT  18.170 1.520 18.410 3.460 ;
        RECT  16.570 2.540 18.410 2.780 ;
        RECT  16.570 1.830 16.810 2.780 ;
        RECT  17.760 1.520 18.410 1.760 ;
        RECT  14.390 2.800 14.630 3.200 ;
        RECT  14.390 2.800 15.610 3.040 ;
        RECT  15.370 1.340 15.610 3.040 ;
        RECT  15.190 1.340 15.610 1.580 ;
        RECT  13.520 1.500 13.760 3.200 ;
        RECT  10.330 1.100 10.570 3.200 ;
        RECT  12.450 2.260 12.810 2.660 ;
        RECT  12.450 2.340 13.760 2.580 ;
        RECT  12.450 1.100 12.690 2.660 ;
        RECT  10.330 1.100 12.690 1.340 ;
        RECT  8.890 3.520 11.770 3.760 ;
        RECT  11.530 2.960 11.770 3.760 ;
        RECT  8.890 1.240 9.130 3.760 ;
        RECT  11.530 2.960 12.130 3.200 ;
        RECT  11.890 1.580 12.130 3.200 ;
        RECT  11.810 1.580 12.210 1.820 ;
        RECT  11.050 1.580 11.290 3.200 ;
        RECT  10.910 2.140 11.290 2.540 ;
        RECT  10.970 1.580 11.370 1.820 ;
        RECT  9.610 0.760 9.850 3.200 ;
        RECT  8.610 0.760 9.850 1.000 ;
        RECT  2.370 0.800 2.610 3.270 ;
        RECT  8.050 1.270 8.290 3.200 ;
        RECT  7.910 1.820 8.290 2.220 ;
        RECT  7.970 1.270 8.370 1.510 ;
        RECT  7.970 0.800 8.210 1.510 ;
        RECT  2.370 0.800 8.210 1.040 ;
        RECT  3.810 1.280 4.050 3.270 ;
        RECT  4.720 1.840 4.960 2.730 ;
        RECT  6.950 1.840 7.190 2.720 ;
        RECT  3.810 2.410 4.960 2.650 ;
        RECT  4.720 1.840 7.190 2.080 ;
        RECT  0.720 3.550 3.250 3.790 ;
        RECT  3.010 1.360 3.250 3.790 ;
        RECT  0.720 1.920 0.960 3.790 ;
        RECT  3.010 2.950 3.410 3.190 ;
        RECT  0.690 1.870 0.930 2.270 ;
        RECT  3.010 1.360 3.410 1.600 ;
        RECT  1.570 2.870 1.970 3.110 ;
        RECT  1.650 1.320 1.890 3.110 ;
        RECT  1.650 1.880 2.030 2.280 ;
        RECT  1.570 1.320 1.970 1.560 ;
    END
END FA2

MACRO FA2P
    CLASS CORE ;
    FOREIGN FA2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.420 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.200 1.580 11.600 1.820 ;
        RECT  11.330 3.020 11.610 4.240 ;
        RECT  11.330 3.020 11.680 3.420 ;
        RECT  12.720 1.100 12.960 1.820 ;
        RECT  12.640 1.580 13.040 1.820 ;
        RECT  12.880 3.020 13.120 4.240 ;
        RECT  11.280 1.100 14.320 1.340 ;
        RECT  14.080 1.100 14.320 4.240 ;
        RECT  18.170 3.520 18.410 4.240 ;
        RECT  11.330 4.000 18.410 4.240 ;
        RECT  21.520 1.330 21.760 3.760 ;
        RECT  18.170 3.520 21.760 3.760 ;
        RECT  21.520 2.790 21.900 3.280 ;
        RECT  21.520 1.330 23.280 1.570 ;
        RECT  21.520 3.040 23.280 3.280 ;
        RECT  11.280 1.100 11.520 1.820 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.250 3.990 7.200 4.230 ;
        RECT  6.960 3.520 7.200 4.230 ;
        RECT  6.960 3.520 10.370 3.760 ;
        RECT  10.090 3.020 10.370 4.140 ;
        RECT  10.090 3.020 10.400 3.420 ;
        RECT  3.740 4.060 4.830 4.340 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.240 1.100 1.640 ;
        RECT  0.790 2.790 1.100 3.190 ;
        RECT  0.790 1.020 1.070 3.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  18.740 0.620 18.980 1.260 ;
        RECT  18.740 1.020 20.600 1.260 ;
        RECT  20.360 0.850 20.600 2.200 ;
        RECT  20.360 0.850 23.990 1.090 ;
        RECT  23.750 0.850 23.990 2.300 ;
        RECT  23.750 2.060 24.150 2.300 ;
        RECT  17.390 0.620 18.980 0.860 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  19.010 4.000 24.010 4.240 ;
        RECT  23.730 3.020 24.010 4.240 ;
        RECT  23.730 3.520 25.030 3.760 ;
        RECT  24.630 3.520 25.030 3.990 ;
        RECT  18.880 4.080 19.650 4.320 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 -0.380 2.720 0.720 ;
        RECT  5.070 -0.380 5.470 0.560 ;
        RECT  7.440 -0.380 7.840 0.560 ;
        RECT  9.080 -0.380 9.480 0.560 ;
        RECT  16.690 -0.380 17.090 0.700 ;
        RECT  19.220 -0.380 19.460 0.640 ;
        RECT  22.230 -0.380 22.630 0.560 ;
        RECT  23.600 -0.380 25.260 0.560 ;
        RECT  0.000 -0.380 25.420 0.380 ;
        RECT  0.160 -0.380 0.560 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.470 4.180 1.870 5.420 ;
        RECT  2.320 4.120 2.720 5.420 ;
        RECT  5.270 4.480 5.670 5.420 ;
        RECT  7.440 4.260 7.840 5.420 ;
        RECT  8.900 4.260 9.300 5.420 ;
        RECT  16.690 4.480 17.090 5.420 ;
        RECT  18.220 4.480 18.620 5.420 ;
        RECT  19.980 4.480 21.260 5.420 ;
        RECT  22.230 4.480 22.630 5.420 ;
        RECT  23.600 4.480 24.000 5.420 ;
        RECT  24.720 4.630 25.120 5.420 ;
        RECT  0.000 4.660 25.420 5.420 ;
        RECT  0.160 4.180 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  24.940 1.560 25.180 3.200 ;
        RECT  22.340 2.540 25.180 2.780 ;
        RECT  22.340 1.830 22.580 2.780 ;
        RECT  22.340 1.830 22.700 2.230 ;
        RECT  24.540 1.560 25.180 1.800 ;
        RECT  24.540 1.400 24.780 1.800 ;
        RECT  20.060 2.800 20.300 3.200 ;
        RECT  20.060 2.800 21.280 3.040 ;
        RECT  21.040 1.340 21.280 3.040 ;
        RECT  20.860 1.340 21.280 1.580 ;
        RECT  19.090 1.500 19.330 3.200 ;
        RECT  16.050 1.100 16.290 3.200 ;
        RECT  18.090 2.260 18.410 2.660 ;
        RECT  18.170 1.100 18.410 2.660 ;
        RECT  18.090 2.340 19.330 2.580 ;
        RECT  16.050 1.100 18.410 1.340 ;
        RECT  14.610 3.520 17.490 3.760 ;
        RECT  17.250 2.960 17.490 3.760 ;
        RECT  14.610 1.240 14.850 3.760 ;
        RECT  17.250 2.960 17.850 3.200 ;
        RECT  17.610 1.580 17.850 3.200 ;
        RECT  17.530 1.580 17.930 1.820 ;
        RECT  16.770 1.580 17.010 3.200 ;
        RECT  16.630 2.140 17.010 2.540 ;
        RECT  16.690 1.580 17.090 1.820 ;
        RECT  15.330 0.620 15.570 3.200 ;
        RECT  6.420 0.950 9.960 1.190 ;
        RECT  9.720 0.620 9.960 1.190 ;
        RECT  5.630 0.750 6.660 0.990 ;
        RECT  9.720 0.620 15.570 0.860 ;
        RECT  13.600 2.540 13.840 3.270 ;
        RECT  12.160 2.540 12.400 3.270 ;
        RECT  10.720 2.540 10.960 3.270 ;
        RECT  9.600 2.540 9.840 3.270 ;
        RECT  8.250 2.870 8.490 3.270 ;
        RECT  6.900 2.870 7.140 3.270 ;
        RECT  6.900 2.950 9.840 3.190 ;
        RECT  9.600 2.540 13.840 2.780 ;
        RECT  10.640 2.060 13.600 2.300 ;
        RECT  13.360 1.580 13.600 2.300 ;
        RECT  12.000 1.580 12.240 2.300 ;
        RECT  10.640 1.430 10.880 2.300 ;
        RECT  13.360 1.580 13.760 1.820 ;
        RECT  11.920 1.580 12.320 1.820 ;
        RECT  10.480 1.430 10.880 1.820 ;
        RECT  6.820 1.430 10.880 1.670 ;
        RECT  4.550 3.510 6.660 3.750 ;
        RECT  6.420 2.390 6.660 3.750 ;
        RECT  4.550 1.280 4.790 3.750 ;
        RECT  4.550 2.870 4.800 3.270 ;
        RECT  6.420 2.390 7.710 2.630 ;
        RECT  4.550 1.280 4.800 1.680 ;
        RECT  5.940 1.280 6.180 3.270 ;
        RECT  3.120 0.800 3.360 3.270 ;
        RECT  5.030 1.820 5.280 2.220 ;
        RECT  5.040 0.800 5.280 2.220 ;
        RECT  5.940 1.900 6.450 2.140 ;
        RECT  5.040 1.280 6.180 1.520 ;
        RECT  3.120 0.800 5.290 1.040 ;
        RECT  1.450 3.550 3.840 3.790 ;
        RECT  3.600 1.360 3.840 3.790 ;
        RECT  1.450 1.920 1.690 3.790 ;
        RECT  3.600 2.950 4.160 3.190 ;
        RECT  1.420 1.870 1.660 2.270 ;
        RECT  3.600 1.360 4.160 1.600 ;
        RECT  2.320 2.870 2.720 3.110 ;
        RECT  2.400 1.320 2.640 3.110 ;
        RECT  2.400 1.880 2.780 2.280 ;
        RECT  2.320 1.320 2.720 1.560 ;
    END
END FA2P

MACRO FA2S
    CLASS CORE ;
    FOREIGN FA2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.170 2.870 7.450 3.270 ;
        RECT  7.210 1.240 7.450 4.320 ;
        RECT  7.210 4.080 9.670 4.320 ;
        RECT  9.220 4.000 11.610 4.240 ;
        RECT  11.330 3.340 11.610 4.240 ;
        RECT  14.850 1.280 15.090 3.760 ;
        RECT  11.330 3.520 15.090 3.760 ;
        RECT  14.850 3.060 15.230 3.460 ;
        RECT  14.850 1.310 15.310 1.550 ;
        RECT  7.170 1.240 7.450 1.640 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.990 4.060 4.290 4.340 ;
        RECT  6.390 1.280 6.630 2.080 ;
        RECT  6.390 1.790 6.970 2.080 ;
        RECT  3.500 4.000 6.930 4.240 ;
        RECT  6.690 1.790 6.930 4.240 ;
        RECT  6.690 1.790 6.970 2.190 ;
        RECT  3.500 3.810 3.900 4.340 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.420 0.480 1.820 ;
        RECT  0.170 2.790 0.480 3.190 ;
        RECT  0.170 0.620 0.450 3.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.690 0.800 13.930 2.200 ;
        RECT  11.930 0.800 17.170 1.040 ;
        RECT  16.930 0.800 17.170 2.320 ;
        RECT  16.110 2.080 17.170 2.320 ;
        RECT  10.740 0.620 12.170 0.860 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 3.040 16.570 4.240 ;
        RECT  12.330 4.000 16.970 4.240 ;
        RECT  16.380 4.060 17.050 4.340 ;
        RECT  12.330 4.000 12.830 4.320 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.600 -0.380 6.000 0.560 ;
        RECT  9.970 -0.380 10.370 0.700 ;
        RECT  12.420 -0.380 12.820 0.560 ;
        RECT  14.850 -0.380 16.920 0.560 ;
        RECT  0.000 -0.380 17.360 0.380 ;
        RECT  0.700 -0.380 1.640 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.520 4.480 6.090 5.420 ;
        RECT  9.970 4.480 10.370 5.420 ;
        RECT  11.700 4.480 12.100 5.420 ;
        RECT  13.240 4.480 15.800 5.420 ;
        RECT  0.000 4.660 17.360 5.420 ;
        RECT  0.160 4.280 1.640 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  16.880 2.560 17.120 3.460 ;
        RECT  15.570 2.560 17.120 2.800 ;
        RECT  15.570 1.600 15.810 2.800 ;
        RECT  15.330 1.830 15.810 2.230 ;
        RECT  16.420 1.440 16.660 1.840 ;
        RECT  15.570 1.600 16.660 1.840 ;
        RECT  13.390 2.800 13.630 3.200 ;
        RECT  13.390 2.800 14.610 3.040 ;
        RECT  14.370 1.340 14.610 3.040 ;
        RECT  14.190 1.340 14.610 1.580 ;
        RECT  12.520 1.500 12.760 3.200 ;
        RECT  9.330 1.100 9.570 3.200 ;
        RECT  11.450 2.260 11.810 2.660 ;
        RECT  11.450 2.340 12.760 2.580 ;
        RECT  11.450 1.100 11.690 2.660 ;
        RECT  9.330 1.100 11.690 1.340 ;
        RECT  7.890 3.520 10.770 3.760 ;
        RECT  10.530 2.960 10.770 3.760 ;
        RECT  7.890 1.240 8.130 3.760 ;
        RECT  10.530 2.960 11.130 3.200 ;
        RECT  10.890 1.580 11.130 3.200 ;
        RECT  10.810 1.580 11.210 1.820 ;
        RECT  10.050 1.580 10.290 3.200 ;
        RECT  9.910 2.140 10.290 2.540 ;
        RECT  9.970 1.580 10.370 1.820 ;
        RECT  8.610 0.760 8.850 3.200 ;
        RECT  4.880 0.800 6.760 1.040 ;
        RECT  6.520 0.760 8.850 1.000 ;
        RECT  4.140 3.450 6.300 3.690 ;
        RECT  6.060 2.330 6.300 3.690 ;
        RECT  3.780 3.230 4.380 3.470 ;
        RECT  3.780 2.830 4.050 3.470 ;
        RECT  3.780 1.280 4.020 3.470 ;
        RECT  6.060 2.330 6.310 2.730 ;
        RECT  3.780 1.280 4.050 1.680 ;
        RECT  2.370 0.800 2.610 3.230 ;
        RECT  5.110 2.870 5.620 3.110 ;
        RECT  5.380 1.280 5.620 3.110 ;
        RECT  4.280 1.820 4.520 2.220 ;
        RECT  4.280 1.820 5.620 2.060 ;
        RECT  5.230 1.280 5.620 2.060 ;
        RECT  4.290 0.800 4.530 2.060 ;
        RECT  2.370 0.800 4.530 1.040 ;
        RECT  0.720 3.550 3.090 3.790 ;
        RECT  2.850 1.360 3.090 3.790 ;
        RECT  0.720 2.130 0.960 3.790 ;
        RECT  2.850 2.830 3.330 3.230 ;
        RECT  0.690 2.080 0.930 2.480 ;
        RECT  2.850 1.360 3.410 1.600 ;
        RECT  1.570 2.870 1.970 3.110 ;
        RECT  1.650 1.500 1.890 3.110 ;
        RECT  1.650 2.190 2.080 2.590 ;
        RECT  1.570 1.500 1.970 1.740 ;
    END
END FA2S

MACRO FA3
    CLASS CORE ;
    FOREIGN FA3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.600 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.830 1.360 7.670 1.600 ;
        RECT  5.980 2.960 7.670 3.200 ;
        RECT  7.430 1.360 7.670 4.240 ;
        RECT  12.970 3.520 13.210 4.240 ;
        RECT  7.430 4.000 13.210 4.240 ;
        RECT  16.090 1.310 16.330 3.760 ;
        RECT  16.090 1.310 16.550 1.550 ;
        RECT  16.090 2.470 16.570 3.760 ;
        RECT  12.970 3.520 16.570 3.760 ;
        RECT  5.980 2.870 6.220 3.270 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.990 4.060 4.130 4.340 ;
        RECT  3.500 4.000 4.790 4.240 ;
        RECT  4.510 3.030 4.790 4.240 ;
        RECT  5.470 2.390 5.710 3.270 ;
        RECT  4.510 3.030 5.710 3.270 ;
        RECT  5.470 2.390 5.870 2.630 ;
        RECT  3.500 3.810 3.900 4.340 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.420 0.480 1.820 ;
        RECT  0.170 2.790 0.480 3.190 ;
        RECT  0.170 0.620 0.450 3.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.330 2.240 12.850 2.640 ;
        RECT  12.570 1.420 12.850 2.640 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.420 13.470 2.640 ;
        RECT  13.130 2.210 13.470 2.610 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.520 -0.380 4.920 0.560 ;
        RECT  7.180 -0.380 9.210 0.560 ;
        RECT  11.600 -0.380 12.000 0.700 ;
        RECT  12.670 -0.380 13.070 0.560 ;
        RECT  16.800 -0.380 17.200 0.560 ;
        RECT  17.760 -0.380 18.160 0.560 ;
        RECT  0.000 -0.380 18.600 0.380 ;
        RECT  1.030 -0.380 1.970 0.720 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.570 4.080 1.970 5.420 ;
        RECT  4.370 4.480 4.770 5.420 ;
        RECT  7.140 4.480 9.160 5.420 ;
        RECT  11.600 4.480 12.000 5.420 ;
        RECT  12.560 4.480 12.960 5.420 ;
        RECT  14.460 4.480 15.940 5.420 ;
        RECT  16.990 4.480 17.390 5.420 ;
        RECT  0.000 4.660 18.600 5.420 ;
        RECT  0.740 4.170 1.140 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  16.870 3.140 18.440 3.380 ;
        RECT  16.870 1.650 17.110 3.380 ;
        RECT  16.570 1.830 17.110 2.230 ;
        RECT  17.660 1.440 17.900 1.890 ;
        RECT  16.870 1.650 17.900 1.890 ;
        RECT  9.210 3.440 9.610 3.730 ;
        RECT  9.210 3.440 12.400 3.680 ;
        RECT  12.160 2.960 12.400 3.680 ;
        RECT  10.960 1.240 11.200 3.680 ;
        RECT  12.160 2.960 14.030 3.200 ;
        RECT  13.710 1.350 13.950 3.200 ;
        RECT  17.350 2.130 18.410 2.370 ;
        RECT  18.170 0.800 18.410 2.370 ;
        RECT  13.710 1.960 15.150 2.200 ;
        RECT  14.910 0.800 15.150 2.200 ;
        RECT  14.910 0.800 18.410 1.040 ;
        RECT  13.800 4.000 18.210 4.240 ;
        RECT  14.610 2.800 14.850 3.200 ;
        RECT  14.610 2.800 15.830 3.040 ;
        RECT  15.590 1.340 15.830 3.040 ;
        RECT  15.410 1.340 15.830 1.580 ;
        RECT  11.540 2.800 11.920 3.200 ;
        RECT  11.540 0.940 11.780 3.200 ;
        RECT  11.540 1.580 12.000 1.820 ;
        RECT  11.540 0.940 12.810 1.180 ;
        RECT  12.570 0.800 14.310 1.040 ;
        RECT  10.240 0.840 10.480 3.200 ;
        RECT  8.610 0.840 8.850 2.350 ;
        RECT  8.610 0.840 10.480 1.080 ;
        RECT  9.520 1.320 9.760 3.200 ;
        RECT  9.440 1.320 9.840 1.560 ;
        RECT  2.360 2.870 2.610 3.270 ;
        RECT  8.050 1.340 8.290 3.200 ;
        RECT  2.360 0.800 2.600 3.270 ;
        RECT  7.910 1.820 8.290 2.220 ;
        RECT  2.360 1.280 2.610 1.680 ;
        RECT  7.970 1.340 8.370 1.580 ;
        RECT  7.970 0.800 8.210 1.580 ;
        RECT  2.360 0.800 8.210 1.040 ;
        RECT  3.960 0.760 4.360 1.040 ;
        RECT  3.810 1.280 4.050 3.270 ;
        RECT  4.720 1.840 4.960 2.730 ;
        RECT  6.950 1.840 7.190 2.720 ;
        RECT  3.810 2.410 4.960 2.650 ;
        RECT  4.720 1.840 7.190 2.080 ;
        RECT  0.720 3.550 3.090 3.790 ;
        RECT  2.850 1.360 3.090 3.790 ;
        RECT  0.720 2.130 0.960 3.790 ;
        RECT  2.850 2.950 3.410 3.190 ;
        RECT  0.690 2.080 0.930 2.480 ;
        RECT  2.850 1.360 3.410 1.600 ;
        RECT  1.570 2.870 1.970 3.110 ;
        RECT  1.650 1.570 1.890 3.110 ;
        RECT  1.650 2.190 2.090 2.590 ;
        RECT  1.570 1.570 1.970 1.810 ;
    END
END FA3

MACRO FA3P
    CLASS CORE ;
    FOREIGN FA3P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.420 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.780 1.580 11.180 1.820 ;
        RECT  11.420 3.020 11.660 4.240 ;
        RECT  12.300 1.100 12.540 1.820 ;
        RECT  12.220 1.580 12.620 1.820 ;
        RECT  12.860 3.020 13.100 4.240 ;
        RECT  10.860 1.100 13.820 1.340 ;
        RECT  13.580 1.100 13.820 2.290 ;
        RECT  13.580 2.050 14.310 2.290 ;
        RECT  14.070 2.050 14.310 4.240 ;
        RECT  18.790 3.520 19.030 4.240 ;
        RECT  11.420 4.000 19.030 4.240 ;
        RECT  21.860 2.790 22.150 3.280 ;
        RECT  21.870 1.330 22.150 3.760 ;
        RECT  18.790 3.520 22.150 3.760 ;
        RECT  21.780 1.330 23.480 1.570 ;
        RECT  21.860 3.040 23.480 3.280 ;
        RECT  10.860 1.100 11.100 1.820 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.230 3.990 7.180 4.230 ;
        RECT  6.940 3.520 7.180 4.230 ;
        RECT  6.940 3.520 10.370 3.760 ;
        RECT  10.090 3.020 10.370 4.420 ;
        RECT  10.090 3.020 10.380 3.420 ;
        RECT  3.720 4.060 4.760 4.340 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.240 1.100 1.640 ;
        RECT  0.790 2.790 1.100 3.190 ;
        RECT  0.790 1.020 1.070 3.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.980 2.240 18.430 2.640 ;
        RECT  18.150 1.420 18.430 2.640 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  18.770 1.420 19.050 2.640 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.760 -0.380 2.700 0.720 ;
        RECT  5.050 -0.380 5.450 0.560 ;
        RECT  7.420 -0.380 7.820 0.560 ;
        RECT  9.060 -0.380 9.460 0.560 ;
        RECT  14.540 -0.380 14.940 0.560 ;
        RECT  17.250 -0.380 17.650 0.700 ;
        RECT  18.320 -0.380 18.720 0.560 ;
        RECT  22.430 -0.380 22.830 0.560 ;
        RECT  23.800 -0.380 25.260 0.560 ;
        RECT  0.000 -0.380 25.420 0.380 ;
        RECT  0.160 -0.380 0.560 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.470 4.180 1.870 5.420 ;
        RECT  2.300 4.080 2.700 5.420 ;
        RECT  5.000 4.480 6.480 5.420 ;
        RECT  7.420 4.260 7.820 5.420 ;
        RECT  8.880 4.260 9.280 5.420 ;
        RECT  14.460 4.480 14.860 5.420 ;
        RECT  17.250 4.480 17.650 5.420 ;
        RECT  18.210 4.480 18.610 5.420 ;
        RECT  19.980 4.480 21.460 5.420 ;
        RECT  22.430 4.480 22.830 5.420 ;
        RECT  23.800 4.480 24.200 5.420 ;
        RECT  24.720 4.630 25.120 5.420 ;
        RECT  0.000 4.660 25.420 5.420 ;
        RECT  0.160 4.180 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  24.940 1.560 25.180 3.200 ;
        RECT  22.540 2.560 25.180 2.800 ;
        RECT  22.540 1.830 22.780 2.800 ;
        RECT  22.540 1.830 22.900 2.230 ;
        RECT  24.540 1.560 25.180 1.800 ;
        RECT  24.540 1.400 24.780 1.800 ;
        RECT  19.440 4.000 24.630 4.240 ;
        RECT  24.390 3.750 24.630 4.240 ;
        RECT  24.390 3.750 25.030 3.990 ;
        RECT  14.860 3.440 15.260 3.730 ;
        RECT  14.860 3.440 18.050 3.680 ;
        RECT  17.810 2.960 18.050 3.680 ;
        RECT  16.610 1.240 16.850 3.680 ;
        RECT  17.810 2.960 19.680 3.200 ;
        RECT  19.360 1.350 19.600 3.200 ;
        RECT  23.720 2.080 24.240 2.320 ;
        RECT  19.360 1.960 20.800 2.200 ;
        RECT  20.560 0.800 20.800 2.200 ;
        RECT  23.720 0.800 23.960 2.320 ;
        RECT  20.560 0.800 23.960 1.040 ;
        RECT  20.260 2.800 20.500 3.200 ;
        RECT  20.260 2.800 21.480 3.040 ;
        RECT  21.240 1.340 21.480 3.040 ;
        RECT  21.060 1.340 21.480 1.580 ;
        RECT  17.190 2.800 17.570 3.200 ;
        RECT  17.190 0.940 17.430 3.200 ;
        RECT  17.190 1.580 17.650 1.820 ;
        RECT  17.190 0.940 18.460 1.180 ;
        RECT  18.220 0.800 19.960 1.040 ;
        RECT  15.890 0.840 16.130 3.200 ;
        RECT  14.060 0.840 16.130 1.080 ;
        RECT  5.610 0.800 10.030 1.040 ;
        RECT  9.790 0.620 14.300 0.860 ;
        RECT  15.170 1.320 15.410 3.200 ;
        RECT  15.090 1.320 15.490 1.560 ;
        RECT  13.580 2.540 13.820 3.270 ;
        RECT  12.140 2.540 12.380 3.270 ;
        RECT  10.700 2.540 10.940 3.270 ;
        RECT  9.580 2.540 9.820 3.270 ;
        RECT  8.230 2.870 8.470 3.270 ;
        RECT  6.880 2.870 7.120 3.270 ;
        RECT  6.880 2.950 9.820 3.190 ;
        RECT  9.580 2.540 13.820 2.780 ;
        RECT  10.090 2.060 13.180 2.300 ;
        RECT  12.940 1.580 13.180 2.300 ;
        RECT  11.530 1.580 11.770 2.300 ;
        RECT  10.090 1.430 10.330 2.300 ;
        RECT  12.940 1.580 13.340 1.820 ;
        RECT  11.500 1.580 11.900 1.820 ;
        RECT  6.800 1.430 10.410 1.670 ;
        RECT  4.530 3.510 6.640 3.750 ;
        RECT  6.400 2.390 6.640 3.750 ;
        RECT  4.530 1.280 4.770 3.750 ;
        RECT  4.530 2.870 4.780 3.270 ;
        RECT  6.400 2.390 7.690 2.630 ;
        RECT  4.530 1.280 4.780 1.680 ;
        RECT  5.920 1.280 6.160 3.270 ;
        RECT  3.090 2.870 3.340 3.270 ;
        RECT  3.090 0.800 3.330 3.270 ;
        RECT  5.010 1.820 5.260 2.220 ;
        RECT  5.020 0.800 5.260 2.220 ;
        RECT  5.920 1.900 6.430 2.140 ;
        RECT  3.090 1.280 3.340 1.680 ;
        RECT  5.020 1.280 6.160 1.520 ;
        RECT  3.090 0.800 5.260 1.040 ;
        RECT  1.450 3.550 3.820 3.790 ;
        RECT  3.580 1.360 3.820 3.790 ;
        RECT  1.450 2.130 1.690 3.790 ;
        RECT  3.580 2.950 4.140 3.190 ;
        RECT  1.420 1.870 1.660 2.270 ;
        RECT  3.580 1.360 4.140 1.600 ;
        RECT  2.300 2.870 2.700 3.110 ;
        RECT  2.380 1.570 2.620 3.110 ;
        RECT  2.380 2.190 2.820 2.590 ;
        RECT  2.300 1.570 2.700 1.810 ;
    END
END FA3P

MACRO FA3S
    CLASS CORE ;
    FOREIGN FA3S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.210 2.870 7.870 3.270 ;
        RECT  7.630 1.320 7.870 4.240 ;
        RECT  11.970 3.520 12.210 4.240 ;
        RECT  7.630 4.000 12.210 4.240 ;
        RECT  14.850 1.310 15.090 3.760 ;
        RECT  14.850 1.310 15.310 1.550 ;
        RECT  14.850 2.470 15.310 3.760 ;
        RECT  11.970 3.520 15.310 3.760 ;
        RECT  7.130 1.320 7.870 1.560 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.990 4.060 4.290 4.340 ;
        RECT  6.390 1.320 6.630 2.080 ;
        RECT  6.390 1.780 6.970 2.080 ;
        RECT  3.500 4.000 6.930 4.240 ;
        RECT  6.690 1.780 6.930 4.240 ;
        RECT  6.690 1.780 6.970 2.180 ;
        RECT  3.500 3.810 3.900 4.340 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.420 0.480 1.820 ;
        RECT  0.170 2.790 0.480 3.190 ;
        RECT  0.170 0.620 0.450 3.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.220 2.240 11.610 2.640 ;
        RECT  11.330 1.420 11.610 2.640 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.290 12.410 2.530 ;
        RECT  11.950 1.420 12.230 2.640 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.670 -0.380 6.070 0.560 ;
        RECT  7.850 -0.380 8.250 0.560 ;
        RECT  10.600 -0.380 11.000 0.700 ;
        RECT  11.670 -0.380 12.070 0.560 ;
        RECT  14.850 -0.380 16.920 0.560 ;
        RECT  0.000 -0.380 17.360 0.380 ;
        RECT  0.700 -0.380 1.640 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.520 4.480 6.090 5.420 ;
        RECT  7.700 4.480 8.100 5.420 ;
        RECT  10.600 4.480 11.000 5.420 ;
        RECT  11.560 4.480 11.960 5.420 ;
        RECT  13.240 4.480 15.800 5.420 ;
        RECT  0.000 4.660 17.360 5.420 ;
        RECT  0.160 4.280 1.640 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  15.630 3.140 17.200 3.380 ;
        RECT  15.630 1.650 15.870 3.380 ;
        RECT  15.330 1.830 15.870 2.230 ;
        RECT  16.420 1.440 16.660 1.890 ;
        RECT  15.630 1.650 16.660 1.890 ;
        RECT  8.210 3.440 8.610 3.730 ;
        RECT  8.210 3.440 11.730 3.680 ;
        RECT  11.490 3.030 11.730 3.680 ;
        RECT  9.960 1.240 10.200 3.680 ;
        RECT  11.490 3.030 12.950 3.270 ;
        RECT  12.710 1.350 12.950 3.270 ;
        RECT  12.440 2.960 12.950 3.270 ;
        RECT  16.110 2.130 17.170 2.370 ;
        RECT  16.930 0.800 17.170 2.370 ;
        RECT  12.710 1.960 13.930 2.200 ;
        RECT  13.690 0.800 13.930 2.200 ;
        RECT  12.520 1.350 12.950 1.750 ;
        RECT  13.690 0.800 17.170 1.040 ;
        RECT  12.580 4.000 16.970 4.240 ;
        RECT  13.390 2.800 13.630 3.200 ;
        RECT  13.390 2.800 14.610 3.040 ;
        RECT  14.370 1.340 14.610 3.040 ;
        RECT  14.190 1.340 14.610 1.580 ;
        RECT  10.540 2.800 10.920 3.200 ;
        RECT  10.540 0.940 10.780 3.200 ;
        RECT  10.540 1.580 11.000 1.820 ;
        RECT  10.540 0.940 11.810 1.180 ;
        RECT  11.570 0.800 13.090 1.040 ;
        RECT  9.240 0.840 9.480 3.200 ;
        RECT  6.520 0.840 9.480 1.080 ;
        RECT  4.880 0.800 6.760 1.040 ;
        RECT  8.520 1.320 8.760 3.200 ;
        RECT  8.440 1.320 8.840 1.560 ;
        RECT  4.140 3.450 6.300 3.690 ;
        RECT  6.060 2.330 6.300 3.690 ;
        RECT  3.780 3.230 4.380 3.470 ;
        RECT  3.780 2.830 4.050 3.470 ;
        RECT  3.780 1.280 4.020 3.470 ;
        RECT  6.060 2.330 6.310 2.730 ;
        RECT  3.780 1.280 4.050 1.680 ;
        RECT  2.370 0.800 2.610 3.230 ;
        RECT  5.110 2.870 5.620 3.110 ;
        RECT  5.380 1.280 5.620 3.110 ;
        RECT  4.280 1.820 4.520 2.220 ;
        RECT  4.280 1.820 5.620 2.060 ;
        RECT  5.230 1.280 5.620 2.060 ;
        RECT  4.290 0.800 4.530 2.060 ;
        RECT  2.370 0.800 4.530 1.040 ;
        RECT  0.720 3.550 3.090 3.790 ;
        RECT  2.850 1.360 3.090 3.790 ;
        RECT  0.720 2.130 0.960 3.790 ;
        RECT  2.850 2.910 3.410 3.150 ;
        RECT  0.690 2.080 0.930 2.480 ;
        RECT  2.850 1.360 3.410 1.600 ;
        RECT  1.570 2.870 1.970 3.110 ;
        RECT  1.650 1.500 1.890 3.110 ;
        RECT  1.650 2.190 2.080 2.590 ;
        RECT  1.570 1.500 1.970 1.740 ;
    END
END FA3S

MACRO FACS1
    CLASS CORE ;
    FOREIGN FACS1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 50.220 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.210 2.080 7.160 2.320 ;
        RECT  6.920 2.050 8.340 2.290 ;
        RECT  9.660 1.200 9.900 2.320 ;
        RECT  8.100 2.080 9.900 2.320 ;
        RECT  9.660 1.200 13.160 1.440 ;
        RECT  12.920 1.200 13.160 2.080 ;
        RECT  14.010 1.920 14.650 2.160 ;
        RECT  12.920 1.840 14.250 2.080 ;
        RECT  14.250 1.920 14.650 2.220 ;
        RECT  6.210 2.080 6.610 2.380 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  35.730 1.840 37.200 2.080 ;
        RECT  36.960 1.200 37.200 2.080 ;
        RECT  36.960 1.200 40.450 1.440 ;
        RECT  40.210 1.200 40.450 2.300 ;
        RECT  40.210 2.060 41.430 2.300 ;
        RECT  41.190 2.050 43.150 2.290 ;
        RECT  42.910 2.120 43.920 2.360 ;
        RECT  35.420 1.980 35.970 2.220 ;
        END
    END CI0
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.010 1.300 2.290 1.700 ;
        RECT  2.010 2.800 2.360 3.200 ;
        RECT  4.360 1.100 4.600 2.550 ;
        RECT  4.530 2.310 4.770 3.940 ;
        RECT  2.010 3.520 4.770 3.760 ;
        RECT  4.360 1.100 5.960 1.340 ;
        RECT  5.850 3.100 6.090 3.940 ;
        RECT  4.530 3.700 6.090 3.940 ;
        RECT  5.770 3.100 6.170 3.340 ;
        RECT  2.010 1.300 2.250 3.760 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  43.960 3.100 44.360 3.340 ;
        RECT  44.190 1.100 45.800 1.340 ;
        RECT  45.450 2.520 45.690 3.940 ;
        RECT  44.040 3.700 45.690 3.940 ;
        RECT  45.560 1.100 45.800 2.760 ;
        RECT  47.870 1.300 48.240 1.700 ;
        RECT  47.850 2.800 48.240 3.200 ;
        RECT  45.450 3.520 48.240 3.760 ;
        RECT  48.000 1.300 48.240 3.760 ;
        RECT  44.040 3.100 44.280 3.940 ;
        END
    END CO0
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  23.130 1.500 23.370 3.280 ;
        RECT  22.930 3.040 23.370 3.280 ;
        RECT  23.030 1.500 23.370 1.900 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 1.800 0.480 2.200 ;
        RECT  0.190 4.000 4.070 4.240 ;
        RECT  6.850 3.580 7.090 4.420 ;
        RECT  3.830 4.180 7.090 4.420 ;
        RECT  6.850 3.580 9.670 3.820 ;
        RECT  9.430 3.580 9.670 4.420 ;
        RECT  9.430 4.180 10.750 4.420 ;
        RECT  10.510 4.000 16.250 4.240 ;
        RECT  16.010 4.180 19.030 4.420 ;
        RECT  18.790 4.000 20.150 4.240 ;
        RECT  21.140 4.080 21.540 4.420 ;
        RECT  19.910 4.180 22.620 4.420 ;
        RECT  22.380 4.000 25.590 4.240 ;
        RECT  27.170 4.080 27.570 4.420 ;
        RECT  25.350 4.180 30.120 4.420 ;
        RECT  29.880 4.000 31.350 4.240 ;
        RECT  31.110 4.180 34.020 4.420 ;
        RECT  33.780 4.000 39.610 4.240 ;
        RECT  40.460 3.580 40.700 4.420 ;
        RECT  39.370 4.180 40.700 4.420 ;
        RECT  40.460 3.580 43.460 3.820 ;
        RECT  43.220 3.580 43.460 4.420 ;
        RECT  43.220 4.180 46.400 4.420 ;
        RECT  46.160 4.000 50.030 4.240 ;
        RECT  49.790 2.290 50.030 4.240 ;
        RECT  49.660 2.520 50.060 2.760 ;
        RECT  0.190 1.800 0.430 4.240 ;
        END
    END B
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  24.350 2.060 24.630 2.800 ;
        RECT  24.290 2.060 24.630 2.460 ;
        END
    END CS
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.740 2.520 1.140 2.760 ;
        RECT  0.770 0.800 4.120 1.040 ;
        RECT  3.880 0.620 4.120 2.310 ;
        RECT  3.090 2.070 4.120 2.310 ;
        RECT  3.880 0.620 6.780 0.860 ;
        RECT  6.540 0.800 9.340 1.040 ;
        RECT  9.100 0.720 13.640 0.960 ;
        RECT  14.360 0.620 14.600 1.200 ;
        RECT  13.400 0.960 14.600 1.200 ;
        RECT  14.360 0.620 18.250 0.860 ;
        RECT  18.010 0.620 18.250 1.250 ;
        RECT  18.970 0.620 19.210 1.250 ;
        RECT  18.010 1.010 19.210 1.250 ;
        RECT  18.970 0.620 22.020 0.860 ;
        RECT  21.780 0.620 22.020 1.130 ;
        RECT  22.900 0.620 23.140 1.130 ;
        RECT  21.780 0.890 23.140 1.130 ;
        RECT  22.900 0.620 26.830 0.860 ;
        RECT  26.590 0.620 26.830 1.130 ;
        RECT  27.880 0.620 28.120 1.130 ;
        RECT  26.590 0.890 28.120 1.130 ;
        RECT  27.880 0.620 32.180 0.860 ;
        RECT  31.940 0.720 35.670 0.960 ;
        RECT  35.430 0.960 36.630 1.200 ;
        RECT  36.390 0.720 40.930 0.960 ;
        RECT  40.690 0.800 43.590 1.040 ;
        RECT  46.040 0.620 46.280 2.300 ;
        RECT  43.350 0.620 46.310 0.860 ;
        RECT  46.040 2.060 47.070 2.300 ;
        RECT  46.040 0.800 49.430 1.040 ;
        RECT  49.150 0.800 49.430 2.280 ;
        RECT  49.080 1.880 49.480 2.120 ;
        RECT  0.770 0.800 1.010 2.760 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.760 -0.380 3.160 0.560 ;
        RECT  7.020 -0.380 7.420 0.560 ;
        RECT  8.480 -0.380 8.880 0.560 ;
        RECT  13.880 -0.380 14.120 0.640 ;
        RECT  18.490 -0.380 18.730 0.640 ;
        RECT  22.310 -0.380 22.550 0.650 ;
        RECT  27.070 -0.380 27.310 0.650 ;
        RECT  35.910 -0.380 36.150 0.640 ;
        RECT  41.250 -0.380 41.650 0.560 ;
        RECT  42.710 -0.380 43.110 0.560 ;
        RECT  47.000 -0.380 47.400 0.560 ;
        RECT  48.600 -0.380 49.000 0.560 ;
        RECT  0.000 -0.380 50.220 0.380 ;
        RECT  1.230 -0.380 1.630 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.850 4.480 3.250 5.420 ;
        RECT  7.330 4.180 7.730 5.420 ;
        RECT  8.790 4.180 9.190 5.420 ;
        RECT  10.990 4.480 11.390 5.420 ;
        RECT  13.070 4.480 13.470 5.420 ;
        RECT  15.370 4.480 15.770 5.420 ;
        RECT  19.270 4.480 19.670 5.420 ;
        RECT  23.940 4.480 24.880 5.420 ;
        RECT  30.470 4.480 30.870 5.420 ;
        RECT  34.290 4.480 34.690 5.420 ;
        RECT  36.560 4.480 36.960 5.420 ;
        RECT  38.730 4.480 39.130 5.420 ;
        RECT  40.940 4.180 41.340 5.420 ;
        RECT  42.400 4.180 42.800 5.420 ;
        RECT  46.970 4.480 47.370 5.420 ;
        RECT  48.500 4.480 49.780 5.420 ;
        RECT  0.000 4.660 50.220 5.420 ;
        RECT  0.440 4.480 1.720 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  48.590 3.060 49.550 3.300 ;
        RECT  48.590 1.340 48.830 3.300 ;
        RECT  48.480 1.860 48.830 2.260 ;
        RECT  48.510 1.340 48.910 1.580 ;
        RECT  45.930 3.030 47.610 3.270 ;
        RECT  47.370 1.580 47.610 3.270 ;
        RECT  47.370 1.840 47.670 2.240 ;
        RECT  46.520 1.580 47.610 1.820 ;
        RECT  46.520 1.300 46.760 1.820 ;
        RECT  45.000 1.580 45.240 1.980 ;
        RECT  43.330 1.580 45.240 1.820 ;
        RECT  40.690 1.420 40.930 1.820 ;
        RECT  40.690 1.570 43.570 1.810 ;
        RECT  44.680 3.100 45.130 3.340 ;
        RECT  44.890 2.620 45.130 3.340 ;
        RECT  40.320 3.100 43.640 3.340 ;
        RECT  43.400 2.620 43.640 3.340 ;
        RECT  43.400 2.620 45.130 2.860 ;
        RECT  39.570 2.980 39.970 3.220 ;
        RECT  39.730 1.680 39.970 3.220 ;
        RECT  39.730 2.540 42.670 2.780 ;
        RECT  42.270 2.530 42.670 2.780 ;
        RECT  39.570 1.680 39.970 1.920 ;
        RECT  39.850 3.520 40.090 3.920 ;
        RECT  38.320 3.520 40.090 3.760 ;
        RECT  38.320 1.680 38.560 3.760 ;
        RECT  38.160 2.980 38.560 3.220 ;
        RECT  38.160 1.680 38.560 1.920 ;
        RECT  33.650 3.520 37.760 3.760 ;
        RECT  37.520 1.680 37.760 3.760 ;
        RECT  33.650 1.680 33.890 3.760 ;
        RECT  37.440 2.980 37.840 3.220 ;
        RECT  36.100 2.440 37.760 2.680 ;
        RECT  37.440 1.680 37.840 1.920 ;
        RECT  33.570 1.680 33.970 1.920 ;
        RECT  32.130 3.220 32.610 3.460 ;
        RECT  32.370 1.200 32.610 3.460 ;
        RECT  34.940 2.980 35.530 3.220 ;
        RECT  34.940 1.200 35.180 3.220 ;
        RECT  32.130 1.680 32.610 1.920 ;
        RECT  34.940 1.440 35.530 1.680 ;
        RECT  32.370 1.200 35.180 1.440 ;
        RECT  34.290 3.040 34.690 3.280 ;
        RECT  34.340 1.680 34.580 3.280 ;
        RECT  34.230 2.240 34.580 2.640 ;
        RECT  34.290 1.680 34.690 1.920 ;
        RECT  31.590 3.700 33.170 3.940 ;
        RECT  32.930 1.680 33.170 3.940 ;
        RECT  30.500 3.520 31.830 3.760 ;
        RECT  30.500 2.710 30.740 3.760 ;
        RECT  32.850 3.220 33.250 3.460 ;
        RECT  30.440 2.710 30.740 3.110 ;
        RECT  32.850 1.680 33.250 1.920 ;
        RECT  28.430 3.120 28.830 3.360 ;
        RECT  31.410 3.040 31.810 3.280 ;
        RECT  28.510 1.100 28.750 3.360 ;
        RECT  31.460 1.490 31.700 3.280 ;
        RECT  30.510 1.490 31.700 1.730 ;
        RECT  30.510 1.100 30.750 1.730 ;
        RECT  28.510 1.100 30.750 1.340 ;
        RECT  29.940 3.360 30.260 3.760 ;
        RECT  29.940 1.580 30.180 3.760 ;
        RECT  30.980 2.040 31.220 2.440 ;
        RECT  29.940 2.120 31.220 2.360 ;
        RECT  29.870 1.580 30.270 1.820 ;
        RECT  26.950 3.600 29.470 3.840 ;
        RECT  29.230 1.580 29.470 3.840 ;
        RECT  26.950 1.500 27.190 3.840 ;
        RECT  29.150 1.580 29.550 1.820 ;
        RECT  27.690 2.880 28.110 3.120 ;
        RECT  27.690 1.580 27.930 3.120 ;
        RECT  27.690 2.140 28.170 2.540 ;
        RECT  27.690 1.580 28.110 1.820 ;
        RECT  26.110 3.040 26.470 3.440 ;
        RECT  26.110 1.100 26.350 3.440 ;
        RECT  23.610 2.310 23.870 2.710 ;
        RECT  23.630 1.100 23.870 2.710 ;
        RECT  26.110 1.500 26.470 1.900 ;
        RECT  23.630 1.100 26.350 1.340 ;
        RECT  20.810 3.600 22.200 3.840 ;
        RECT  25.630 1.580 25.870 3.760 ;
        RECT  21.960 3.520 25.870 3.760 ;
        RECT  25.510 3.040 25.870 3.760 ;
        RECT  20.810 1.580 21.050 3.840 ;
        RECT  20.730 3.040 21.050 3.440 ;
        RECT  25.430 1.580 25.870 1.820 ;
        RECT  20.650 1.580 21.050 1.820 ;
        RECT  24.510 3.040 25.110 3.280 ;
        RECT  24.870 1.580 25.110 3.280 ;
        RECT  24.870 2.320 25.210 2.720 ;
        RECT  24.510 1.580 25.110 1.820 ;
        RECT  22.090 2.970 22.490 3.210 ;
        RECT  22.150 1.580 22.390 3.210 ;
        RECT  21.960 2.330 22.390 2.730 ;
        RECT  22.090 1.580 22.490 1.820 ;
        RECT  21.370 3.120 21.770 3.360 ;
        RECT  18.190 3.040 18.740 3.280 ;
        RECT  21.450 1.500 21.690 3.360 ;
        RECT  18.190 1.490 18.430 3.280 ;
        RECT  21.290 1.100 21.530 1.920 ;
        RECT  18.190 1.490 18.580 1.900 ;
        RECT  18.190 1.490 19.690 1.730 ;
        RECT  19.450 1.100 19.690 1.730 ;
        RECT  19.450 1.100 21.530 1.340 ;
        RECT  19.860 3.520 20.260 3.760 ;
        RECT  20.020 1.580 20.260 3.760 ;
        RECT  18.960 2.040 19.200 2.440 ;
        RECT  18.960 2.040 20.260 2.280 ;
        RECT  19.930 1.580 20.260 2.280 ;
        RECT  19.930 1.580 20.330 1.820 ;
        RECT  16.890 3.700 18.550 3.940 ;
        RECT  19.380 2.710 19.620 3.760 ;
        RECT  18.310 3.520 19.620 3.760 ;
        RECT  16.890 1.680 17.130 3.940 ;
        RECT  16.810 3.220 17.210 3.460 ;
        RECT  19.380 2.710 19.710 3.110 ;
        RECT  16.810 1.680 17.210 1.920 ;
        RECT  17.530 3.220 17.930 3.460 ;
        RECT  14.530 2.980 15.130 3.220 ;
        RECT  14.890 1.200 15.130 3.220 ;
        RECT  17.530 1.200 17.770 3.460 ;
        RECT  17.530 1.680 17.930 1.920 ;
        RECT  14.530 1.440 15.130 1.680 ;
        RECT  14.890 1.200 17.770 1.440 ;
        RECT  12.300 3.520 16.410 3.760 ;
        RECT  16.170 1.680 16.410 3.760 ;
        RECT  12.300 2.980 12.540 3.760 ;
        RECT  12.280 2.980 12.680 3.220 ;
        RECT  12.290 1.680 12.530 3.220 ;
        RECT  12.290 2.440 13.940 2.680 ;
        RECT  16.090 1.680 16.490 1.920 ;
        RECT  12.280 1.680 12.680 1.920 ;
        RECT  15.370 3.040 15.770 3.280 ;
        RECT  15.450 1.680 15.690 3.280 ;
        RECT  15.450 2.240 15.830 2.640 ;
        RECT  15.370 1.680 15.770 1.920 ;
        RECT  10.030 3.460 10.270 3.860 ;
        RECT  10.030 3.520 11.800 3.760 ;
        RECT  11.560 1.680 11.800 3.760 ;
        RECT  11.560 2.980 11.960 3.220 ;
        RECT  11.560 1.680 11.960 1.920 ;
        RECT  10.140 2.980 10.540 3.220 ;
        RECT  10.140 1.680 10.380 3.220 ;
        RECT  7.460 2.560 10.380 2.800 ;
        RECT  7.460 2.530 7.860 2.800 ;
        RECT  10.140 1.680 10.540 1.920 ;
        RECT  6.490 3.100 9.810 3.340 ;
        RECT  5.050 3.100 5.450 3.340 ;
        RECT  6.490 2.620 6.730 3.340 ;
        RECT  5.050 2.620 5.290 3.340 ;
        RECT  5.050 2.620 6.730 2.860 ;
        RECT  9.180 1.440 9.420 1.840 ;
        RECT  4.840 1.600 6.680 1.840 ;
        RECT  6.440 1.570 9.420 1.810 ;
        RECT  2.600 3.030 4.280 3.270 ;
        RECT  2.600 1.380 2.840 3.270 ;
        RECT  2.490 1.840 2.840 2.240 ;
        RECT  3.400 1.300 3.640 1.700 ;
        RECT  2.600 1.380 3.640 1.620 ;
        RECT  0.670 3.060 1.770 3.300 ;
        RECT  1.530 1.340 1.770 3.300 ;
        RECT  1.250 1.340 1.770 1.580 ;
    END
END FACS1

MACRO FACS1P
    CLASS CORE ;
    FOREIGN FACS1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.620 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.090 2.050 14.680 2.290 ;
        RECT  15.380 1.200 15.620 2.320 ;
        RECT  14.440 2.080 15.620 2.320 ;
        RECT  15.380 1.200 18.880 1.440 ;
        RECT  18.640 1.200 18.880 2.080 ;
        RECT  18.640 1.840 19.860 2.080 ;
        RECT  19.620 1.980 20.370 2.160 ;
        RECT  18.640 1.920 20.260 2.080 ;
        RECT  19.970 1.980 20.370 2.220 ;
        RECT  8.650 2.140 11.330 2.380 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  42.350 1.840 43.760 2.080 ;
        RECT  43.520 1.200 43.760 2.080 ;
        RECT  43.520 1.200 47.020 1.440 ;
        RECT  46.780 1.200 47.020 2.380 ;
        RECT  46.780 2.140 48.050 2.380 ;
        RECT  47.810 2.050 51.440 2.290 ;
        RECT  51.200 2.120 53.880 2.360 ;
        RECT  53.480 2.120 53.880 2.380 ;
        RECT  41.980 1.980 42.590 2.220 ;
        END
    END CI0
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.170 2.800 2.410 3.200 ;
        RECT  2.670 1.360 2.910 3.760 ;
        RECT  2.170 2.880 3.650 3.120 ;
        RECT  2.050 1.440 3.670 1.680 ;
        RECT  3.410 2.800 3.650 3.200 ;
        RECT  3.430 1.360 3.670 1.760 ;
        RECT  5.700 1.100 5.940 2.550 ;
        RECT  5.860 2.310 6.100 3.940 ;
        RECT  2.670 3.520 6.100 3.760 ;
        RECT  7.060 3.100 7.300 3.940 ;
        RECT  6.980 3.100 7.380 3.340 ;
        RECT  8.500 3.100 8.740 3.940 ;
        RECT  5.860 3.700 8.740 3.940 ;
        RECT  5.700 1.100 8.770 1.340 ;
        RECT  8.420 3.100 8.820 3.340 ;
        RECT  2.050 1.360 2.290 1.760 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  53.710 3.100 54.110 3.340 ;
        RECT  55.230 3.100 55.470 3.940 ;
        RECT  55.150 3.100 55.550 3.340 ;
        RECT  53.640 1.100 56.700 1.340 ;
        RECT  56.430 2.520 56.670 3.940 ;
        RECT  53.790 3.700 56.670 3.940 ;
        RECT  56.460 1.100 56.700 2.760 ;
        RECT  58.890 1.360 59.130 1.760 ;
        RECT  58.910 2.800 59.150 3.200 ;
        RECT  56.430 3.520 59.950 3.760 ;
        RECT  59.710 1.440 59.950 3.760 ;
        RECT  58.890 1.440 60.510 1.680 ;
        RECT  58.910 2.880 60.470 3.120 ;
        RECT  60.270 1.360 60.510 1.760 ;
        RECT  53.790 3.100 54.030 3.940 ;
        END
    END CO0
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  29.330 1.500 29.830 1.900 ;
        RECT  29.330 3.040 29.890 3.280 ;
        RECT  29.330 1.500 29.570 3.280 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 1.800 0.480 2.200 ;
        RECT  0.190 4.000 5.410 4.240 ;
        RECT  9.380 3.580 9.620 4.420 ;
        RECT  5.170 4.180 9.620 4.420 ;
        RECT  9.380 3.580 15.500 3.820 ;
        RECT  15.260 3.580 15.500 4.420 ;
        RECT  15.260 4.180 16.470 4.420 ;
        RECT  16.230 4.000 21.970 4.240 ;
        RECT  21.730 4.180 24.750 4.420 ;
        RECT  24.510 4.000 25.870 4.240 ;
        RECT  26.860 4.080 27.260 4.420 ;
        RECT  25.630 4.180 28.340 4.420 ;
        RECT  28.100 4.000 32.150 4.240 ;
        RECT  33.730 4.080 34.130 4.420 ;
        RECT  31.910 4.180 36.680 4.420 ;
        RECT  36.440 4.000 37.910 4.240 ;
        RECT  37.670 4.180 40.580 4.420 ;
        RECT  40.340 4.000 46.170 4.240 ;
        RECT  46.890 3.580 47.130 4.420 ;
        RECT  45.930 4.180 47.130 4.420 ;
        RECT  46.890 3.580 53.270 3.820 ;
        RECT  53.030 3.580 53.270 4.420 ;
        RECT  53.030 4.180 57.460 4.420 ;
        RECT  57.220 4.000 62.430 4.240 ;
        RECT  62.190 2.290 62.430 4.240 ;
        RECT  62.060 2.520 62.460 2.760 ;
        RECT  0.190 1.800 0.430 4.240 ;
        END
    END B
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  30.550 2.060 31.070 2.460 ;
        RECT  30.550 2.060 30.830 2.800 ;
        END
    END CS
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.740 2.520 1.140 2.760 ;
        RECT  0.770 0.800 5.460 1.040 ;
        RECT  5.220 0.620 5.460 2.310 ;
        RECT  4.430 2.070 5.460 2.310 ;
        RECT  5.220 0.620 9.560 0.860 ;
        RECT  9.320 0.800 15.170 1.040 ;
        RECT  14.930 0.720 19.360 0.960 ;
        RECT  20.080 0.620 20.320 1.200 ;
        RECT  19.120 0.960 20.320 1.200 ;
        RECT  20.080 0.620 23.970 0.860 ;
        RECT  23.730 0.620 23.970 1.250 ;
        RECT  24.690 0.620 24.930 1.250 ;
        RECT  23.730 1.010 24.930 1.250 ;
        RECT  24.690 0.620 27.740 0.860 ;
        RECT  27.500 0.620 27.740 1.130 ;
        RECT  29.460 0.620 29.700 1.130 ;
        RECT  27.500 0.890 29.700 1.130 ;
        RECT  29.460 0.620 33.390 0.860 ;
        RECT  33.150 0.620 33.390 1.130 ;
        RECT  34.440 0.620 34.680 1.130 ;
        RECT  33.150 0.890 34.680 1.130 ;
        RECT  34.440 0.620 38.740 0.860 ;
        RECT  38.500 0.720 42.230 0.960 ;
        RECT  41.990 0.960 43.190 1.200 ;
        RECT  42.950 0.720 47.590 0.960 ;
        RECT  47.350 0.800 53.330 1.040 ;
        RECT  53.090 0.620 57.260 0.860 ;
        RECT  57.020 0.620 57.260 2.300 ;
        RECT  57.020 2.060 58.050 2.300 ;
        RECT  57.020 0.800 61.830 1.040 ;
        RECT  61.550 0.800 61.830 2.280 ;
        RECT  61.480 1.880 61.880 2.120 ;
        RECT  0.770 0.800 1.010 2.760 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.070 -0.380 4.470 0.560 ;
        RECT  9.820 -0.380 10.220 0.560 ;
        RECT  11.280 -0.380 11.680 0.560 ;
        RECT  12.740 -0.380 13.140 0.560 ;
        RECT  14.200 -0.380 14.600 0.560 ;
        RECT  19.600 -0.380 19.840 0.640 ;
        RECT  24.210 -0.380 24.450 0.640 ;
        RECT  27.980 -0.380 28.970 0.650 ;
        RECT  33.630 -0.380 33.870 0.650 ;
        RECT  42.470 -0.380 42.710 0.640 ;
        RECT  47.800 -0.380 48.200 0.560 ;
        RECT  49.260 -0.380 49.660 0.560 ;
        RECT  50.720 -0.380 51.120 0.560 ;
        RECT  52.180 -0.380 52.580 0.560 ;
        RECT  58.090 -0.380 58.490 0.560 ;
        RECT  61.000 -0.380 61.400 0.560 ;
        RECT  0.000 -0.380 62.620 0.380 ;
        RECT  1.230 -0.380 1.630 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.750 4.480 3.150 5.420 ;
        RECT  4.090 4.480 4.490 5.420 ;
        RECT  9.980 4.180 10.380 5.420 ;
        RECT  11.440 4.180 11.840 5.420 ;
        RECT  12.900 4.180 13.300 5.420 ;
        RECT  14.360 4.180 14.760 5.420 ;
        RECT  16.710 4.480 17.110 5.420 ;
        RECT  18.790 4.480 19.190 5.420 ;
        RECT  21.090 4.480 21.490 5.420 ;
        RECT  24.990 4.480 25.390 5.420 ;
        RECT  30.500 4.480 31.440 5.420 ;
        RECT  37.030 4.480 37.430 5.420 ;
        RECT  40.850 4.480 41.250 5.420 ;
        RECT  43.120 4.480 43.520 5.420 ;
        RECT  45.290 4.480 45.690 5.420 ;
        RECT  47.770 4.180 48.170 5.420 ;
        RECT  49.230 4.180 49.630 5.420 ;
        RECT  50.690 4.180 51.090 5.420 ;
        RECT  52.150 4.180 52.550 5.420 ;
        RECT  58.110 4.480 58.510 5.420 ;
        RECT  59.410 4.480 59.810 5.420 ;
        RECT  60.900 4.480 62.180 5.420 ;
        RECT  0.000 4.660 62.620 5.420 ;
        RECT  0.440 4.480 1.720 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  60.990 3.060 61.950 3.300 ;
        RECT  60.990 1.340 61.230 3.300 ;
        RECT  60.880 1.920 61.230 2.320 ;
        RECT  60.910 1.340 61.310 1.580 ;
        RECT  56.990 3.030 58.650 3.270 ;
        RECT  58.410 1.580 58.650 3.270 ;
        RECT  58.410 1.900 58.680 2.300 ;
        RECT  57.500 1.580 58.650 1.820 ;
        RECT  57.500 1.300 57.740 1.820 ;
        RECT  47.260 1.500 47.500 1.900 ;
        RECT  52.800 1.600 56.220 1.840 ;
        RECT  47.260 1.570 53.040 1.810 ;
        RECT  55.950 2.620 56.190 3.420 ;
        RECT  54.430 3.100 54.830 3.340 ;
        RECT  47.150 3.100 53.280 3.340 ;
        RECT  53.040 2.620 53.280 3.340 ;
        RECT  54.510 2.620 54.750 3.340 ;
        RECT  53.040 2.620 56.190 2.860 ;
        RECT  46.140 2.980 46.540 3.220 ;
        RECT  46.300 1.680 46.540 3.220 ;
        RECT  46.300 2.620 50.960 2.860 ;
        RECT  50.560 2.530 50.960 2.860 ;
        RECT  46.140 1.680 46.540 1.920 ;
        RECT  46.410 3.520 46.650 3.920 ;
        RECT  44.880 3.520 46.650 3.760 ;
        RECT  44.880 1.680 45.120 3.760 ;
        RECT  44.720 2.980 45.120 3.220 ;
        RECT  44.720 1.680 45.120 1.920 ;
        RECT  40.210 3.520 44.320 3.760 ;
        RECT  44.080 1.680 44.320 3.760 ;
        RECT  40.210 1.680 40.450 3.760 ;
        RECT  44.000 2.980 44.400 3.220 ;
        RECT  42.840 2.440 44.320 2.680 ;
        RECT  44.000 1.680 44.400 1.920 ;
        RECT  40.130 1.680 40.530 1.920 ;
        RECT  38.690 3.220 39.170 3.460 ;
        RECT  38.930 1.200 39.170 3.460 ;
        RECT  41.500 2.980 42.090 3.220 ;
        RECT  41.500 1.200 41.740 3.220 ;
        RECT  38.690 1.680 39.170 1.920 ;
        RECT  41.500 1.440 42.090 1.680 ;
        RECT  38.930 1.200 41.740 1.440 ;
        RECT  40.850 3.040 41.250 3.280 ;
        RECT  40.900 1.680 41.140 3.280 ;
        RECT  40.790 2.240 41.140 2.640 ;
        RECT  40.850 1.680 41.250 1.920 ;
        RECT  38.150 3.700 39.730 3.940 ;
        RECT  39.490 1.680 39.730 3.940 ;
        RECT  37.060 3.520 38.390 3.760 ;
        RECT  37.060 2.710 37.300 3.760 ;
        RECT  39.410 3.220 39.810 3.460 ;
        RECT  37.000 2.710 37.300 3.110 ;
        RECT  39.410 1.680 39.810 1.920 ;
        RECT  34.990 3.120 35.390 3.360 ;
        RECT  37.970 3.040 38.370 3.280 ;
        RECT  35.070 1.100 35.310 3.360 ;
        RECT  38.020 1.490 38.260 3.280 ;
        RECT  37.070 1.490 38.260 1.730 ;
        RECT  37.070 1.100 37.310 1.730 ;
        RECT  35.070 1.100 37.310 1.340 ;
        RECT  36.500 3.360 36.820 3.760 ;
        RECT  36.500 1.580 36.740 3.760 ;
        RECT  37.540 2.040 37.780 2.440 ;
        RECT  36.500 2.120 37.780 2.360 ;
        RECT  36.430 1.580 36.830 1.820 ;
        RECT  33.510 3.600 36.030 3.840 ;
        RECT  35.790 1.580 36.030 3.840 ;
        RECT  33.510 1.500 33.750 3.840 ;
        RECT  35.710 1.580 36.110 1.820 ;
        RECT  34.250 2.880 34.670 3.120 ;
        RECT  34.250 1.580 34.490 3.120 ;
        RECT  34.250 2.140 34.730 2.540 ;
        RECT  34.250 1.580 34.670 1.820 ;
        RECT  32.670 3.040 33.030 3.440 ;
        RECT  32.670 1.100 32.910 3.440 ;
        RECT  29.970 2.310 30.310 2.710 ;
        RECT  30.070 1.100 30.310 2.710 ;
        RECT  32.670 1.500 33.030 1.900 ;
        RECT  30.070 1.100 32.910 1.340 ;
        RECT  26.530 3.600 27.920 3.840 ;
        RECT  32.190 1.580 32.430 3.760 ;
        RECT  27.680 3.520 32.430 3.760 ;
        RECT  32.070 3.040 32.430 3.760 ;
        RECT  26.530 1.580 26.770 3.840 ;
        RECT  26.450 3.040 26.770 3.440 ;
        RECT  31.990 1.580 32.430 1.820 ;
        RECT  26.370 1.580 26.770 1.820 ;
        RECT  31.070 3.040 31.670 3.280 ;
        RECT  31.430 1.580 31.670 3.280 ;
        RECT  31.430 2.320 31.770 2.720 ;
        RECT  31.070 1.580 31.670 1.820 ;
        RECT  27.810 2.970 28.210 3.210 ;
        RECT  27.870 1.580 28.110 3.210 ;
        RECT  27.680 2.330 28.110 2.730 ;
        RECT  27.810 1.580 28.210 1.820 ;
        RECT  27.090 3.120 27.490 3.360 ;
        RECT  23.910 3.040 24.460 3.280 ;
        RECT  27.170 1.500 27.410 3.360 ;
        RECT  23.910 1.490 24.150 3.280 ;
        RECT  27.010 1.100 27.250 1.920 ;
        RECT  23.910 1.490 24.300 1.900 ;
        RECT  23.910 1.490 25.410 1.730 ;
        RECT  25.170 1.100 25.410 1.730 ;
        RECT  25.170 1.100 27.250 1.340 ;
        RECT  25.580 3.520 25.980 3.760 ;
        RECT  25.740 1.580 25.980 3.760 ;
        RECT  24.680 2.040 24.920 2.440 ;
        RECT  24.680 2.040 25.980 2.280 ;
        RECT  25.650 1.580 25.980 2.280 ;
        RECT  25.650 1.580 26.050 1.820 ;
        RECT  22.610 3.700 24.270 3.940 ;
        RECT  25.100 2.710 25.340 3.760 ;
        RECT  24.030 3.520 25.340 3.760 ;
        RECT  22.610 1.680 22.850 3.940 ;
        RECT  22.530 3.220 22.930 3.460 ;
        RECT  25.100 2.710 25.430 3.110 ;
        RECT  22.530 1.680 22.930 1.920 ;
        RECT  23.250 3.220 23.650 3.460 ;
        RECT  20.250 2.980 20.850 3.220 ;
        RECT  20.610 1.200 20.850 3.220 ;
        RECT  23.250 1.200 23.490 3.460 ;
        RECT  23.250 1.680 23.650 1.920 ;
        RECT  20.250 1.440 20.850 1.680 ;
        RECT  20.610 1.200 23.490 1.440 ;
        RECT  18.020 3.520 22.130 3.760 ;
        RECT  21.890 1.680 22.130 3.760 ;
        RECT  18.020 2.980 18.260 3.760 ;
        RECT  18.000 2.980 18.400 3.220 ;
        RECT  18.010 1.680 18.250 3.220 ;
        RECT  18.010 2.440 19.660 2.680 ;
        RECT  21.810 1.680 22.210 1.920 ;
        RECT  18.000 1.680 18.400 1.920 ;
        RECT  21.090 3.040 21.490 3.280 ;
        RECT  21.170 1.680 21.410 3.280 ;
        RECT  21.170 2.240 21.550 2.640 ;
        RECT  21.090 1.680 21.490 1.920 ;
        RECT  15.750 3.460 15.990 3.860 ;
        RECT  15.750 3.520 17.520 3.760 ;
        RECT  17.280 1.680 17.520 3.760 ;
        RECT  17.280 2.980 17.680 3.220 ;
        RECT  17.280 1.680 17.680 1.920 ;
        RECT  15.860 2.980 16.260 3.220 ;
        RECT  15.860 1.680 16.100 3.220 ;
        RECT  11.570 2.560 16.100 2.800 ;
        RECT  11.570 2.530 11.970 2.800 ;
        RECT  15.860 1.680 16.260 1.920 ;
        RECT  6.340 2.620 6.580 3.420 ;
        RECT  9.250 3.100 15.380 3.340 ;
        RECT  7.700 3.100 8.100 3.340 ;
        RECT  9.250 2.620 9.490 3.340 ;
        RECT  7.780 2.620 8.020 3.340 ;
        RECT  6.340 2.620 9.490 2.860 ;
        RECT  14.900 1.440 15.140 1.840 ;
        RECT  6.180 1.600 9.660 1.840 ;
        RECT  9.140 1.570 15.140 1.810 ;
        RECT  3.940 3.030 5.620 3.270 ;
        RECT  3.940 1.380 4.180 3.270 ;
        RECT  3.830 1.960 4.180 2.360 ;
        RECT  4.740 1.300 4.980 1.700 ;
        RECT  3.940 1.380 4.980 1.620 ;
        RECT  0.670 3.060 1.770 3.300 ;
        RECT  1.530 1.340 1.770 3.300 ;
        RECT  1.250 1.340 1.770 1.580 ;
    END
END FACS1P

MACRO FACS1S
    CLASS CORE ;
    FOREIGN FACS1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 45.260 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 1.200 7.540 2.320 ;
        RECT  5.120 2.080 7.540 2.320 ;
        RECT  7.300 1.200 10.800 1.440 ;
        RECT  10.560 1.200 10.800 2.200 ;
        RECT  10.560 1.960 12.290 2.200 ;
        RECT  11.890 1.960 12.290 2.220 ;
        RECT  5.130 2.020 5.410 2.860 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  33.200 1.840 34.640 2.080 ;
        RECT  34.400 1.200 34.640 2.080 ;
        RECT  34.400 1.200 37.900 1.440 ;
        RECT  37.660 1.200 37.900 2.320 ;
        RECT  37.660 2.080 40.100 2.320 ;
        RECT  32.860 1.980 33.440 2.220 ;
        END
    END CI0
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.050 2.800 2.360 3.200 ;
        RECT  2.010 1.320 2.410 1.560 ;
        RECT  4.530 1.460 4.770 3.760 ;
        RECT  2.050 3.520 4.770 3.760 ;
        RECT  4.530 1.460 4.880 1.860 ;
        RECT  4.530 3.100 5.120 3.340 ;
        RECT  2.050 1.320 2.290 3.760 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  40.080 3.100 40.730 3.340 ;
        RECT  40.490 1.460 40.730 3.760 ;
        RECT  42.890 2.800 43.210 3.200 ;
        RECT  42.970 1.380 43.210 3.760 ;
        RECT  40.490 3.520 43.210 3.760 ;
        RECT  42.830 1.380 43.230 1.620 ;
        RECT  40.320 1.460 40.730 1.860 ;
        END
    END CO0
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  20.650 1.500 20.890 3.280 ;
        RECT  20.570 3.040 20.970 3.280 ;
        RECT  20.270 2.380 20.890 2.660 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 1.800 0.480 2.200 ;
        RECT  0.190 4.000 13.890 4.240 ;
        RECT  13.650 4.180 16.670 4.420 ;
        RECT  16.430 4.000 17.790 4.240 ;
        RECT  18.780 4.080 19.180 4.420 ;
        RECT  17.550 4.180 20.260 4.420 ;
        RECT  20.020 4.000 23.030 4.240 ;
        RECT  24.610 4.080 25.010 4.420 ;
        RECT  22.790 4.180 27.560 4.420 ;
        RECT  27.320 4.000 28.790 4.240 ;
        RECT  28.550 4.180 31.460 4.420 ;
        RECT  31.220 4.000 45.070 4.240 ;
        RECT  44.830 2.520 45.070 4.240 ;
        RECT  44.700 2.520 45.100 2.760 ;
        RECT  0.190 1.800 0.430 4.240 ;
        END
    END B
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  21.870 2.060 22.150 2.800 ;
        RECT  21.810 2.040 22.050 2.440 ;
        END
    END CS
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.740 2.520 1.140 2.760 ;
        RECT  0.770 0.800 4.290 1.040 ;
        RECT  4.050 0.620 4.290 2.310 ;
        RECT  3.210 2.070 4.290 2.310 ;
        RECT  4.050 0.620 5.390 0.860 ;
        RECT  5.150 0.800 6.980 1.040 ;
        RECT  6.740 0.720 11.280 0.960 ;
        RECT  12.000 0.620 12.240 1.200 ;
        RECT  11.040 0.960 12.240 1.200 ;
        RECT  12.000 0.620 15.890 0.860 ;
        RECT  15.650 0.620 15.890 1.250 ;
        RECT  16.610 0.620 16.850 1.250 ;
        RECT  15.650 1.010 16.850 1.250 ;
        RECT  16.610 0.620 19.660 0.860 ;
        RECT  19.420 0.620 19.660 1.130 ;
        RECT  20.540 0.620 20.780 1.130 ;
        RECT  19.420 0.890 20.780 1.130 ;
        RECT  20.540 0.620 24.230 0.860 ;
        RECT  23.990 0.620 24.230 1.130 ;
        RECT  24.950 0.620 25.190 1.130 ;
        RECT  23.990 0.890 25.190 1.130 ;
        RECT  24.950 0.620 29.620 0.860 ;
        RECT  29.380 0.720 33.110 0.960 ;
        RECT  32.870 0.960 34.070 1.200 ;
        RECT  33.830 0.720 38.380 0.960 ;
        RECT  38.140 0.800 39.970 1.040 ;
        RECT  39.730 0.720 41.210 0.960 ;
        RECT  40.970 0.720 41.210 2.310 ;
        RECT  40.970 2.070 42.050 2.310 ;
        RECT  40.960 0.800 44.470 1.040 ;
        RECT  44.190 0.800 44.470 2.120 ;
        RECT  44.120 1.880 44.520 2.120 ;
        RECT  0.770 0.800 1.010 2.760 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.060 -0.380 6.460 0.560 ;
        RECT  11.520 -0.380 11.760 0.640 ;
        RECT  16.130 -0.380 16.370 0.640 ;
        RECT  19.950 -0.380 20.190 0.650 ;
        RECT  24.470 -0.380 24.710 0.650 ;
        RECT  33.350 -0.380 33.590 0.640 ;
        RECT  38.740 -0.380 39.140 0.560 ;
        RECT  42.040 -0.380 42.440 0.560 ;
        RECT  43.640 -0.380 44.040 0.560 ;
        RECT  0.000 -0.380 45.260 0.380 ;
        RECT  1.680 -0.380 3.160 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.850 4.480 3.250 5.420 ;
        RECT  6.280 4.480 6.680 5.420 ;
        RECT  8.410 4.480 8.810 5.420 ;
        RECT  10.710 4.480 11.110 5.420 ;
        RECT  13.010 4.480 13.410 5.420 ;
        RECT  16.910 4.480 17.310 5.420 ;
        RECT  20.500 4.480 22.520 5.420 ;
        RECT  27.910 4.480 28.310 5.420 ;
        RECT  31.730 4.480 32.130 5.420 ;
        RECT  34.000 4.480 34.400 5.420 ;
        RECT  36.390 4.480 36.790 5.420 ;
        RECT  38.520 4.480 38.920 5.420 ;
        RECT  42.010 4.480 42.410 5.420 ;
        RECT  43.540 4.480 44.820 5.420 ;
        RECT  0.000 4.660 45.260 5.420 ;
        RECT  0.440 4.480 1.720 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  43.630 3.060 44.590 3.300 ;
        RECT  43.630 1.340 43.870 3.300 ;
        RECT  43.520 1.860 43.870 2.260 ;
        RECT  43.550 1.340 43.950 1.580 ;
        RECT  40.970 3.030 42.590 3.270 ;
        RECT  42.350 1.590 42.590 3.270 ;
        RECT  42.350 1.840 42.660 2.240 ;
        RECT  41.450 1.590 42.590 1.830 ;
        RECT  41.450 1.300 41.690 1.830 ;
        RECT  38.140 1.440 38.380 1.840 ;
        RECT  38.140 1.540 39.870 1.780 ;
        RECT  37.900 3.100 39.650 3.340 ;
        RECT  37.020 2.980 37.420 3.220 ;
        RECT  37.180 1.680 37.420 3.220 ;
        RECT  37.180 2.560 39.310 2.800 ;
        RECT  37.020 1.680 37.420 1.920 ;
        RECT  35.760 3.520 37.610 3.760 ;
        RECT  35.760 1.680 36.000 3.760 ;
        RECT  35.600 2.980 36.000 3.220 ;
        RECT  35.600 1.680 36.000 1.920 ;
        RECT  31.090 3.520 35.200 3.760 ;
        RECT  34.960 1.680 35.200 3.760 ;
        RECT  31.090 1.680 31.330 3.760 ;
        RECT  34.880 2.980 35.280 3.220 ;
        RECT  33.540 2.440 35.200 2.680 ;
        RECT  34.880 1.680 35.280 1.920 ;
        RECT  31.010 1.680 31.410 1.920 ;
        RECT  29.570 3.220 30.050 3.460 ;
        RECT  29.810 1.200 30.050 3.460 ;
        RECT  32.380 2.980 32.970 3.220 ;
        RECT  32.380 1.200 32.620 3.220 ;
        RECT  29.570 1.680 30.050 1.920 ;
        RECT  32.380 1.440 32.970 1.680 ;
        RECT  29.810 1.200 32.620 1.440 ;
        RECT  31.730 3.040 32.130 3.280 ;
        RECT  31.780 1.680 32.020 3.280 ;
        RECT  31.670 2.240 32.020 2.640 ;
        RECT  31.730 1.680 32.130 1.920 ;
        RECT  29.030 3.700 30.610 3.940 ;
        RECT  30.370 1.680 30.610 3.940 ;
        RECT  27.940 3.520 29.270 3.760 ;
        RECT  27.940 2.710 28.180 3.760 ;
        RECT  30.290 3.220 30.690 3.460 ;
        RECT  27.880 2.710 28.180 3.110 ;
        RECT  30.290 1.680 30.690 1.920 ;
        RECT  25.870 3.120 26.270 3.360 ;
        RECT  28.850 3.040 29.250 3.280 ;
        RECT  25.950 1.100 26.190 3.360 ;
        RECT  28.900 1.490 29.140 3.280 ;
        RECT  27.950 1.490 29.140 1.730 ;
        RECT  27.950 1.100 28.190 1.730 ;
        RECT  25.950 1.100 28.190 1.340 ;
        RECT  27.380 3.360 27.700 3.760 ;
        RECT  27.380 1.580 27.620 3.760 ;
        RECT  28.420 2.040 28.660 2.440 ;
        RECT  27.380 2.120 28.660 2.360 ;
        RECT  27.310 1.580 27.710 1.820 ;
        RECT  24.390 3.600 26.910 3.840 ;
        RECT  26.670 1.580 26.910 3.840 ;
        RECT  24.390 1.500 24.630 3.840 ;
        RECT  26.590 1.580 26.990 1.820 ;
        RECT  25.130 2.880 25.550 3.120 ;
        RECT  25.130 1.580 25.370 3.120 ;
        RECT  25.130 2.140 25.610 2.540 ;
        RECT  25.130 1.580 25.550 1.820 ;
        RECT  23.510 3.040 23.910 3.440 ;
        RECT  23.510 1.100 23.750 3.440 ;
        RECT  21.130 2.420 21.510 2.820 ;
        RECT  21.270 1.100 21.510 2.820 ;
        RECT  23.510 1.500 23.910 1.900 ;
        RECT  21.270 1.100 23.750 1.340 ;
        RECT  18.450 3.600 19.840 3.840 ;
        RECT  22.970 1.580 23.210 3.760 ;
        RECT  19.600 3.520 23.210 3.760 ;
        RECT  22.950 3.040 23.210 3.760 ;
        RECT  18.450 1.580 18.690 3.840 ;
        RECT  18.370 3.040 18.690 3.440 ;
        RECT  22.870 1.580 23.270 1.820 ;
        RECT  18.290 1.580 18.690 1.820 ;
        RECT  22.150 3.040 22.630 3.280 ;
        RECT  22.390 1.580 22.630 3.280 ;
        RECT  22.390 2.320 22.730 2.720 ;
        RECT  22.150 1.580 22.630 1.820 ;
        RECT  19.730 2.970 20.130 3.210 ;
        RECT  19.790 1.580 20.030 3.210 ;
        RECT  19.600 2.330 20.030 2.730 ;
        RECT  19.730 1.580 20.130 1.820 ;
        RECT  19.010 3.120 19.410 3.360 ;
        RECT  15.830 3.040 16.380 3.280 ;
        RECT  19.090 1.500 19.330 3.360 ;
        RECT  15.830 1.490 16.070 3.280 ;
        RECT  18.930 1.100 19.170 1.920 ;
        RECT  15.830 1.490 16.220 1.900 ;
        RECT  15.830 1.490 17.330 1.730 ;
        RECT  17.090 1.100 17.330 1.730 ;
        RECT  17.090 1.100 19.170 1.340 ;
        RECT  17.500 3.520 17.900 3.760 ;
        RECT  17.660 1.580 17.900 3.760 ;
        RECT  16.600 2.040 16.840 2.440 ;
        RECT  16.600 2.040 17.900 2.280 ;
        RECT  17.570 1.580 17.900 2.280 ;
        RECT  17.570 1.580 17.970 1.820 ;
        RECT  14.530 3.700 16.190 3.940 ;
        RECT  17.020 2.710 17.260 3.760 ;
        RECT  15.950 3.520 17.260 3.760 ;
        RECT  14.530 1.680 14.770 3.940 ;
        RECT  14.450 3.220 14.850 3.460 ;
        RECT  17.020 2.710 17.350 3.110 ;
        RECT  14.450 1.680 14.850 1.920 ;
        RECT  15.170 3.220 15.570 3.460 ;
        RECT  12.170 2.980 12.770 3.220 ;
        RECT  12.530 1.200 12.770 3.220 ;
        RECT  15.170 1.200 15.410 3.460 ;
        RECT  15.170 1.680 15.570 1.920 ;
        RECT  12.170 1.440 12.770 1.680 ;
        RECT  12.530 1.200 15.410 1.440 ;
        RECT  9.940 3.520 14.050 3.760 ;
        RECT  13.810 1.680 14.050 3.760 ;
        RECT  9.940 2.980 10.180 3.760 ;
        RECT  9.920 2.980 10.320 3.220 ;
        RECT  9.930 1.680 10.170 3.220 ;
        RECT  9.930 2.440 11.580 2.680 ;
        RECT  13.730 1.680 14.130 1.920 ;
        RECT  9.920 1.680 10.320 1.920 ;
        RECT  13.010 3.040 13.410 3.280 ;
        RECT  13.090 1.680 13.330 3.280 ;
        RECT  13.090 2.240 13.470 2.640 ;
        RECT  13.010 1.680 13.410 1.920 ;
        RECT  7.590 3.520 9.440 3.760 ;
        RECT  9.200 1.680 9.440 3.760 ;
        RECT  9.200 2.980 9.600 3.220 ;
        RECT  9.200 1.680 9.600 1.920 ;
        RECT  7.780 2.980 8.180 3.220 ;
        RECT  7.780 1.680 8.020 3.220 ;
        RECT  5.890 2.560 8.020 2.800 ;
        RECT  7.780 1.680 8.180 1.920 ;
        RECT  5.550 3.100 7.300 3.340 ;
        RECT  6.820 1.440 7.060 1.840 ;
        RECT  5.330 1.540 7.060 1.780 ;
        RECT  2.670 3.030 4.280 3.270 ;
        RECT  2.670 1.320 2.910 3.270 ;
        RECT  2.570 1.840 2.910 2.240 ;
        RECT  2.670 1.320 3.810 1.560 ;
        RECT  0.670 3.060 1.770 3.300 ;
        RECT  1.530 1.340 1.770 3.300 ;
        RECT  1.250 1.340 1.770 1.580 ;
    END
END FACS1S

MACRO FACS2
    CLASS CORE ;
    FOREIGN FACS2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 54.560 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.210 2.080 7.250 2.320 ;
        RECT  7.010 2.050 8.490 2.290 ;
        RECT  9.660 1.200 9.900 2.320 ;
        RECT  8.250 2.080 9.900 2.320 ;
        RECT  9.660 1.200 15.310 1.440 ;
        RECT  15.070 1.200 15.310 2.080 ;
        RECT  16.150 1.920 16.790 2.160 ;
        RECT  15.070 1.840 16.390 2.080 ;
        RECT  16.390 1.920 16.790 2.220 ;
        RECT  6.210 2.080 6.610 2.380 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  38.010 1.840 39.350 2.080 ;
        RECT  39.110 1.200 39.350 2.080 ;
        RECT  39.110 1.200 44.730 1.440 ;
        RECT  44.490 1.200 44.730 2.300 ;
        RECT  44.490 2.060 45.710 2.300 ;
        RECT  45.470 2.050 47.430 2.290 ;
        RECT  47.190 2.120 48.200 2.360 ;
        RECT  37.560 1.980 38.250 2.220 ;
        END
    END CI0
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.010 1.300 2.290 1.700 ;
        RECT  2.010 2.800 2.360 3.200 ;
        RECT  4.360 1.100 4.600 2.550 ;
        RECT  4.530 2.310 4.770 3.940 ;
        RECT  2.010 3.520 4.770 3.760 ;
        RECT  4.360 1.100 5.960 1.340 ;
        RECT  5.850 3.100 6.090 3.940 ;
        RECT  4.530 3.700 6.090 3.940 ;
        RECT  5.770 3.100 6.170 3.340 ;
        RECT  2.010 1.300 2.250 3.760 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  48.240 3.100 48.640 3.340 ;
        RECT  48.470 1.100 50.030 1.340 ;
        RECT  49.790 1.100 50.030 3.940 ;
        RECT  48.320 3.700 50.030 3.940 ;
        RECT  52.210 1.300 52.580 1.700 ;
        RECT  52.190 2.800 52.580 3.200 ;
        RECT  49.790 3.520 52.580 3.760 ;
        RECT  52.340 1.300 52.580 3.760 ;
        RECT  48.320 3.100 48.560 3.940 ;
        END
    END CO0
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  24.990 1.500 25.410 1.900 ;
        RECT  24.990 3.040 25.470 3.280 ;
        RECT  24.990 1.500 25.230 3.280 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.470 4.000 18.410 4.240 ;
        RECT  18.170 4.180 21.170 4.420 ;
        RECT  20.930 4.000 22.750 4.240 ;
        RECT  22.510 4.080 24.760 4.320 ;
        RECT  24.520 4.000 27.710 4.240 ;
        RECT  27.470 4.080 32.260 4.320 ;
        RECT  32.020 4.000 33.490 4.240 ;
        RECT  33.250 4.180 36.160 4.420 ;
        RECT  35.920 4.000 40.760 4.240 ;
        RECT  40.480 3.460 40.760 4.240 ;
        RECT  13.810 3.460 14.090 4.240 ;
        END
    END B
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  26.210 2.060 26.670 2.460 ;
        RECT  26.210 2.060 26.490 2.800 ;
        END
    END CS
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.510 0.620 16.750 1.200 ;
        RECT  15.550 0.960 16.750 1.200 ;
        RECT  16.510 0.620 20.390 0.860 ;
        RECT  20.150 0.620 20.390 1.250 ;
        RECT  21.110 0.620 21.350 1.250 ;
        RECT  20.150 1.010 21.350 1.250 ;
        RECT  21.110 0.620 24.160 0.860 ;
        RECT  23.920 0.620 24.160 1.130 ;
        RECT  25.040 0.620 25.280 1.130 ;
        RECT  23.920 0.890 25.280 1.130 ;
        RECT  25.040 0.620 28.970 0.860 ;
        RECT  28.730 0.620 28.970 1.130 ;
        RECT  29.950 0.620 30.190 1.130 ;
        RECT  28.730 0.890 30.190 1.130 ;
        RECT  33.180 0.620 33.790 0.980 ;
        RECT  29.950 0.620 33.910 0.860 ;
        RECT  33.180 0.720 37.810 0.960 ;
        RECT  37.570 0.960 38.870 1.200 ;
        RECT  38.630 0.620 38.870 1.590 ;
        RECT  38.630 0.720 43.070 0.960 ;
        RECT  11.330 0.720 15.790 0.960 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.760 -0.380 3.160 0.560 ;
        RECT  7.020 -0.380 7.420 0.560 ;
        RECT  8.480 -0.380 8.880 0.560 ;
        RECT  16.030 -0.380 16.270 0.640 ;
        RECT  20.630 -0.380 20.870 0.640 ;
        RECT  24.450 -0.380 24.690 0.650 ;
        RECT  29.210 -0.380 29.450 0.650 ;
        RECT  38.050 -0.380 38.290 0.640 ;
        RECT  45.530 -0.380 45.930 0.560 ;
        RECT  46.990 -0.380 47.390 0.560 ;
        RECT  51.340 -0.380 51.740 0.560 ;
        RECT  52.940 -0.380 53.340 0.560 ;
        RECT  0.000 -0.380 54.560 0.380 ;
        RECT  1.230 -0.380 1.630 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.850 4.480 3.250 5.420 ;
        RECT  7.330 4.180 7.730 5.420 ;
        RECT  8.790 4.180 9.190 5.420 ;
        RECT  10.990 4.480 11.390 5.420 ;
        RECT  12.850 4.480 13.250 5.420 ;
        RECT  15.210 4.480 15.610 5.420 ;
        RECT  17.510 4.480 17.910 5.420 ;
        RECT  21.410 4.480 21.810 5.420 ;
        RECT  26.080 4.480 27.020 5.420 ;
        RECT  32.610 4.480 33.010 5.420 ;
        RECT  36.430 4.480 36.830 5.420 ;
        RECT  38.700 4.480 39.100 5.420 ;
        RECT  40.870 4.480 41.270 5.420 ;
        RECT  43.010 4.480 43.410 5.420 ;
        RECT  45.220 4.180 45.620 5.420 ;
        RECT  46.680 4.180 47.080 5.420 ;
        RECT  51.310 4.480 51.710 5.420 ;
        RECT  52.840 4.480 54.120 5.420 ;
        RECT  0.000 4.660 54.560 5.420 ;
        RECT  0.440 4.480 1.720 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  47.500 4.180 50.740 4.420 ;
        RECT  43.650 4.180 44.980 4.420 ;
        RECT  44.740 3.580 44.980 4.420 ;
        RECT  54.130 2.520 54.370 4.240 ;
        RECT  41.490 4.000 43.890 4.240 ;
        RECT  50.500 4.000 54.370 4.240 ;
        RECT  47.500 3.580 47.740 4.420 ;
        RECT  44.740 3.580 47.740 3.820 ;
        RECT  54.000 2.520 54.400 2.760 ;
        RECT  52.930 3.060 53.890 3.300 ;
        RECT  52.930 1.340 53.170 3.300 ;
        RECT  52.820 1.860 53.170 2.260 ;
        RECT  52.850 1.340 53.250 1.580 ;
        RECT  50.380 2.060 51.410 2.300 ;
        RECT  53.420 1.880 53.820 2.120 ;
        RECT  50.380 0.620 50.620 2.300 ;
        RECT  53.490 0.800 53.770 2.120 ;
        RECT  50.380 0.800 53.770 1.040 ;
        RECT  44.970 0.800 47.870 1.040 ;
        RECT  43.620 0.720 45.210 0.960 ;
        RECT  47.630 0.620 50.620 0.860 ;
        RECT  50.270 3.030 51.950 3.270 ;
        RECT  51.710 1.580 51.950 3.270 ;
        RECT  51.710 1.840 52.010 2.240 ;
        RECT  50.860 1.580 51.950 1.820 ;
        RECT  50.860 1.300 51.100 1.820 ;
        RECT  49.280 1.580 49.520 1.980 ;
        RECT  47.610 1.580 49.520 1.820 ;
        RECT  44.970 1.420 45.210 1.820 ;
        RECT  44.970 1.570 47.850 1.810 ;
        RECT  48.960 3.100 49.410 3.340 ;
        RECT  49.170 2.620 49.410 3.340 ;
        RECT  44.600 3.100 47.920 3.340 ;
        RECT  47.680 2.620 47.920 3.340 ;
        RECT  47.680 2.620 49.410 2.860 ;
        RECT  43.850 2.980 44.250 3.220 ;
        RECT  44.010 1.680 44.250 3.220 ;
        RECT  44.010 2.540 46.950 2.780 ;
        RECT  46.550 2.530 46.950 2.780 ;
        RECT  43.850 1.680 44.250 1.920 ;
        RECT  44.130 3.520 44.370 3.920 ;
        RECT  41.800 3.520 44.370 3.760 ;
        RECT  41.800 1.680 42.040 3.760 ;
        RECT  41.720 2.980 42.120 3.220 ;
        RECT  41.720 1.680 42.120 1.920 ;
        RECT  42.440 2.980 42.840 3.220 ;
        RECT  42.520 1.680 42.760 3.220 ;
        RECT  42.520 2.320 43.750 2.560 ;
        RECT  42.440 1.680 42.840 1.920 ;
        RECT  40.310 2.980 40.710 3.220 ;
        RECT  40.390 1.680 40.630 3.220 ;
        RECT  41.300 2.240 41.540 2.640 ;
        RECT  40.390 2.320 41.540 2.560 ;
        RECT  40.310 1.680 40.710 1.920 ;
        RECT  35.790 3.520 39.910 3.760 ;
        RECT  39.670 1.680 39.910 3.760 ;
        RECT  35.790 1.680 36.030 3.760 ;
        RECT  39.590 2.980 39.990 3.220 ;
        RECT  38.510 2.440 39.910 2.680 ;
        RECT  39.590 1.680 39.990 1.920 ;
        RECT  35.710 1.680 36.110 1.920 ;
        RECT  34.270 3.220 34.750 3.460 ;
        RECT  34.510 1.200 34.750 3.460 ;
        RECT  37.080 2.980 37.670 3.220 ;
        RECT  37.080 1.200 37.320 3.220 ;
        RECT  34.270 1.680 34.750 1.920 ;
        RECT  37.080 1.440 37.670 1.680 ;
        RECT  34.510 1.200 37.320 1.440 ;
        RECT  36.430 3.040 36.830 3.280 ;
        RECT  36.480 1.680 36.720 3.280 ;
        RECT  36.370 2.240 36.720 2.640 ;
        RECT  36.430 1.680 36.830 1.920 ;
        RECT  33.730 3.700 35.310 3.940 ;
        RECT  35.070 1.680 35.310 3.940 ;
        RECT  32.640 3.520 33.970 3.760 ;
        RECT  32.640 2.710 32.880 3.760 ;
        RECT  34.990 3.220 35.390 3.460 ;
        RECT  32.580 2.710 32.880 3.110 ;
        RECT  34.990 1.680 35.390 1.920 ;
        RECT  30.570 3.120 30.970 3.360 ;
        RECT  33.550 3.040 33.950 3.280 ;
        RECT  30.650 1.100 30.890 3.360 ;
        RECT  33.600 1.490 33.840 3.280 ;
        RECT  32.650 1.490 33.840 1.730 ;
        RECT  32.650 1.100 32.890 1.730 ;
        RECT  30.650 1.100 32.890 1.340 ;
        RECT  32.080 3.360 32.400 3.760 ;
        RECT  32.080 1.580 32.320 3.760 ;
        RECT  33.120 2.040 33.360 2.440 ;
        RECT  32.080 2.120 33.360 2.360 ;
        RECT  32.010 1.580 32.410 1.820 ;
        RECT  29.090 3.600 31.610 3.840 ;
        RECT  31.370 1.580 31.610 3.840 ;
        RECT  29.090 1.500 29.330 3.840 ;
        RECT  31.290 1.580 31.690 1.820 ;
        RECT  29.830 2.880 30.250 3.120 ;
        RECT  29.830 1.580 30.070 3.120 ;
        RECT  29.830 2.140 30.310 2.540 ;
        RECT  29.830 1.580 30.250 1.820 ;
        RECT  28.250 3.040 28.610 3.440 ;
        RECT  28.250 1.100 28.490 3.440 ;
        RECT  25.650 2.310 25.970 2.710 ;
        RECT  25.650 1.100 25.890 2.710 ;
        RECT  28.250 1.500 28.610 1.900 ;
        RECT  25.650 1.100 28.490 1.340 ;
        RECT  22.950 3.600 24.340 3.840 ;
        RECT  27.770 1.580 28.010 3.760 ;
        RECT  24.100 3.520 28.010 3.760 ;
        RECT  27.650 3.040 28.010 3.760 ;
        RECT  22.950 1.580 23.190 3.840 ;
        RECT  22.870 3.040 23.190 3.440 ;
        RECT  27.570 1.580 28.010 1.820 ;
        RECT  22.790 1.580 23.190 1.820 ;
        RECT  26.650 3.040 27.250 3.280 ;
        RECT  27.010 1.580 27.250 3.280 ;
        RECT  27.010 2.320 27.350 2.720 ;
        RECT  26.650 1.580 27.250 1.820 ;
        RECT  24.230 2.970 24.630 3.210 ;
        RECT  24.290 1.580 24.530 3.210 ;
        RECT  24.100 2.330 24.530 2.730 ;
        RECT  24.230 1.580 24.630 1.820 ;
        RECT  23.510 3.120 23.910 3.360 ;
        RECT  20.330 3.040 20.880 3.280 ;
        RECT  23.590 1.500 23.830 3.360 ;
        RECT  20.330 1.490 20.570 3.280 ;
        RECT  23.430 1.100 23.670 1.920 ;
        RECT  20.330 1.490 20.720 1.900 ;
        RECT  20.330 1.490 21.830 1.730 ;
        RECT  21.590 1.100 21.830 1.730 ;
        RECT  21.590 1.100 23.670 1.340 ;
        RECT  22.000 3.520 22.400 3.760 ;
        RECT  22.160 1.580 22.400 3.760 ;
        RECT  21.100 2.040 21.340 2.440 ;
        RECT  21.100 2.040 22.400 2.280 ;
        RECT  22.070 1.580 22.400 2.280 ;
        RECT  22.070 1.580 22.470 1.820 ;
        RECT  19.030 3.700 20.690 3.940 ;
        RECT  21.520 2.710 21.760 3.760 ;
        RECT  20.450 3.520 21.760 3.760 ;
        RECT  19.030 1.680 19.270 3.940 ;
        RECT  18.950 3.220 19.350 3.460 ;
        RECT  21.520 2.710 21.850 3.110 ;
        RECT  18.950 1.680 19.350 1.920 ;
        RECT  19.670 3.220 20.070 3.460 ;
        RECT  16.670 2.980 17.270 3.220 ;
        RECT  17.030 1.200 17.270 3.220 ;
        RECT  19.670 1.200 19.910 3.460 ;
        RECT  19.670 1.680 20.070 1.920 ;
        RECT  16.670 1.440 17.270 1.680 ;
        RECT  17.030 1.200 19.910 1.440 ;
        RECT  14.440 3.520 18.550 3.760 ;
        RECT  18.310 1.680 18.550 3.760 ;
        RECT  14.440 2.980 14.680 3.760 ;
        RECT  14.420 2.980 14.820 3.220 ;
        RECT  14.430 1.680 14.670 3.220 ;
        RECT  14.430 2.440 16.080 2.680 ;
        RECT  18.230 1.680 18.630 1.920 ;
        RECT  14.420 1.680 14.820 1.920 ;
        RECT  17.510 3.040 17.910 3.280 ;
        RECT  17.590 1.680 17.830 3.280 ;
        RECT  17.590 2.240 17.970 2.640 ;
        RECT  17.510 1.680 17.910 1.920 ;
        RECT  13.700 2.980 14.100 3.220 ;
        RECT  13.780 1.680 14.020 3.220 ;
        RECT  12.870 2.240 13.110 2.640 ;
        RECT  12.870 2.320 14.020 2.560 ;
        RECT  13.700 1.680 14.100 1.920 ;
        RECT  9.430 4.180 10.750 4.420 ;
        RECT  3.830 4.180 7.090 4.420 ;
        RECT  6.850 3.580 7.090 4.420 ;
        RECT  10.510 4.000 12.690 4.240 ;
        RECT  0.190 4.000 4.070 4.240 ;
        RECT  9.430 3.580 9.670 4.420 ;
        RECT  0.190 1.800 0.430 4.240 ;
        RECT  6.850 3.580 9.670 3.820 ;
        RECT  0.190 1.800 0.480 2.200 ;
        RECT  10.030 3.460 10.270 3.860 ;
        RECT  10.030 3.520 12.600 3.760 ;
        RECT  12.360 1.680 12.600 3.760 ;
        RECT  12.280 2.980 12.680 3.220 ;
        RECT  12.280 1.680 12.680 1.920 ;
        RECT  11.560 2.980 11.960 3.220 ;
        RECT  11.640 1.680 11.880 3.220 ;
        RECT  10.650 2.320 11.880 2.560 ;
        RECT  11.560 1.680 11.960 1.920 ;
        RECT  0.740 2.520 1.140 2.760 ;
        RECT  0.770 0.800 1.010 2.760 ;
        RECT  3.090 2.070 4.120 2.310 ;
        RECT  3.880 0.620 4.120 2.310 ;
        RECT  6.540 0.800 9.340 1.040 ;
        RECT  0.770 0.800 4.120 1.040 ;
        RECT  9.100 0.720 10.770 0.960 ;
        RECT  3.880 0.620 6.780 0.860 ;
        RECT  10.140 2.980 10.540 3.220 ;
        RECT  10.140 1.680 10.380 3.220 ;
        RECT  7.460 2.560 10.380 2.800 ;
        RECT  7.460 2.530 7.860 2.800 ;
        RECT  10.140 1.680 10.540 1.920 ;
        RECT  6.490 3.100 9.810 3.340 ;
        RECT  5.050 3.100 5.450 3.340 ;
        RECT  6.490 2.620 6.730 3.340 ;
        RECT  5.050 2.620 5.290 3.340 ;
        RECT  5.050 2.620 6.730 2.860 ;
        RECT  9.180 1.440 9.420 1.840 ;
        RECT  4.840 1.600 6.680 1.840 ;
        RECT  6.440 1.570 9.420 1.810 ;
        RECT  2.600 3.030 4.280 3.270 ;
        RECT  2.600 1.380 2.840 3.270 ;
        RECT  2.490 1.840 2.840 2.240 ;
        RECT  3.400 1.300 3.640 1.700 ;
        RECT  2.600 1.380 3.640 1.620 ;
        RECT  0.670 3.060 1.770 3.300 ;
        RECT  1.530 1.340 1.770 3.300 ;
        RECT  1.250 1.340 1.770 1.580 ;
    END
END FACS2

MACRO FACS2P
    CLASS CORE ;
    FOREIGN FACS2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 66.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.090 2.050 14.680 2.290 ;
        RECT  15.380 1.200 15.620 2.320 ;
        RECT  14.440 2.080 15.620 2.320 ;
        RECT  15.380 1.200 21.020 1.440 ;
        RECT  20.780 1.200 21.020 2.080 ;
        RECT  21.890 1.920 22.510 2.160 ;
        RECT  20.780 1.840 22.130 2.080 ;
        RECT  22.110 1.920 22.510 2.220 ;
        RECT  8.650 2.140 11.330 2.380 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  44.120 1.980 44.520 2.220 ;
        RECT  44.120 1.980 45.070 2.160 ;
        RECT  44.830 1.840 45.900 2.080 ;
        RECT  44.130 1.920 45.900 2.080 ;
        RECT  45.660 1.200 45.900 2.080 ;
        RECT  45.660 1.200 51.300 1.440 ;
        RECT  51.060 1.200 51.300 2.380 ;
        RECT  51.060 2.140 52.330 2.380 ;
        RECT  52.090 2.050 55.720 2.290 ;
        RECT  55.480 2.120 58.160 2.360 ;
        RECT  57.760 2.120 58.160 2.380 ;
        RECT  44.190 1.920 44.470 2.740 ;
        END
    END CI0
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.170 2.800 2.410 3.200 ;
        RECT  2.670 1.440 2.910 3.760 ;
        RECT  2.170 2.880 3.650 3.120 ;
        RECT  2.050 1.440 3.670 1.680 ;
        RECT  3.410 2.800 3.650 3.200 ;
        RECT  3.430 1.360 3.670 1.760 ;
        RECT  5.700 1.100 5.940 2.550 ;
        RECT  5.860 2.310 6.100 3.940 ;
        RECT  2.670 3.520 6.100 3.760 ;
        RECT  7.060 3.100 7.300 3.940 ;
        RECT  6.980 3.100 7.380 3.340 ;
        RECT  8.500 3.100 8.740 3.940 ;
        RECT  5.860 3.700 8.740 3.940 ;
        RECT  5.700 1.100 8.770 1.340 ;
        RECT  8.420 3.100 8.820 3.340 ;
        RECT  2.050 1.360 2.290 1.760 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  57.990 3.100 58.390 3.340 ;
        RECT  59.510 3.100 59.750 3.940 ;
        RECT  59.430 3.100 59.830 3.340 ;
        RECT  57.920 1.100 60.980 1.340 ;
        RECT  60.710 2.520 60.950 3.940 ;
        RECT  58.070 3.700 60.950 3.940 ;
        RECT  60.740 1.100 60.980 2.760 ;
        RECT  63.230 1.360 63.470 1.760 ;
        RECT  63.250 2.800 63.490 3.200 ;
        RECT  60.710 3.520 64.290 3.760 ;
        RECT  64.050 1.440 64.290 3.760 ;
        RECT  63.230 1.440 64.850 1.680 ;
        RECT  63.250 2.880 64.810 3.120 ;
        RECT  64.610 1.360 64.850 1.760 ;
        RECT  58.070 3.100 58.310 3.940 ;
        END
    END CO0
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  31.170 1.500 31.970 1.900 ;
        RECT  31.170 3.040 32.030 3.280 ;
        RECT  31.170 1.500 31.450 3.280 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  19.190 4.000 24.110 4.240 ;
        RECT  23.870 4.180 26.890 4.420 ;
        RECT  26.650 4.000 28.010 4.240 ;
        RECT  29.000 4.080 29.400 4.420 ;
        RECT  27.770 4.180 30.480 4.420 ;
        RECT  30.240 4.000 34.290 4.240 ;
        RECT  35.870 4.080 36.270 4.420 ;
        RECT  34.050 4.180 38.820 4.420 ;
        RECT  38.580 4.000 40.050 4.240 ;
        RECT  39.810 4.180 42.720 4.420 ;
        RECT  42.480 4.000 47.270 4.240 ;
        RECT  19.390 3.460 19.670 4.240 ;
        END
    END B
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  33.030 2.060 33.310 2.800 ;
        RECT  32.970 2.060 33.310 2.460 ;
        END
    END CS
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  21.870 0.900 22.150 1.600 ;
        RECT  22.220 0.620 22.460 1.140 ;
        RECT  21.260 0.900 22.460 1.140 ;
        RECT  22.220 0.620 26.110 0.860 ;
        RECT  25.870 0.620 26.110 1.250 ;
        RECT  26.830 0.620 27.070 1.250 ;
        RECT  25.870 1.010 27.070 1.250 ;
        RECT  26.830 0.620 29.880 0.860 ;
        RECT  29.640 0.620 29.880 1.130 ;
        RECT  31.600 0.620 31.840 1.130 ;
        RECT  29.640 0.890 31.840 1.130 ;
        RECT  31.600 0.620 35.530 0.860 ;
        RECT  35.290 0.620 35.530 1.130 ;
        RECT  36.580 0.620 36.820 1.130 ;
        RECT  35.290 0.890 36.820 1.130 ;
        RECT  36.580 0.620 40.730 0.860 ;
        RECT  40.490 0.720 44.460 0.960 ;
        RECT  44.220 0.960 45.420 1.200 ;
        RECT  45.180 0.720 49.650 0.960 ;
        RECT  17.050 0.720 21.500 0.960 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.070 -0.380 4.470 0.560 ;
        RECT  9.820 -0.380 10.220 0.560 ;
        RECT  11.280 -0.380 11.680 0.560 ;
        RECT  12.740 -0.380 13.140 0.560 ;
        RECT  14.200 -0.380 14.600 0.560 ;
        RECT  21.740 -0.380 21.980 0.640 ;
        RECT  26.350 -0.380 26.590 0.640 ;
        RECT  30.120 -0.380 31.110 0.650 ;
        RECT  35.770 -0.380 36.010 0.650 ;
        RECT  44.700 -0.380 44.940 0.640 ;
        RECT  52.080 -0.380 52.480 0.560 ;
        RECT  53.540 -0.380 53.940 0.560 ;
        RECT  55.000 -0.380 55.400 0.560 ;
        RECT  56.460 -0.380 56.860 0.560 ;
        RECT  62.430 -0.380 62.830 0.560 ;
        RECT  65.340 -0.380 65.740 0.560 ;
        RECT  0.000 -0.380 66.960 0.380 ;
        RECT  1.230 -0.380 1.630 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.750 4.480 3.150 5.420 ;
        RECT  4.090 4.480 4.490 5.420 ;
        RECT  9.980 4.180 10.380 5.420 ;
        RECT  11.440 4.180 11.840 5.420 ;
        RECT  12.900 4.180 13.300 5.420 ;
        RECT  14.360 4.180 14.760 5.420 ;
        RECT  16.570 4.480 16.970 5.420 ;
        RECT  18.630 4.480 19.030 5.420 ;
        RECT  20.930 4.480 21.330 5.420 ;
        RECT  23.230 4.480 23.630 5.420 ;
        RECT  27.130 4.480 27.530 5.420 ;
        RECT  32.640 4.480 33.580 5.420 ;
        RECT  39.170 4.480 39.570 5.420 ;
        RECT  42.990 4.480 43.390 5.420 ;
        RECT  45.260 4.480 45.660 5.420 ;
        RECT  47.430 4.480 47.830 5.420 ;
        RECT  49.570 4.480 49.970 5.420 ;
        RECT  52.050 4.180 52.450 5.420 ;
        RECT  53.510 4.180 53.910 5.420 ;
        RECT  54.970 4.180 55.370 5.420 ;
        RECT  56.430 4.180 56.830 5.420 ;
        RECT  62.450 4.480 62.850 5.420 ;
        RECT  63.750 4.480 64.150 5.420 ;
        RECT  65.240 4.480 66.520 5.420 ;
        RECT  0.000 4.660 66.960 5.420 ;
        RECT  0.440 4.480 1.720 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  57.310 4.180 61.800 4.420 ;
        RECT  50.210 4.180 51.410 4.420 ;
        RECT  51.170 3.580 51.410 4.420 ;
        RECT  66.530 2.520 66.770 4.240 ;
        RECT  48.050 4.000 50.450 4.240 ;
        RECT  61.560 4.000 66.770 4.240 ;
        RECT  57.310 3.580 57.550 4.420 ;
        RECT  51.170 3.580 57.550 3.820 ;
        RECT  66.400 2.520 66.800 2.760 ;
        RECT  65.330 3.060 66.290 3.300 ;
        RECT  65.330 1.340 65.570 3.300 ;
        RECT  65.220 1.920 65.570 2.320 ;
        RECT  65.250 1.340 65.650 1.580 ;
        RECT  61.360 2.060 62.390 2.300 ;
        RECT  65.820 1.880 66.220 2.120 ;
        RECT  61.360 0.620 61.600 2.300 ;
        RECT  65.890 0.800 66.170 2.120 ;
        RECT  61.360 0.800 66.170 1.040 ;
        RECT  51.630 0.800 57.610 1.040 ;
        RECT  50.170 0.720 51.870 0.960 ;
        RECT  57.370 0.620 61.600 0.860 ;
        RECT  61.330 3.030 62.990 3.270 ;
        RECT  62.750 1.580 62.990 3.270 ;
        RECT  62.750 1.900 63.020 2.300 ;
        RECT  61.840 1.580 62.990 1.820 ;
        RECT  61.840 1.300 62.080 1.820 ;
        RECT  51.540 1.500 51.780 1.900 ;
        RECT  57.080 1.600 60.500 1.840 ;
        RECT  51.540 1.570 57.320 1.810 ;
        RECT  60.230 2.620 60.470 3.420 ;
        RECT  58.710 3.100 59.110 3.340 ;
        RECT  51.430 3.100 57.560 3.340 ;
        RECT  57.320 2.620 57.560 3.340 ;
        RECT  58.790 2.620 59.030 3.340 ;
        RECT  57.320 2.620 60.470 2.860 ;
        RECT  50.420 2.980 50.820 3.220 ;
        RECT  50.580 1.680 50.820 3.220 ;
        RECT  50.580 2.620 55.240 2.860 ;
        RECT  54.840 2.530 55.240 2.860 ;
        RECT  50.420 1.680 50.820 1.920 ;
        RECT  50.690 3.520 50.930 3.920 ;
        RECT  48.360 3.520 50.930 3.760 ;
        RECT  48.360 1.680 48.600 3.760 ;
        RECT  48.280 2.980 48.680 3.220 ;
        RECT  48.280 1.680 48.680 1.920 ;
        RECT  49.000 2.980 49.400 3.220 ;
        RECT  49.080 1.680 49.320 3.220 ;
        RECT  49.080 2.320 50.310 2.560 ;
        RECT  49.000 1.680 49.400 1.920 ;
        RECT  46.860 2.980 47.260 3.220 ;
        RECT  46.940 1.680 47.180 3.220 ;
        RECT  47.850 2.240 48.090 2.640 ;
        RECT  46.940 2.320 48.090 2.560 ;
        RECT  46.860 1.680 47.260 1.920 ;
        RECT  42.350 3.520 46.460 3.760 ;
        RECT  46.220 1.680 46.460 3.760 ;
        RECT  42.350 1.680 42.590 3.760 ;
        RECT  46.140 2.980 46.540 3.220 ;
        RECT  44.980 2.440 46.460 2.680 ;
        RECT  46.140 1.680 46.540 1.920 ;
        RECT  42.270 1.680 42.670 1.920 ;
        RECT  40.830 3.220 41.310 3.460 ;
        RECT  41.070 1.200 41.310 3.460 ;
        RECT  43.640 2.980 44.230 3.220 ;
        RECT  43.640 1.200 43.880 3.220 ;
        RECT  40.830 1.680 41.310 1.920 ;
        RECT  43.640 1.440 44.230 1.680 ;
        RECT  41.070 1.200 43.880 1.440 ;
        RECT  42.990 3.040 43.390 3.280 ;
        RECT  43.040 1.680 43.280 3.280 ;
        RECT  42.930 2.240 43.280 2.640 ;
        RECT  42.990 1.680 43.390 1.920 ;
        RECT  40.290 3.700 41.870 3.940 ;
        RECT  41.630 1.680 41.870 3.940 ;
        RECT  39.200 3.520 40.530 3.760 ;
        RECT  39.200 2.710 39.440 3.760 ;
        RECT  41.550 3.220 41.950 3.460 ;
        RECT  39.140 2.710 39.440 3.110 ;
        RECT  41.550 1.680 41.950 1.920 ;
        RECT  37.130 3.120 37.530 3.360 ;
        RECT  40.110 3.040 40.510 3.280 ;
        RECT  37.210 1.100 37.450 3.360 ;
        RECT  40.160 1.540 40.400 3.280 ;
        RECT  40.080 1.580 40.480 1.820 ;
        RECT  39.210 1.540 40.400 1.780 ;
        RECT  39.210 1.100 39.450 1.780 ;
        RECT  37.210 1.100 39.450 1.340 ;
        RECT  38.640 3.360 38.960 3.760 ;
        RECT  38.640 1.580 38.880 3.760 ;
        RECT  39.660 2.040 39.900 2.440 ;
        RECT  38.640 2.120 39.900 2.360 ;
        RECT  38.570 1.580 38.970 1.820 ;
        RECT  35.650 3.600 38.170 3.840 ;
        RECT  37.930 1.580 38.170 3.840 ;
        RECT  35.650 1.500 35.890 3.840 ;
        RECT  37.850 1.580 38.250 1.820 ;
        RECT  36.390 2.880 36.810 3.120 ;
        RECT  36.390 1.580 36.630 3.120 ;
        RECT  36.390 2.140 36.870 2.540 ;
        RECT  36.390 1.580 36.810 1.820 ;
        RECT  34.810 3.040 35.170 3.440 ;
        RECT  34.810 1.100 35.050 3.440 ;
        RECT  32.110 2.310 32.450 2.710 ;
        RECT  32.210 1.100 32.450 2.710 ;
        RECT  34.810 1.500 35.170 1.900 ;
        RECT  32.210 1.100 35.050 1.340 ;
        RECT  28.670 3.600 30.060 3.840 ;
        RECT  34.330 1.580 34.570 3.760 ;
        RECT  29.820 3.520 34.570 3.760 ;
        RECT  34.210 3.040 34.570 3.760 ;
        RECT  28.670 1.580 28.910 3.840 ;
        RECT  28.590 3.040 28.910 3.440 ;
        RECT  34.130 1.580 34.570 1.820 ;
        RECT  28.510 1.580 28.910 1.820 ;
        RECT  33.210 3.040 33.810 3.280 ;
        RECT  33.570 1.580 33.810 3.280 ;
        RECT  33.570 2.320 33.910 2.720 ;
        RECT  33.210 1.580 33.810 1.820 ;
        RECT  29.950 2.970 30.350 3.210 ;
        RECT  30.010 1.580 30.250 3.210 ;
        RECT  29.820 2.330 30.250 2.730 ;
        RECT  29.950 1.580 30.350 1.820 ;
        RECT  29.230 3.120 29.630 3.360 ;
        RECT  26.050 3.040 26.600 3.280 ;
        RECT  29.310 1.500 29.550 3.360 ;
        RECT  26.050 1.490 26.290 3.280 ;
        RECT  29.150 1.100 29.390 1.920 ;
        RECT  26.050 1.490 26.440 1.900 ;
        RECT  26.050 1.490 27.550 1.730 ;
        RECT  27.310 1.100 27.550 1.730 ;
        RECT  27.310 1.100 29.390 1.340 ;
        RECT  27.720 3.520 28.120 3.760 ;
        RECT  27.880 1.580 28.120 3.760 ;
        RECT  26.820 2.040 27.060 2.440 ;
        RECT  26.820 2.040 28.120 2.280 ;
        RECT  27.790 1.580 28.120 2.280 ;
        RECT  27.790 1.580 28.190 1.820 ;
        RECT  24.750 3.700 26.410 3.940 ;
        RECT  27.240 2.710 27.480 3.760 ;
        RECT  26.170 3.520 27.480 3.760 ;
        RECT  24.750 1.680 24.990 3.940 ;
        RECT  24.670 3.220 25.070 3.460 ;
        RECT  27.240 2.710 27.570 3.110 ;
        RECT  24.670 1.680 25.070 1.920 ;
        RECT  25.390 3.220 25.790 3.460 ;
        RECT  22.390 2.980 22.990 3.220 ;
        RECT  22.750 1.200 22.990 3.220 ;
        RECT  25.390 1.200 25.630 3.460 ;
        RECT  25.390 1.680 25.790 1.920 ;
        RECT  22.390 1.440 22.990 1.680 ;
        RECT  22.750 1.200 25.630 1.440 ;
        RECT  20.160 3.520 24.270 3.760 ;
        RECT  24.030 1.680 24.270 3.760 ;
        RECT  20.160 2.980 20.400 3.760 ;
        RECT  20.140 2.980 20.540 3.220 ;
        RECT  20.150 1.680 20.390 3.220 ;
        RECT  20.150 2.440 21.800 2.680 ;
        RECT  23.950 1.680 24.350 1.920 ;
        RECT  20.140 1.680 20.540 1.920 ;
        RECT  23.230 3.040 23.630 3.280 ;
        RECT  23.310 1.680 23.550 3.280 ;
        RECT  23.310 2.240 23.690 2.640 ;
        RECT  23.230 1.680 23.630 1.920 ;
        RECT  19.420 2.980 19.820 3.220 ;
        RECT  19.580 1.680 19.820 3.220 ;
        RECT  18.590 2.240 18.830 2.640 ;
        RECT  18.590 2.320 19.820 2.560 ;
        RECT  19.420 1.680 19.820 1.920 ;
        RECT  5.170 4.180 9.620 4.420 ;
        RECT  9.380 3.580 9.620 4.420 ;
        RECT  15.000 4.000 18.410 4.240 ;
        RECT  0.190 4.000 5.410 4.240 ;
        RECT  15.000 3.580 15.240 4.240 ;
        RECT  0.190 1.800 0.430 4.240 ;
        RECT  9.380 3.580 15.240 3.820 ;
        RECT  0.190 1.800 0.480 2.200 ;
        RECT  15.670 3.520 18.320 3.760 ;
        RECT  18.080 1.680 18.320 3.760 ;
        RECT  18.000 2.980 18.400 3.220 ;
        RECT  18.000 1.680 18.400 1.920 ;
        RECT  17.280 2.980 17.680 3.220 ;
        RECT  17.360 1.680 17.600 3.220 ;
        RECT  16.370 2.320 17.600 2.560 ;
        RECT  17.280 1.680 17.680 1.920 ;
        RECT  0.740 2.520 1.140 2.760 ;
        RECT  0.770 0.800 1.010 2.760 ;
        RECT  4.430 2.070 5.460 2.310 ;
        RECT  5.220 0.620 5.460 2.310 ;
        RECT  9.320 0.800 15.170 1.040 ;
        RECT  0.770 0.800 5.460 1.040 ;
        RECT  14.930 0.720 16.490 0.960 ;
        RECT  5.220 0.620 9.560 0.860 ;
        RECT  15.860 2.980 16.260 3.220 ;
        RECT  15.860 1.680 16.100 3.220 ;
        RECT  11.570 2.560 16.100 2.800 ;
        RECT  11.570 2.530 11.970 2.800 ;
        RECT  15.860 1.680 16.260 1.920 ;
        RECT  6.340 2.620 6.580 3.420 ;
        RECT  9.250 3.100 15.380 3.340 ;
        RECT  7.700 3.100 8.100 3.340 ;
        RECT  9.250 2.620 9.490 3.340 ;
        RECT  7.780 2.620 8.020 3.340 ;
        RECT  6.340 2.620 9.490 2.860 ;
        RECT  14.900 1.440 15.140 1.840 ;
        RECT  6.180 1.600 9.660 1.840 ;
        RECT  9.140 1.570 15.140 1.810 ;
        RECT  3.940 3.030 5.620 3.270 ;
        RECT  3.940 1.380 4.180 3.270 ;
        RECT  3.830 1.960 4.180 2.360 ;
        RECT  4.740 1.300 4.980 1.700 ;
        RECT  3.940 1.380 4.980 1.620 ;
        RECT  0.670 3.060 1.770 3.300 ;
        RECT  1.530 1.340 1.770 3.300 ;
        RECT  1.250 1.340 1.770 1.580 ;
    END
END FACS2P

MACRO FACS2S
    CLASS CORE ;
    FOREIGN FACS2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 49.600 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.280 1.200 7.520 2.320 ;
        RECT  5.100 2.080 7.520 2.320 ;
        RECT  7.280 1.200 12.920 1.440 ;
        RECT  12.680 1.200 12.920 2.200 ;
        RECT  12.680 1.960 14.410 2.200 ;
        RECT  14.010 1.960 14.410 2.220 ;
        RECT  5.130 2.080 5.410 2.860 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  35.350 1.820 36.710 2.100 ;
        RECT  36.470 1.200 36.710 2.100 ;
        RECT  36.470 1.200 42.220 1.440 ;
        RECT  41.980 1.200 42.220 2.320 ;
        RECT  41.980 2.080 44.420 2.320 ;
        RECT  35.040 1.980 35.590 2.220 ;
        END
    END CI0
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.050 2.800 2.360 3.200 ;
        RECT  2.010 1.320 2.410 1.560 ;
        RECT  4.530 1.460 4.770 3.760 ;
        RECT  2.050 3.520 4.770 3.760 ;
        RECT  4.530 1.460 4.860 1.860 ;
        RECT  4.530 3.100 5.100 3.340 ;
        RECT  2.050 1.320 2.290 3.760 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  44.400 3.100 45.070 3.340 ;
        RECT  44.830 1.460 45.070 3.760 ;
        RECT  47.230 2.800 47.550 3.200 ;
        RECT  47.310 1.380 47.550 3.760 ;
        RECT  44.830 3.520 47.550 3.760 ;
        RECT  47.170 1.380 47.570 1.620 ;
        RECT  44.640 1.460 45.070 1.860 ;
        END
    END CO0
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  22.510 1.500 23.010 1.900 ;
        RECT  22.510 3.040 23.090 3.280 ;
        RECT  22.510 1.500 22.750 3.280 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.710 4.000 16.010 4.240 ;
        RECT  15.770 4.180 18.790 4.420 ;
        RECT  18.550 4.000 19.910 4.240 ;
        RECT  20.900 4.080 21.300 4.420 ;
        RECT  19.670 4.180 22.380 4.420 ;
        RECT  22.140 4.000 25.230 4.240 ;
        RECT  22.140 4.060 26.000 4.240 ;
        RECT  26.790 4.080 27.190 4.420 ;
        RECT  24.990 4.180 29.740 4.420 ;
        RECT  29.500 4.000 30.970 4.240 ;
        RECT  30.730 4.180 33.640 4.420 ;
        RECT  33.400 4.000 38.410 4.240 ;
        RECT  10.710 2.840 10.990 4.240 ;
        END
    END B
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  23.730 2.420 24.210 2.820 ;
        RECT  23.730 1.760 24.010 3.080 ;
        END
    END CS
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.210 0.620 13.450 1.720 ;
        RECT  14.170 0.620 14.410 1.200 ;
        RECT  13.210 0.960 14.410 1.200 ;
        RECT  14.170 0.620 18.010 0.860 ;
        RECT  17.770 0.620 18.010 1.250 ;
        RECT  18.730 0.620 18.970 1.250 ;
        RECT  17.770 1.010 18.970 1.250 ;
        RECT  18.730 0.620 21.780 0.860 ;
        RECT  21.540 0.620 21.780 1.130 ;
        RECT  22.680 0.620 22.920 1.130 ;
        RECT  21.540 0.890 22.920 1.130 ;
        RECT  22.680 0.620 26.410 0.860 ;
        RECT  26.170 0.620 26.410 1.130 ;
        RECT  27.130 0.620 27.370 1.130 ;
        RECT  26.170 0.890 27.370 1.130 ;
        RECT  30.610 0.620 31.680 0.980 ;
        RECT  27.130 0.620 31.800 0.860 ;
        RECT  30.610 0.720 35.270 0.960 ;
        RECT  35.030 0.960 36.230 1.200 ;
        RECT  35.990 0.720 40.550 0.960 ;
        RECT  8.950 0.720 13.450 0.960 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.040 -0.380 6.440 0.560 ;
        RECT  13.690 -0.380 13.930 0.640 ;
        RECT  18.250 -0.380 18.490 0.640 ;
        RECT  22.070 -0.380 22.310 0.650 ;
        RECT  26.650 -0.380 26.890 0.650 ;
        RECT  35.510 -0.380 35.750 0.640 ;
        RECT  43.060 -0.380 43.460 0.560 ;
        RECT  46.380 -0.380 46.780 0.560 ;
        RECT  47.980 -0.380 48.380 0.560 ;
        RECT  0.000 -0.380 49.600 0.380 ;
        RECT  1.680 -0.380 3.160 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.850 4.480 3.250 5.420 ;
        RECT  6.260 4.480 6.660 5.420 ;
        RECT  8.390 4.480 8.790 5.420 ;
        RECT  10.690 4.480 11.090 5.420 ;
        RECT  12.830 4.480 13.230 5.420 ;
        RECT  15.130 4.480 15.530 5.420 ;
        RECT  19.030 4.480 19.430 5.420 ;
        RECT  22.680 4.480 24.700 5.420 ;
        RECT  30.090 4.480 30.490 5.420 ;
        RECT  33.910 4.480 34.310 5.420 ;
        RECT  36.180 4.480 36.580 5.420 ;
        RECT  38.570 4.480 38.970 5.420 ;
        RECT  40.710 4.480 41.110 5.420 ;
        RECT  42.840 4.480 43.240 5.420 ;
        RECT  46.350 4.480 46.750 5.420 ;
        RECT  47.880 4.480 49.160 5.420 ;
        RECT  0.000 4.660 49.600 5.420 ;
        RECT  0.440 4.480 1.720 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  39.130 4.000 49.410 4.240 ;
        RECT  49.170 2.520 49.410 4.240 ;
        RECT  49.040 2.520 49.440 2.760 ;
        RECT  47.970 3.060 48.930 3.300 ;
        RECT  47.970 1.340 48.210 3.300 ;
        RECT  47.860 1.860 48.210 2.260 ;
        RECT  47.890 1.340 48.290 1.580 ;
        RECT  45.310 2.070 46.390 2.310 ;
        RECT  48.460 1.880 48.860 2.120 ;
        RECT  45.310 0.720 45.550 2.310 ;
        RECT  48.530 0.800 48.810 2.120 ;
        RECT  45.300 0.800 48.810 1.040 ;
        RECT  42.460 0.800 44.290 1.040 ;
        RECT  44.050 0.720 45.550 0.960 ;
        RECT  41.110 0.720 42.700 0.960 ;
        RECT  45.310 3.030 46.930 3.270 ;
        RECT  46.690 1.590 46.930 3.270 ;
        RECT  46.690 1.840 47.000 2.240 ;
        RECT  45.790 1.590 46.930 1.830 ;
        RECT  45.790 1.300 46.030 1.830 ;
        RECT  42.460 1.440 42.700 1.840 ;
        RECT  42.460 1.540 44.190 1.780 ;
        RECT  42.220 3.100 43.970 3.340 ;
        RECT  41.340 2.980 41.740 3.220 ;
        RECT  41.500 1.680 41.740 3.220 ;
        RECT  41.500 2.560 43.630 2.800 ;
        RECT  41.340 1.680 41.740 1.920 ;
        RECT  39.280 3.520 41.930 3.760 ;
        RECT  39.280 1.680 39.520 3.760 ;
        RECT  39.200 2.980 39.600 3.220 ;
        RECT  39.200 1.680 39.600 1.920 ;
        RECT  39.920 2.980 40.320 3.220 ;
        RECT  39.990 1.680 40.230 3.220 ;
        RECT  39.990 2.280 41.230 2.520 ;
        RECT  39.920 1.680 40.320 1.920 ;
        RECT  37.780 2.980 38.180 3.220 ;
        RECT  37.860 1.680 38.100 3.220 ;
        RECT  38.770 2.200 39.010 2.600 ;
        RECT  37.860 2.280 39.010 2.520 ;
        RECT  37.780 1.680 38.180 1.920 ;
        RECT  33.270 3.520 37.380 3.760 ;
        RECT  37.140 1.680 37.380 3.760 ;
        RECT  33.270 1.680 33.510 3.760 ;
        RECT  37.060 2.980 37.460 3.220 ;
        RECT  35.720 2.440 37.380 2.680 ;
        RECT  37.060 1.680 37.460 1.920 ;
        RECT  33.190 1.680 33.590 1.920 ;
        RECT  31.750 3.220 32.230 3.460 ;
        RECT  31.990 1.200 32.230 3.460 ;
        RECT  34.550 2.980 35.150 3.220 ;
        RECT  34.550 1.200 34.790 3.220 ;
        RECT  31.750 1.680 32.230 1.920 ;
        RECT  34.550 1.440 35.150 1.680 ;
        RECT  31.990 1.200 34.790 1.440 ;
        RECT  33.910 3.040 34.310 3.280 ;
        RECT  33.960 1.680 34.200 3.280 ;
        RECT  33.850 2.240 34.200 2.640 ;
        RECT  33.910 1.680 34.310 1.920 ;
        RECT  31.210 3.700 32.790 3.940 ;
        RECT  32.550 1.680 32.790 3.940 ;
        RECT  30.120 3.520 31.450 3.760 ;
        RECT  30.120 2.710 30.360 3.760 ;
        RECT  32.470 3.220 32.870 3.460 ;
        RECT  30.060 2.710 30.360 3.110 ;
        RECT  32.470 1.680 32.870 1.920 ;
        RECT  28.050 3.120 28.450 3.360 ;
        RECT  31.030 3.040 31.430 3.280 ;
        RECT  28.130 1.100 28.370 3.360 ;
        RECT  31.080 1.490 31.320 3.280 ;
        RECT  30.130 1.490 31.320 1.730 ;
        RECT  30.130 1.100 30.370 1.730 ;
        RECT  28.130 1.100 30.370 1.340 ;
        RECT  29.560 3.360 29.880 3.760 ;
        RECT  29.560 1.580 29.800 3.760 ;
        RECT  30.600 2.040 30.840 2.440 ;
        RECT  29.560 2.120 30.840 2.360 ;
        RECT  29.490 1.580 29.890 1.820 ;
        RECT  26.570 3.600 29.090 3.840 ;
        RECT  28.850 1.580 29.090 3.840 ;
        RECT  26.570 1.500 26.810 3.840 ;
        RECT  28.770 1.580 29.170 1.820 ;
        RECT  27.310 2.880 27.730 3.120 ;
        RECT  27.310 1.580 27.550 3.120 ;
        RECT  27.310 2.140 27.790 2.540 ;
        RECT  27.310 1.580 27.730 1.820 ;
        RECT  25.690 3.040 26.090 3.440 ;
        RECT  25.690 1.100 25.930 3.440 ;
        RECT  23.250 1.100 23.490 2.440 ;
        RECT  25.690 1.500 26.090 1.900 ;
        RECT  23.250 1.100 25.930 1.340 ;
        RECT  20.570 3.600 21.960 3.840 ;
        RECT  25.150 1.580 25.390 3.760 ;
        RECT  21.720 3.520 25.390 3.760 ;
        RECT  25.130 3.040 25.390 3.760 ;
        RECT  20.570 1.580 20.810 3.840 ;
        RECT  20.490 3.040 20.810 3.440 ;
        RECT  25.050 1.580 25.450 1.820 ;
        RECT  20.410 1.580 20.810 1.820 ;
        RECT  24.330 3.040 24.810 3.280 ;
        RECT  24.570 1.580 24.810 3.280 ;
        RECT  24.570 2.320 24.910 2.720 ;
        RECT  24.330 1.580 24.810 1.820 ;
        RECT  21.850 2.970 22.250 3.210 ;
        RECT  21.910 1.580 22.150 3.210 ;
        RECT  21.720 2.330 22.150 2.730 ;
        RECT  21.850 1.580 22.250 1.820 ;
        RECT  21.130 3.120 21.530 3.360 ;
        RECT  17.950 3.040 18.500 3.280 ;
        RECT  21.210 1.500 21.450 3.360 ;
        RECT  17.950 1.490 18.190 3.280 ;
        RECT  21.050 1.100 21.290 1.920 ;
        RECT  17.950 1.490 18.340 1.900 ;
        RECT  17.950 1.490 19.450 1.730 ;
        RECT  19.210 1.100 19.450 1.730 ;
        RECT  19.210 1.100 21.290 1.340 ;
        RECT  19.620 3.520 20.020 3.760 ;
        RECT  19.780 1.580 20.020 3.760 ;
        RECT  18.720 2.040 18.960 2.440 ;
        RECT  18.720 2.040 20.020 2.280 ;
        RECT  19.690 1.580 20.020 2.280 ;
        RECT  19.690 1.580 20.090 1.820 ;
        RECT  16.650 3.700 18.310 3.940 ;
        RECT  19.140 2.710 19.380 3.760 ;
        RECT  18.070 3.520 19.380 3.760 ;
        RECT  16.650 1.680 16.890 3.940 ;
        RECT  16.570 3.220 16.970 3.460 ;
        RECT  19.140 2.710 19.470 3.110 ;
        RECT  16.570 1.680 16.970 1.920 ;
        RECT  17.290 3.220 17.690 3.460 ;
        RECT  14.290 2.980 14.890 3.220 ;
        RECT  14.650 1.200 14.890 3.220 ;
        RECT  17.290 1.200 17.530 3.460 ;
        RECT  17.290 1.680 17.690 1.920 ;
        RECT  14.290 1.440 14.890 1.680 ;
        RECT  14.650 1.200 17.530 1.440 ;
        RECT  12.060 3.520 16.170 3.760 ;
        RECT  15.930 1.680 16.170 3.760 ;
        RECT  12.060 2.980 12.300 3.760 ;
        RECT  12.040 2.980 12.440 3.220 ;
        RECT  12.050 1.680 12.290 3.220 ;
        RECT  12.050 2.440 13.700 2.680 ;
        RECT  15.850 1.680 16.250 1.920 ;
        RECT  12.040 1.680 12.440 1.920 ;
        RECT  15.130 3.040 15.530 3.280 ;
        RECT  15.210 1.680 15.450 3.280 ;
        RECT  15.210 2.240 15.590 2.640 ;
        RECT  15.130 1.680 15.530 1.920 ;
        RECT  11.320 2.980 11.720 3.220 ;
        RECT  11.400 1.680 11.640 3.220 ;
        RECT  10.490 2.200 10.730 2.600 ;
        RECT  10.490 2.280 11.640 2.520 ;
        RECT  11.320 1.680 11.720 1.920 ;
        RECT  0.190 4.000 10.470 4.240 ;
        RECT  0.190 1.800 0.430 4.240 ;
        RECT  0.190 1.800 0.480 2.200 ;
        RECT  7.570 3.520 10.220 3.760 ;
        RECT  9.980 1.680 10.220 3.760 ;
        RECT  9.900 2.980 10.300 3.220 ;
        RECT  9.900 1.680 10.300 1.920 ;
        RECT  9.180 2.980 9.580 3.220 ;
        RECT  9.260 1.680 9.500 3.220 ;
        RECT  8.350 2.200 8.590 2.600 ;
        RECT  8.350 2.280 9.500 2.520 ;
        RECT  9.180 1.680 9.580 1.920 ;
        RECT  0.740 2.520 1.140 2.760 ;
        RECT  0.770 0.800 1.010 2.760 ;
        RECT  3.210 2.070 4.290 2.310 ;
        RECT  4.050 0.620 4.290 2.310 ;
        RECT  5.130 0.800 6.960 1.040 ;
        RECT  0.770 0.800 4.290 1.040 ;
        RECT  6.720 0.720 8.390 0.960 ;
        RECT  4.050 0.620 5.370 0.860 ;
        RECT  7.760 2.980 8.160 3.220 ;
        RECT  7.760 1.680 8.000 3.220 ;
        RECT  5.870 2.560 8.000 2.800 ;
        RECT  7.760 1.680 8.160 1.920 ;
        RECT  5.530 3.100 7.280 3.340 ;
        RECT  6.800 1.440 7.040 1.840 ;
        RECT  5.310 1.540 7.040 1.780 ;
        RECT  2.670 3.030 4.280 3.270 ;
        RECT  2.670 1.320 2.910 3.270 ;
        RECT  2.570 1.840 2.910 2.240 ;
        RECT  2.670 1.320 3.810 1.560 ;
        RECT  0.670 3.060 1.770 3.300 ;
        RECT  1.530 1.340 1.770 3.300 ;
        RECT  1.250 1.340 1.770 1.580 ;
    END
END FACS2S

MACRO FILLER1
    CLASS CORE SPACER ;
    FOREIGN FILLER1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.620 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 0.620 0.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 0.620 5.420 ;
        END
    END VCC
END FILLER1

MACRO FILLER16
    CLASS CORE SPACER ;
    FOREIGN FILLER16 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 9.920 0.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 9.920 5.420 ;
        END
    END VCC
END FILLER16

MACRO FILLER2
    CLASS CORE SPACER ;
    FOREIGN FILLER2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.240 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.240 0.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 1.240 5.420 ;
        END
    END VCC
END FILLER2

MACRO FILLER2C
    CLASS CORE SPACER ;
    FOREIGN FILLER2C 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.240 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.240 0.380 ;
        RECT  0.140 -0.380 0.580 2.530 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 1.240 5.420 ;
        RECT  0.430 2.770 0.870 5.420 ;
        END
    END VCC
END FILLER2C

MACRO FILLER32
    CLASS CORE SPACER ;
    FOREIGN FILLER32 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.840 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 19.840 0.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 19.840 5.420 ;
        END
    END VCC
END FILLER32

MACRO FILLER4
    CLASS CORE SPACER ;
    FOREIGN FILLER4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 2.480 5.420 ;
        END
    END VCC
END FILLER4

MACRO FILLER4C
    CLASS CORE SPACER ;
    FOREIGN FILLER4C 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.140 -0.380 2.340 1.130 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.140 -0.380 0.500 2.650 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.140 3.910 2.340 5.420 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  1.980 1.850 2.340 5.420 ;
        END
    END VCC
END FILLER4C

MACRO FILLER64
    CLASS CORE SPACER ;
    FOREIGN FILLER64 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 39.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 39.680 0.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 39.680 5.420 ;
        END
    END VCC
END FILLER64

MACRO FILLER8
    CLASS CORE SPACER ;
    FOREIGN FILLER8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 4.960 5.420 ;
        END
    END VCC
END FILLER8

MACRO FILLER8C
    CLASS CORE SPACER ;
    FOREIGN FILLER8C 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.730 -0.380 1.130 0.870 ;
        RECT  3.830 -0.380 4.230 0.870 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.190 -0.380 1.130 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.830 4.170 4.230 5.420 ;
        RECT  3.830 4.480 4.770 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.730 4.170 1.130 5.420 ;
        END
    END VCC
END FILLER8C

MACRO FILLERAC
    CLASS CORE SPACER ;
    FOREIGN FILLERAC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.730 -0.380 1.130 0.870 ;
        RECT  8.790 -0.380 9.190 0.870 ;
        RECT  0.000 -0.380 9.920 0.380 ;
        RECT  0.190 -0.380 1.130 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  8.790 4.170 9.190 5.420 ;
        RECT  8.790 4.480 9.730 5.420 ;
        RECT  0.000 4.660 9.920 5.420 ;
        RECT  0.730 4.170 1.130 5.420 ;
        END
    END VCC
END FILLERAC

MACRO FILLERBC
    CLASS CORE SPACER ;
    FOREIGN FILLERBC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.840 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.730 -0.380 1.130 0.870 ;
        RECT  9.410 -0.380 9.810 0.870 ;
        RECT  18.710 -0.380 19.110 0.870 ;
        RECT  18.710 -0.380 19.650 0.560 ;
        RECT  0.000 -0.380 19.840 0.380 ;
        RECT  0.190 -0.380 1.130 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  10.030 3.860 10.430 5.420 ;
        RECT  9.530 4.480 10.430 5.420 ;
        RECT  18.710 4.170 19.110 5.420 ;
        RECT  0.000 4.660 19.840 5.420 ;
        RECT  0.720 4.170 1.120 5.420 ;
        END
    END VCC
END FILLERBC

MACRO FILLERCC
    CLASS CORE SPACER ;
    FOREIGN FILLERCC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 39.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.730 -0.380 1.130 0.870 ;
        RECT  10.030 -0.380 10.430 0.870 ;
        RECT  18.830 -0.380 19.730 0.560 ;
        RECT  19.330 -0.380 19.730 1.180 ;
        RECT  29.250 -0.380 29.650 0.870 ;
        RECT  38.550 -0.380 38.950 0.880 ;
        RECT  38.550 -0.380 39.490 0.570 ;
        RECT  0.000 -0.380 39.680 0.380 ;
        RECT  0.190 -0.380 1.130 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  10.030 3.860 10.430 5.420 ;
        RECT  9.530 4.480 10.430 5.420 ;
        RECT  19.940 4.170 20.340 5.420 ;
        RECT  29.310 3.860 29.710 5.420 ;
        RECT  28.810 4.480 29.710 5.420 ;
        RECT  38.550 4.170 38.950 5.420 ;
        RECT  0.000 4.660 39.680 5.420 ;
        RECT  0.730 4.170 1.130 5.420 ;
        END
    END VCC
END FILLERCC

MACRO GCKETF
    CLASS CORE ;
    FOREIGN GCKETF 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.010 1.600 11.230 1.840 ;
        RECT  10.990 1.600 11.230 2.500 ;
        RECT  10.990 2.100 11.260 2.500 ;
        RECT  7.010 1.600 7.250 2.180 ;
        END
    END CK
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.110 2.080 10.350 2.890 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 2.230 0.480 2.630 ;
        RECT  0.190 2.180 0.430 2.860 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.940 1.490 13.180 4.090 ;
        RECT  12.860 3.150 13.180 4.090 ;
        RECT  14.300 1.200 14.690 1.600 ;
        RECT  12.940 2.280 14.690 2.760 ;
        RECT  14.450 1.200 14.690 4.090 ;
        RECT  14.300 3.150 14.690 4.090 ;
        RECT  12.860 1.490 13.180 1.890 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.160 -0.380 3.560 0.560 ;
        RECT  6.450 -0.380 6.850 0.570 ;
        RECT  8.660 -0.380 9.060 0.570 ;
        RECT  10.080 -0.380 10.480 0.570 ;
        RECT  13.580 -0.380 13.820 1.050 ;
        RECT  15.020 -0.380 15.260 1.050 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.810 4.480 4.210 5.420 ;
        RECT  5.900 4.480 6.300 5.420 ;
        RECT  7.040 4.480 7.440 5.420 ;
        RECT  9.710 4.260 10.110 5.420 ;
        RECT  10.620 3.930 11.020 5.420 ;
        RECT  12.140 2.890 12.380 5.420 ;
        RECT  13.580 3.620 13.820 5.420 ;
        RECT  15.020 3.620 15.260 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.760 3.970 9.210 4.210 ;
        RECT  8.970 3.390 9.210 4.210 ;
        RECT  8.970 3.390 11.790 3.630 ;
        RECT  11.550 1.480 11.790 3.630 ;
        RECT  11.550 2.230 12.700 2.630 ;
        RECT  11.470 1.480 11.870 1.720 ;
        RECT  10.750 1.000 11.150 1.360 ;
        RECT  9.290 1.000 9.690 1.360 ;
        RECT  7.870 1.000 8.270 1.360 ;
        RECT  7.870 1.000 12.670 1.240 ;
        RECT  12.270 0.850 12.670 1.240 ;
        RECT  4.950 3.590 5.290 3.990 ;
        RECT  5.050 1.560 5.290 3.990 ;
        RECT  8.320 2.100 8.560 3.720 ;
        RECT  5.050 3.480 8.560 3.720 ;
        RECT  3.020 1.560 5.290 1.800 ;
        RECT  6.230 2.870 7.640 3.110 ;
        RECT  6.230 1.080 6.470 3.110 ;
        RECT  3.130 1.080 7.550 1.320 ;
        RECT  1.350 0.850 3.370 1.090 ;
        RECT  5.740 1.560 5.980 3.210 ;
        RECT  5.550 2.230 5.980 2.630 ;
        RECT  5.530 1.560 5.980 1.800 ;
        RECT  1.350 4.060 3.650 4.300 ;
        RECT  4.380 2.230 4.620 4.130 ;
        RECT  3.410 3.890 4.620 4.130 ;
        RECT  2.620 2.340 4.620 2.580 ;
        RECT  1.660 3.580 3.170 3.820 ;
        RECT  3.800 2.960 4.040 3.650 ;
        RECT  2.930 3.410 4.040 3.650 ;
        RECT  1.660 1.330 1.900 3.820 ;
        RECT  2.140 2.940 2.690 3.340 ;
        RECT  2.140 1.410 2.380 3.340 ;
        RECT  2.140 1.410 2.700 1.650 ;
        RECT  0.870 1.310 1.110 3.520 ;
    END
END GCKETF

MACRO GCKETN
    CLASS CORE ;
    FOREIGN GCKETN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.010 1.560 10.080 1.800 ;
        RECT  9.840 1.560 10.080 2.450 ;
        RECT  7.010 1.560 7.250 2.180 ;
        END
    END CK
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.860 2.290 9.220 2.890 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 2.320 0.480 2.720 ;
        RECT  0.190 2.180 0.430 2.860 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.970 1.280 12.210 4.090 ;
        RECT  11.920 3.150 12.210 4.090 ;
        RECT  11.920 1.280 12.210 1.680 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.350 -0.380 3.750 0.560 ;
        RECT  6.410 -0.380 6.810 0.620 ;
        RECT  8.780 -0.380 9.180 0.570 ;
        RECT  11.200 -0.380 11.440 1.680 ;
        RECT  0.000 -0.380 12.400 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.130 4.480 4.530 5.420 ;
        RECT  5.860 4.480 6.260 5.420 ;
        RECT  7.000 4.480 7.400 5.420 ;
        RECT  9.410 4.000 9.810 5.420 ;
        RECT  11.200 3.620 11.440 5.420 ;
        RECT  0.000 4.660 12.400 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.920 3.970 9.110 4.210 ;
        RECT  8.870 3.520 9.110 4.210 ;
        RECT  10.320 3.520 10.560 3.980 ;
        RECT  8.870 3.520 10.720 3.760 ;
        RECT  10.480 0.810 10.720 3.760 ;
        RECT  10.480 2.230 10.880 2.630 ;
        RECT  7.920 1.080 9.970 1.320 ;
        RECT  5.200 3.480 5.440 4.120 ;
        RECT  4.990 3.480 8.360 3.720 ;
        RECT  8.120 2.590 8.360 3.720 ;
        RECT  4.990 1.560 5.230 3.720 ;
        RECT  3.180 1.560 5.230 1.800 ;
        RECT  6.190 2.870 7.600 3.110 ;
        RECT  6.190 1.080 6.430 3.110 ;
        RECT  3.290 1.080 7.600 1.320 ;
        RECT  1.510 0.850 3.530 1.090 ;
        RECT  5.700 1.560 5.940 3.210 ;
        RECT  5.510 2.230 5.940 2.630 ;
        RECT  5.490 1.560 5.940 1.800 ;
        RECT  1.510 4.060 3.810 4.300 ;
        RECT  4.500 2.230 4.740 4.130 ;
        RECT  3.570 3.890 4.740 4.130 ;
        RECT  2.780 2.340 4.740 2.580 ;
        RECT  1.820 3.580 3.330 3.820 ;
        RECT  4.020 3.230 4.260 3.650 ;
        RECT  3.090 3.410 4.260 3.650 ;
        RECT  1.820 1.330 2.060 3.820 ;
        RECT  2.300 2.940 2.850 3.340 ;
        RECT  2.300 1.410 2.540 3.340 ;
        RECT  2.300 1.410 2.860 1.650 ;
        RECT  1.030 1.310 1.270 3.520 ;
    END
END GCKETN

MACRO GCKETP
    CLASS CORE ;
    FOREIGN GCKETP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.010 1.560 10.080 1.800 ;
        RECT  9.840 1.560 10.080 2.860 ;
        RECT  7.010 1.560 7.250 2.180 ;
        END
    END CK
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.870 2.310 9.220 2.710 ;
        RECT  8.870 2.290 9.110 2.890 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 2.230 0.480 2.630 ;
        RECT  0.190 2.180 0.430 2.860 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.970 1.490 12.210 4.090 ;
        RECT  11.820 3.150 12.210 4.090 ;
        RECT  11.820 1.490 12.210 1.890 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.350 -0.380 3.750 0.560 ;
        RECT  6.410 -0.380 6.810 0.620 ;
        RECT  8.710 -0.380 9.110 0.570 ;
        RECT  11.040 -0.380 11.280 1.910 ;
        RECT  11.040 1.490 11.340 1.890 ;
        RECT  12.540 -0.380 12.780 1.800 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.130 4.480 4.530 5.420 ;
        RECT  5.860 4.480 6.260 5.420 ;
        RECT  7.000 4.480 7.400 5.420 ;
        RECT  9.220 4.260 9.620 5.420 ;
        RECT  11.100 2.790 11.340 5.420 ;
        RECT  12.540 3.620 12.780 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.920 3.970 8.850 4.210 ;
        RECT  8.610 3.520 8.850 4.210 ;
        RECT  10.320 3.520 10.560 3.980 ;
        RECT  8.610 3.520 10.720 3.760 ;
        RECT  10.480 0.810 10.720 3.760 ;
        RECT  10.480 2.230 10.820 2.630 ;
        RECT  7.920 1.080 9.970 1.320 ;
        RECT  5.200 3.480 5.440 4.120 ;
        RECT  4.990 3.480 8.360 3.720 ;
        RECT  8.120 2.690 8.360 3.720 ;
        RECT  4.990 1.560 5.230 3.720 ;
        RECT  3.180 1.560 5.230 1.800 ;
        RECT  6.190 2.870 7.600 3.110 ;
        RECT  6.190 1.080 6.430 3.110 ;
        RECT  3.290 1.080 7.600 1.320 ;
        RECT  1.510 0.850 3.530 1.090 ;
        RECT  5.700 1.560 5.940 3.210 ;
        RECT  5.510 2.230 5.940 2.630 ;
        RECT  5.490 1.560 5.940 1.800 ;
        RECT  1.510 4.060 3.810 4.300 ;
        RECT  4.500 2.230 4.740 4.130 ;
        RECT  3.570 3.890 4.740 4.130 ;
        RECT  2.780 2.340 4.740 2.580 ;
        RECT  1.820 3.580 3.330 3.820 ;
        RECT  4.020 3.230 4.260 3.650 ;
        RECT  3.090 3.410 4.260 3.650 ;
        RECT  1.820 1.330 2.060 3.820 ;
        RECT  2.300 2.940 2.850 3.340 ;
        RECT  2.300 1.410 2.540 3.340 ;
        RECT  2.300 1.410 2.860 1.650 ;
        RECT  1.030 1.310 1.270 3.520 ;
    END
END GCKETP

MACRO GCKETT
    CLASS CORE ;
    FOREIGN GCKETT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.010 1.600 11.250 1.840 ;
        RECT  11.010 1.600 11.250 2.500 ;
        RECT  11.010 2.100 11.280 2.500 ;
        RECT  7.010 1.600 7.250 2.180 ;
        END
    END CK
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.490 2.100 9.820 2.500 ;
        RECT  9.490 2.080 9.730 2.890 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 2.230 0.480 2.630 ;
        RECT  0.190 2.180 0.430 2.860 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.400 1.200 14.690 1.600 ;
        RECT  12.960 2.400 14.690 2.640 ;
        RECT  14.450 1.200 14.690 4.090 ;
        RECT  14.400 3.150 14.690 4.090 ;
        RECT  12.960 1.490 13.200 4.090 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.160 -0.380 3.560 0.560 ;
        RECT  6.190 -0.380 6.590 0.570 ;
        RECT  8.400 -0.380 8.800 0.570 ;
        RECT  9.980 -0.380 10.380 0.570 ;
        RECT  13.680 -0.380 13.920 0.890 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.910 4.480 4.310 5.420 ;
        RECT  5.640 4.480 6.040 5.420 ;
        RECT  6.780 4.480 7.180 5.420 ;
        RECT  10.010 4.260 10.410 5.420 ;
        RECT  12.240 2.890 12.480 5.420 ;
        RECT  13.680 3.620 13.920 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.170 3.270 11.410 4.210 ;
        RECT  7.860 3.970 9.710 4.210 ;
        RECT  9.470 3.270 9.710 4.210 ;
        RECT  9.470 3.270 11.810 3.510 ;
        RECT  11.570 1.480 11.810 3.510 ;
        RECT  11.570 2.230 12.720 2.630 ;
        RECT  11.490 1.480 11.890 1.720 ;
        RECT  10.770 1.000 11.170 1.360 ;
        RECT  9.190 1.000 9.590 1.360 ;
        RECT  7.610 1.000 8.010 1.360 ;
        RECT  7.610 1.000 12.690 1.240 ;
        RECT  12.290 0.870 12.690 1.240 ;
        RECT  4.980 3.480 5.220 4.120 ;
        RECT  4.770 3.480 8.300 3.720 ;
        RECT  8.060 2.100 8.300 3.720 ;
        RECT  4.770 1.560 5.010 3.720 ;
        RECT  3.020 1.560 5.010 1.800 ;
        RECT  5.970 2.870 7.380 3.110 ;
        RECT  5.970 1.080 6.210 3.110 ;
        RECT  3.130 1.080 7.290 1.320 ;
        RECT  1.350 0.850 3.370 1.090 ;
        RECT  5.480 1.560 5.720 3.210 ;
        RECT  5.290 2.230 5.720 2.630 ;
        RECT  5.270 1.560 5.720 1.800 ;
        RECT  1.350 4.060 3.660 4.300 ;
        RECT  4.280 2.230 4.520 4.130 ;
        RECT  3.420 3.890 4.520 4.130 ;
        RECT  2.620 2.340 4.520 2.580 ;
        RECT  1.660 3.580 3.170 3.820 ;
        RECT  3.800 2.960 4.040 3.650 ;
        RECT  2.930 3.410 4.040 3.650 ;
        RECT  1.660 1.330 1.900 3.820 ;
        RECT  2.140 2.940 2.690 3.340 ;
        RECT  2.140 1.410 2.380 3.340 ;
        RECT  2.140 1.410 2.700 1.650 ;
        RECT  0.870 1.310 1.110 3.520 ;
    END
END GCKETT

MACRO HA1
    CLASS CORE ;
    FOREIGN HA1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.060 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 1.180 6.650 3.300 ;
        RECT  6.180 2.900 6.650 3.300 ;
        RECT  6.190 1.460 6.650 1.860 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.610 0.630 7.890 3.260 ;
        RECT  7.570 2.860 7.890 3.260 ;
        RECT  7.570 1.240 7.890 1.640 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.280 1.070 2.840 ;
        RECT  0.790 1.280 1.550 1.520 ;
        RECT  2.310 1.100 2.550 3.840 ;
        RECT  2.310 3.440 2.610 3.840 ;
        RECT  1.310 1.100 4.260 1.340 ;
        RECT  4.020 1.100 4.260 3.200 ;
        RECT  5.150 2.170 5.390 3.200 ;
        RECT  4.020 2.960 5.390 3.200 ;
        RECT  5.150 2.170 5.460 2.570 ;
        RECT  0.740 2.200 1.070 2.600 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 0.620 4.790 2.550 ;
        RECT  2.440 0.620 4.790 0.860 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.050 -0.380 5.450 0.560 ;
        RECT  6.900 -0.380 7.270 0.940 ;
        RECT  0.000 -0.380 8.060 0.380 ;
        RECT  0.720 -0.380 1.120 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 3.080 1.540 5.420 ;
        RECT  4.660 4.470 5.580 5.420 ;
        RECT  6.870 4.090 7.290 5.420 ;
        RECT  0.000 4.660 8.060 5.420 ;
        RECT  1.060 3.080 1.540 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.530 3.990 6.630 4.230 ;
        RECT  6.390 3.580 6.630 4.230 ;
        RECT  4.530 3.520 4.770 4.230 ;
        RECT  6.390 3.580 7.250 3.820 ;
        RECT  7.010 2.140 7.250 3.820 ;
        RECT  2.940 3.520 4.770 3.760 ;
        RECT  2.940 1.580 3.180 3.760 ;
        RECT  2.810 2.880 3.180 3.280 ;
        RECT  7.010 2.140 7.370 2.540 ;
        RECT  2.790 1.580 3.180 1.980 ;
        RECT  5.070 3.450 5.940 3.690 ;
        RECT  5.700 0.850 5.940 3.690 ;
        RECT  5.410 0.850 5.940 1.800 ;
        RECT  1.830 4.180 3.230 4.420 ;
        RECT  3.690 4.020 4.090 4.320 ;
        RECT  2.990 4.080 4.090 4.320 ;
        RECT  1.830 1.580 2.070 4.420 ;
        RECT  3.510 2.880 3.770 3.280 ;
        RECT  3.510 1.580 3.750 3.280 ;
        RECT  0.190 4.080 1.000 4.320 ;
        RECT  0.190 1.490 0.430 4.320 ;
        RECT  0.190 2.880 0.480 3.280 ;
        RECT  0.190 1.490 0.480 1.890 ;
    END
END HA1

MACRO HA1P
    CLASS CORE ;
    FOREIGN HA1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.300 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 0.620 7.270 3.300 ;
        RECT  6.960 2.900 7.270 3.300 ;
        RECT  6.960 1.460 7.270 1.860 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.120 1.260 9.130 1.540 ;
        RECT  8.850 1.260 9.130 3.220 ;
        RECT  8.120 2.940 9.130 3.220 ;
        RECT  8.120 1.260 8.520 1.600 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.390 0.850 1.890 1.130 ;
        RECT  2.410 0.700 2.650 3.750 ;
        RECT  1.610 0.700 3.600 0.980 ;
        RECT  3.200 0.700 3.600 1.150 ;
        RECT  0.790 0.850 1.070 1.780 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.780 1.690 2.880 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.290 -0.380 4.670 1.900 ;
        RECT  6.240 -0.380 6.660 0.930 ;
        RECT  7.510 -0.380 7.900 0.940 ;
        RECT  8.740 -0.380 9.140 0.960 ;
        RECT  0.000 -0.380 9.300 0.380 ;
        RECT  0.960 -0.380 1.360 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 3.150 1.540 5.420 ;
        RECT  4.610 4.000 5.020 5.420 ;
        RECT  6.220 4.090 6.620 5.420 ;
        RECT  7.500 4.090 7.920 5.420 ;
        RECT  8.770 4.100 9.140 5.420 ;
        RECT  0.000 4.660 9.300 5.420 ;
        RECT  1.060 3.150 1.540 3.550 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.390 3.580 7.870 3.820 ;
        RECT  7.630 2.400 7.870 3.820 ;
        RECT  2.960 3.520 6.630 3.760 ;
        RECT  2.960 1.490 3.200 3.760 ;
        RECT  7.630 2.400 8.290 2.640 ;
        RECT  7.890 2.280 8.290 2.640 ;
        RECT  2.890 1.490 3.200 1.890 ;
        RECT  5.150 3.010 5.870 3.250 ;
        RECT  5.150 1.570 5.390 3.250 ;
        RECT  5.150 2.400 6.740 2.640 ;
        RECT  6.500 2.200 6.740 2.640 ;
        RECT  5.000 1.570 5.400 1.810 ;
        RECT  1.930 4.080 4.260 4.320 ;
        RECT  3.860 4.020 4.260 4.320 ;
        RECT  1.930 1.490 2.170 4.320 ;
        RECT  3.710 1.490 3.950 3.190 ;
        RECT  3.610 1.490 3.950 1.890 ;
        RECT  0.190 4.080 1.060 4.320 ;
        RECT  0.190 1.490 0.430 4.320 ;
        RECT  0.190 2.790 0.480 3.190 ;
        RECT  0.190 1.490 0.480 1.890 ;
    END
END HA1P

MACRO HA1S
    CLASS CORE ;
    FOREIGN HA1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.060 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.000 3.540 6.460 3.940 ;
        RECT  6.370 1.470 6.650 3.220 ;
        RECT  6.180 2.940 6.460 3.940 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.610 1.160 7.890 3.830 ;
        RECT  7.570 3.430 7.890 3.830 ;
        RECT  7.150 1.160 7.890 1.400 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.670 2.200 1.070 2.600 ;
        RECT  2.350 1.100 2.590 3.840 ;
        RECT  0.790 1.100 4.270 1.340 ;
        RECT  4.030 1.100 4.270 2.840 ;
        RECT  4.030 2.600 5.270 2.840 ;
        RECT  5.030 2.340 5.460 2.740 ;
        RECT  0.790 0.620 1.070 2.600 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 0.620 4.790 2.350 ;
        RECT  2.100 0.620 4.790 0.860 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.070 -0.380 5.430 1.010 ;
        RECT  6.280 -0.380 6.650 1.150 ;
        RECT  6.280 -0.380 7.590 0.660 ;
        RECT  0.000 -0.380 8.060 0.380 ;
        RECT  1.310 -0.380 1.710 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.200 2.960 1.440 5.420 ;
        RECT  4.250 4.080 4.670 5.420 ;
        RECT  4.250 4.230 5.180 5.420 ;
        RECT  7.190 4.380 7.530 5.420 ;
        RECT  0.000 4.660 8.060 5.420 ;
        RECT  0.960 2.880 1.200 3.280 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.510 4.180 6.940 4.420 ;
        RECT  6.700 3.520 6.940 4.420 ;
        RECT  5.510 3.580 5.750 4.420 ;
        RECT  4.600 3.580 5.750 3.820 ;
        RECT  6.890 2.740 7.130 3.760 ;
        RECT  2.830 3.520 4.840 3.760 ;
        RECT  2.830 1.580 3.070 3.760 ;
        RECT  6.890 2.740 7.320 3.140 ;
        RECT  5.070 3.100 5.710 3.340 ;
        RECT  5.700 0.830 5.940 3.260 ;
        RECT  5.470 3.020 5.940 3.260 ;
        RECT  5.470 1.380 5.940 1.780 ;
        RECT  5.700 0.830 6.030 1.230 ;
        RECT  1.870 4.180 3.410 4.420 ;
        RECT  3.560 4.020 3.960 4.320 ;
        RECT  3.170 4.080 3.960 4.320 ;
        RECT  1.870 1.580 2.110 4.420 ;
        RECT  3.550 1.580 3.790 3.280 ;
        RECT  0.720 3.520 0.960 4.370 ;
        RECT  0.190 3.520 0.960 3.760 ;
        RECT  0.190 0.700 0.430 3.760 ;
        RECT  0.190 2.880 0.480 3.280 ;
        RECT  0.190 0.700 0.480 1.100 ;
    END
END HA1S

MACRO HA1T
    CLASS CORE ;
    FOREIGN HA1T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.880 1.440 8.520 1.680 ;
        RECT  6.880 2.980 8.520 3.220 ;
        RECT  6.990 0.620 7.270 3.300 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.360 1.320 11.000 1.600 ;
        RECT  9.360 2.940 11.000 3.220 ;
        RECT  10.090 1.320 10.370 3.220 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 0.810 1.070 1.720 ;
        RECT  0.400 0.810 1.900 1.090 ;
        RECT  2.410 0.700 2.650 3.750 ;
        RECT  1.620 0.700 3.600 0.980 ;
        RECT  3.200 0.700 3.600 1.150 ;
        RECT  0.400 0.810 1.070 1.150 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.840 ;
        RECT  1.360 2.200 1.690 2.600 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.290 -0.380 4.670 1.900 ;
        RECT  6.240 -0.380 6.660 0.930 ;
        RECT  7.510 -0.380 7.900 0.940 ;
        RECT  8.740 -0.380 9.140 0.960 ;
        RECT  9.980 -0.380 10.380 0.960 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.960 -0.380 1.360 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 3.150 1.540 5.420 ;
        RECT  4.610 4.000 5.020 5.420 ;
        RECT  6.220 4.090 6.620 5.420 ;
        RECT  7.500 4.090 7.920 5.420 ;
        RECT  8.770 4.100 9.140 5.420 ;
        RECT  10.010 4.100 10.380 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  1.060 3.150 1.540 3.550 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.390 3.580 9.020 3.820 ;
        RECT  8.780 2.400 9.020 3.820 ;
        RECT  2.940 3.520 6.630 3.760 ;
        RECT  2.940 1.490 3.180 3.760 ;
        RECT  8.780 2.400 9.530 2.640 ;
        RECT  9.130 2.280 9.530 2.640 ;
        RECT  2.890 1.490 3.180 1.890 ;
        RECT  5.150 3.010 5.810 3.250 ;
        RECT  5.150 1.570 5.390 3.250 ;
        RECT  5.150 2.360 6.740 2.600 ;
        RECT  6.500 2.200 6.740 2.600 ;
        RECT  4.970 1.570 5.390 1.810 ;
        RECT  1.930 4.080 4.260 4.320 ;
        RECT  3.860 4.020 4.260 4.320 ;
        RECT  1.930 1.490 2.170 4.320 ;
        RECT  3.710 1.490 3.950 3.190 ;
        RECT  3.610 1.490 3.950 1.890 ;
        RECT  0.190 4.080 1.060 4.320 ;
        RECT  0.190 1.490 0.430 4.320 ;
        RECT  0.190 2.790 0.480 3.190 ;
        RECT  0.190 1.490 0.480 1.890 ;
    END
END HA1T

MACRO HA2
    CLASS CORE ;
    FOREIGN HA2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.300 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.890 1.280 3.130 ;
        RECT  0.170 1.290 2.530 1.530 ;
        RECT  0.170 1.290 0.450 3.130 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 0.630 9.130 3.260 ;
        RECT  8.810 2.860 9.130 3.260 ;
        RECT  8.810 1.480 9.130 1.880 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.290 0.720 3.530 2.080 ;
        RECT  1.190 1.840 3.530 2.080 ;
        RECT  3.290 0.720 4.240 1.040 ;
        RECT  3.290 0.800 5.480 1.040 ;
        RECT  5.240 0.620 6.250 0.860 ;
        RECT  1.190 1.840 1.470 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.610 3.410 7.890 4.340 ;
        RECT  3.830 4.000 7.890 4.240 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.490 -0.380 4.890 0.560 ;
        RECT  8.040 -0.380 8.440 0.780 ;
        RECT  0.000 -0.380 9.300 0.380 ;
        RECT  0.160 -0.380 2.720 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.490 4.480 4.890 5.420 ;
        RECT  8.190 4.040 8.510 5.420 ;
        RECT  0.000 4.660 9.300 5.420 ;
        RECT  2.220 4.240 2.620 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.800 3.040 6.200 3.280 ;
        RECT  5.960 1.100 6.200 3.280 ;
        RECT  8.330 2.140 8.610 2.540 ;
        RECT  8.330 1.020 8.570 2.540 ;
        RECT  5.800 1.500 6.200 1.740 ;
        RECT  5.960 1.100 6.670 1.340 ;
        RECT  6.430 1.020 8.570 1.260 ;
        RECT  7.320 2.930 7.720 3.170 ;
        RECT  7.320 1.560 7.560 3.170 ;
        RECT  7.210 2.150 7.560 2.550 ;
        RECT  7.320 1.560 7.720 1.800 ;
        RECT  3.780 3.520 6.920 3.760 ;
        RECT  6.680 1.580 6.920 3.760 ;
        RECT  3.780 1.420 4.020 3.760 ;
        RECT  6.600 3.040 7.000 3.280 ;
        RECT  2.360 2.350 4.020 2.590 ;
        RECT  4.690 2.110 4.930 2.510 ;
        RECT  3.780 2.190 4.930 2.430 ;
        RECT  6.600 1.580 7.000 1.820 ;
        RECT  5.080 3.040 5.480 3.280 ;
        RECT  5.170 1.500 5.410 3.280 ;
        RECT  5.080 1.500 5.480 1.740 ;
        RECT  0.160 3.370 3.160 3.610 ;
        RECT  2.920 3.050 3.160 3.610 ;
    END
END HA2

MACRO HA2P
    CLASS CORE ;
    FOREIGN HA2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.890 2.600 3.130 ;
        RECT  0.750 1.290 5.290 1.530 ;
        RECT  0.790 1.290 1.070 3.130 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 0.630 11.610 3.260 ;
        RECT  11.300 2.860 11.610 3.260 ;
        RECT  11.300 1.480 11.610 1.880 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.770 1.050 6.010 2.080 ;
        RECT  2.630 1.840 6.010 2.080 ;
        RECT  7.810 0.630 8.050 1.290 ;
        RECT  5.770 1.050 8.050 1.290 ;
        RECT  7.810 0.630 8.210 0.870 ;
        RECT  2.630 1.840 2.870 2.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 4.060 6.650 4.340 ;
        RECT  6.370 4.030 6.800 4.270 ;
        RECT  6.370 3.550 6.650 4.340 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  7.060 -0.380 7.460 0.810 ;
        RECT  10.530 -0.380 10.930 0.780 ;
        RECT  11.920 -0.380 12.240 1.160 ;
        RECT  0.000 -0.380 12.400 0.380 ;
        RECT  0.160 -0.380 5.480 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.910 4.240 5.310 5.420 ;
        RECT  7.060 4.480 7.460 5.420 ;
        RECT  10.600 4.120 11.000 5.420 ;
        RECT  11.840 4.120 12.240 5.420 ;
        RECT  0.000 4.660 12.400 5.420 ;
        RECT  3.670 4.240 4.070 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.370 3.070 8.770 3.310 ;
        RECT  8.530 1.050 8.770 3.310 ;
        RECT  10.820 2.140 11.090 2.540 ;
        RECT  10.820 1.050 11.060 2.540 ;
        RECT  8.370 1.530 8.770 1.770 ;
        RECT  8.530 1.050 11.060 1.290 ;
        RECT  9.810 2.930 10.210 3.170 ;
        RECT  9.810 1.560 10.050 3.170 ;
        RECT  9.700 2.150 10.050 2.550 ;
        RECT  9.810 1.560 10.210 1.800 ;
        RECT  7.250 3.630 9.410 3.870 ;
        RECT  9.170 1.530 9.410 3.870 ;
        RECT  7.250 2.110 7.490 3.870 ;
        RECT  9.090 3.070 9.490 3.310 ;
        RECT  6.270 3.070 6.670 3.310 ;
        RECT  6.350 1.530 6.590 3.310 ;
        RECT  5.120 2.350 6.590 2.590 ;
        RECT  7.250 2.110 7.500 2.510 ;
        RECT  6.350 2.190 7.500 2.430 ;
        RECT  9.090 1.530 9.490 1.770 ;
        RECT  6.270 1.530 6.670 1.770 ;
        RECT  7.730 2.990 7.980 3.390 ;
        RECT  7.740 1.530 7.980 3.390 ;
        RECT  7.650 1.530 8.050 1.770 ;
        RECT  1.580 3.370 1.820 4.010 ;
        RECT  0.160 3.370 5.850 3.610 ;
        RECT  5.610 3.050 5.850 3.610 ;
        RECT  4.370 3.050 4.610 3.610 ;
    END
END HA2P

MACRO HA2T
    CLASS CORE ;
    FOREIGN HA2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.890 4.020 3.130 ;
        RECT  0.750 1.550 8.050 1.790 ;
        RECT  0.790 1.550 1.070 3.130 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 0.630 14.710 3.260 ;
        RECT  14.400 2.860 14.710 3.260 ;
        RECT  14.400 1.560 15.880 1.800 ;
        RECT  14.400 2.940 15.880 3.180 ;
        RECT  15.640 1.480 15.880 1.880 ;
        RECT  15.640 2.860 15.880 3.260 ;
        RECT  14.400 1.480 14.710 1.880 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.590 1.050 8.830 2.640 ;
        RECT  3.690 2.400 8.830 2.640 ;
        RECT  10.910 0.630 11.150 1.290 ;
        RECT  8.590 1.050 11.150 1.290 ;
        RECT  10.910 0.630 11.310 0.870 ;
        RECT  3.690 2.350 4.090 2.640 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.500 4.030 9.900 4.340 ;
        RECT  8.850 4.060 9.920 4.340 ;
        RECT  8.850 2.910 9.130 4.340 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  10.160 -0.380 10.560 0.810 ;
        RECT  13.630 -0.380 14.030 0.780 ;
        RECT  15.020 -0.380 15.340 1.160 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  0.160 -0.380 8.660 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.430 4.240 6.830 5.420 ;
        RECT  7.670 4.240 8.070 5.420 ;
        RECT  10.160 4.480 10.560 5.420 ;
        RECT  13.700 4.120 14.100 5.420 ;
        RECT  14.940 4.120 15.340 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  5.010 4.240 5.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.470 3.070 11.870 3.310 ;
        RECT  11.630 1.050 11.870 3.310 ;
        RECT  13.920 2.140 14.190 2.540 ;
        RECT  13.920 1.050 14.160 2.540 ;
        RECT  11.470 1.530 11.870 1.770 ;
        RECT  11.630 1.050 14.160 1.290 ;
        RECT  12.910 2.930 13.310 3.170 ;
        RECT  12.910 1.560 13.150 3.170 ;
        RECT  12.800 2.150 13.150 2.550 ;
        RECT  12.910 1.560 13.310 1.800 ;
        RECT  9.450 3.550 12.510 3.790 ;
        RECT  12.270 1.530 12.510 3.790 ;
        RECT  9.450 1.530 9.690 3.790 ;
        RECT  12.190 3.070 12.590 3.310 ;
        RECT  9.230 2.270 9.690 2.670 ;
        RECT  10.360 2.110 10.600 2.510 ;
        RECT  9.450 2.190 10.600 2.430 ;
        RECT  12.190 1.530 12.590 1.770 ;
        RECT  9.370 1.530 9.770 1.770 ;
        RECT  10.750 3.070 11.150 3.310 ;
        RECT  10.840 1.530 11.080 3.310 ;
        RECT  10.750 1.530 11.150 1.770 ;
        RECT  3.000 3.370 3.240 4.010 ;
        RECT  0.240 3.370 0.480 4.010 ;
        RECT  0.240 3.370 8.610 3.610 ;
        RECT  8.370 3.050 8.610 3.610 ;
        RECT  7.130 3.050 7.370 3.610 ;
        RECT  4.470 3.050 4.710 3.610 ;
    END
END HA2T

MACRO HA3
    CLASS CORE ;
    FOREIGN HA3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.860 1.490 7.100 3.200 ;
        RECT  5.100 2.960 7.100 3.200 ;
        RECT  5.100 2.960 5.500 3.740 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.610 0.730 7.890 3.260 ;
        RECT  7.580 2.860 7.890 3.260 ;
        RECT  7.580 1.480 7.890 1.880 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.810 1.630 1.050 4.370 ;
        RECT  0.720 4.130 1.120 4.370 ;
        RECT  0.740 2.200 1.050 2.600 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.180 0.620 3.420 1.390 ;
        RECT  3.180 1.150 4.290 1.390 ;
        RECT  4.050 1.150 4.290 2.080 ;
        RECT  4.050 1.840 5.390 2.080 ;
        RECT  5.150 1.840 5.390 2.430 ;
        RECT  1.440 0.620 3.420 0.860 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.010 -0.380 5.410 0.560 ;
        RECT  8.200 -0.380 8.540 1.160 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  0.720 -0.380 1.120 0.910 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.690 4.480 6.170 5.420 ;
        RECT  8.120 4.120 8.520 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.240 3.660 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.470 3.990 7.720 4.230 ;
        RECT  7.480 3.640 7.720 4.230 ;
        RECT  4.470 3.650 4.710 4.230 ;
        RECT  3.210 3.650 4.710 3.890 ;
        RECT  7.480 3.640 8.370 3.880 ;
        RECT  8.130 2.140 8.370 3.880 ;
        RECT  3.210 3.040 3.450 3.890 ;
        RECT  2.710 3.040 3.450 3.280 ;
        RECT  2.710 2.880 3.010 3.280 ;
        RECT  2.770 1.580 3.010 3.280 ;
        RECT  6.130 0.930 6.370 2.470 ;
        RECT  4.530 0.930 6.370 1.170 ;
        RECT  4.530 0.620 4.770 1.170 ;
        RECT  3.660 0.620 4.060 0.910 ;
        RECT  3.660 0.620 4.770 0.860 ;
        RECT  1.750 4.180 4.060 4.420 ;
        RECT  3.660 4.130 4.060 4.420 ;
        RECT  1.750 1.580 1.990 4.420 ;
        RECT  3.690 2.560 3.930 3.410 ;
        RECT  3.570 1.660 3.810 2.800 ;
        RECT  3.410 1.660 3.810 1.900 ;
        RECT  2.230 3.540 2.970 3.940 ;
        RECT  2.230 2.400 2.470 3.940 ;
        RECT  0.240 1.150 0.480 3.280 ;
        RECT  2.290 1.100 2.530 2.640 ;
        RECT  0.240 1.150 1.600 1.390 ;
        RECT  1.360 1.100 2.530 1.340 ;
    END
END HA3

MACRO HA3P
    CLASS CORE ;
    FOREIGN HA3P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.250 1.440 8.490 3.200 ;
        RECT  5.100 2.960 8.490 3.200 ;
        RECT  7.940 1.440 8.490 1.840 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 0.630 10.370 3.220 ;
        RECT  10.060 2.820 10.370 3.220 ;
        RECT  10.060 1.240 10.370 1.640 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.760 1.070 4.370 ;
        RECT  0.790 4.130 1.190 4.370 ;
        RECT  0.730 2.200 1.070 2.600 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.160 0.620 3.400 1.390 ;
        RECT  3.160 1.150 4.290 1.390 ;
        RECT  4.050 1.150 4.290 2.320 ;
        RECT  4.050 2.080 4.770 2.320 ;
        RECT  4.530 2.080 4.770 2.640 ;
        RECT  4.530 2.380 5.010 2.640 ;
        RECT  1.440 0.620 3.400 0.860 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.010 -0.380 5.350 0.990 ;
        RECT  6.380 -0.380 6.820 1.150 ;
        RECT  9.380 -0.380 9.750 0.960 ;
        RECT  10.680 -0.380 10.920 0.960 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.720 -0.380 1.120 0.910 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.710 4.480 8.960 5.420 ;
        RECT  9.360 4.120 9.760 5.420 ;
        RECT  10.630 4.040 11.000 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.240 3.660 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.560 3.990 9.120 4.230 ;
        RECT  8.880 3.640 9.120 4.230 ;
        RECT  4.560 3.650 4.800 4.230 ;
        RECT  3.210 3.650 4.800 3.890 ;
        RECT  8.880 3.640 9.820 3.880 ;
        RECT  9.580 2.140 9.820 3.880 ;
        RECT  3.210 3.040 3.450 3.890 ;
        RECT  2.710 3.040 3.450 3.280 ;
        RECT  2.710 2.880 3.010 3.280 ;
        RECT  2.770 1.580 3.010 3.280 ;
        RECT  9.580 2.140 9.850 2.540 ;
        RECT  5.730 1.390 7.460 1.630 ;
        RECT  7.220 0.910 7.460 1.630 ;
        RECT  5.730 0.750 5.970 1.630 ;
        RECT  7.220 0.910 8.980 1.150 ;
        RECT  7.580 2.280 7.820 2.680 ;
        RECT  5.250 2.320 7.820 2.560 ;
        RECT  5.250 1.550 5.490 2.560 ;
        RECT  4.530 1.550 5.490 1.790 ;
        RECT  4.530 0.670 4.770 1.790 ;
        RECT  3.640 0.670 4.770 0.910 ;
        RECT  1.750 4.180 4.060 4.420 ;
        RECT  3.660 4.130 4.060 4.420 ;
        RECT  1.750 1.580 1.990 4.420 ;
        RECT  3.690 2.560 3.930 3.410 ;
        RECT  3.410 2.560 3.930 2.800 ;
        RECT  3.410 1.660 3.650 2.800 ;
        RECT  3.410 1.660 3.810 1.900 ;
        RECT  2.230 3.540 2.970 3.940 ;
        RECT  2.230 2.400 2.470 3.940 ;
        RECT  0.190 2.880 0.480 3.280 ;
        RECT  0.190 1.280 0.430 3.280 ;
        RECT  2.290 1.100 2.530 2.640 ;
        RECT  0.190 1.280 0.480 1.890 ;
        RECT  0.190 1.280 1.510 1.520 ;
        RECT  1.270 1.100 2.530 1.340 ;
    END
END HA3P

MACRO HA3T
    CLASS CORE ;
    FOREIGN HA3T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.640 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 1.820 9.750 3.240 ;
        RECT  5.200 3.000 10.460 3.240 ;
        RECT  10.240 1.630 10.640 2.100 ;
        RECT  8.800 1.820 10.640 2.100 ;
        RECT  8.800 1.630 9.200 2.100 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 0.630 12.230 3.350 ;
        RECT  11.920 2.950 12.230 3.350 ;
        RECT  13.160 1.480 13.470 1.880 ;
        RECT  11.950 2.400 13.470 2.640 ;
        RECT  13.190 0.630 13.470 3.350 ;
        RECT  13.160 2.950 13.470 3.350 ;
        RECT  11.920 1.480 12.230 1.880 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.760 1.070 4.370 ;
        RECT  0.790 4.130 1.190 4.370 ;
        RECT  0.730 2.200 1.070 2.600 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.160 0.620 3.400 1.390 ;
        RECT  3.160 1.150 4.290 1.390 ;
        RECT  4.050 1.150 4.290 2.300 ;
        RECT  4.050 2.060 4.770 2.300 ;
        RECT  4.530 2.060 4.770 2.640 ;
        RECT  4.530 2.400 4.930 2.640 ;
        RECT  1.440 0.620 3.400 0.860 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.010 -0.380 5.350 0.990 ;
        RECT  5.640 -0.380 6.070 0.990 ;
        RECT  7.230 -0.380 7.630 0.910 ;
        RECT  11.240 -0.380 11.610 1.160 ;
        RECT  12.540 -0.380 12.780 1.170 ;
        RECT  0.000 -0.380 13.640 0.380 ;
        RECT  0.720 -0.380 1.120 0.910 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.400 4.190 4.800 5.420 ;
        RECT  5.990 4.190 6.390 5.420 ;
        RECT  7.600 4.190 8.000 5.420 ;
        RECT  9.240 4.190 9.640 5.420 ;
        RECT  10.880 4.190 11.280 5.420 ;
        RECT  12.490 4.140 12.860 5.420 ;
        RECT  0.000 4.660 13.640 5.420 ;
        RECT  0.240 3.660 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.210 3.650 11.680 3.890 ;
        RECT  11.440 2.140 11.680 3.890 ;
        RECT  3.210 3.040 3.450 3.890 ;
        RECT  2.710 3.040 3.450 3.280 ;
        RECT  2.710 2.880 3.010 3.280 ;
        RECT  2.770 1.580 3.010 3.280 ;
        RECT  11.440 2.140 11.710 2.540 ;
        RECT  6.440 1.230 8.450 1.470 ;
        RECT  8.210 0.670 8.450 1.470 ;
        RECT  8.210 0.670 9.920 0.910 ;
        RECT  5.170 2.340 8.610 2.580 ;
        RECT  5.170 1.550 5.410 2.580 ;
        RECT  4.530 1.550 5.410 1.790 ;
        RECT  4.530 0.620 4.770 1.790 ;
        RECT  3.640 0.620 4.040 0.910 ;
        RECT  3.640 0.620 4.770 0.860 ;
        RECT  1.750 4.180 4.060 4.420 ;
        RECT  3.660 4.130 4.060 4.420 ;
        RECT  1.750 1.580 1.990 4.420 ;
        RECT  3.690 2.560 3.930 3.410 ;
        RECT  3.410 2.560 3.930 2.800 ;
        RECT  3.410 1.660 3.650 2.800 ;
        RECT  3.410 1.660 3.810 1.900 ;
        RECT  2.230 3.540 2.970 3.940 ;
        RECT  2.230 2.400 2.470 3.940 ;
        RECT  0.190 2.880 0.480 3.280 ;
        RECT  0.190 1.280 0.430 3.280 ;
        RECT  2.290 1.100 2.530 2.640 ;
        RECT  0.190 1.280 0.480 1.890 ;
        RECT  0.190 1.280 1.510 1.520 ;
        RECT  1.270 1.100 2.530 1.340 ;
    END
END HA3T

MACRO INV1
    CLASS CORE ;
    FOREIGN INV1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.860 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.490 0.480 1.890 ;
        RECT  0.170 2.840 0.480 3.240 ;
        RECT  0.170 1.180 0.450 3.300 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.070 2.840 ;
        RECT  0.690 2.220 1.070 2.620 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.860 0.380 ;
        RECT  0.930 -0.380 1.170 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 1.860 5.420 ;
        RECT  0.680 3.910 1.080 5.420 ;
        END
    END VCC
END INV1

MACRO INV12
    CLASS CORE ;
    FOREIGN INV12 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.210 1.280 6.660 3.760 ;
        RECT  0.790 3.080 6.660 3.760 ;
        RECT  0.790 1.280 6.660 1.910 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.070 2.200 2.930 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.460 -0.380 1.860 1.040 ;
        RECT  2.760 -0.380 3.160 1.010 ;
        RECT  4.210 -0.380 4.610 1.040 ;
        RECT  5.540 -0.380 5.940 1.040 ;
        RECT  6.840 -0.380 7.240 1.040 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.160 -0.380 0.560 1.010 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.460 4.110 1.860 5.420 ;
        RECT  2.760 4.140 3.160 5.420 ;
        RECT  4.260 4.140 4.660 5.420 ;
        RECT  5.580 4.100 5.980 5.420 ;
        RECT  6.880 4.110 7.280 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.160 4.110 0.560 5.420 ;
        END
    END VCC
END INV12

MACRO INV12CK
    CLASS CORE ;
    FOREIGN INV12CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.300 0.840 2.740 4.420 ;
        RECT  3.740 0.840 4.180 4.420 ;
        RECT  5.180 0.840 5.620 4.420 ;
        RECT  6.620 0.840 7.060 4.420 ;
        RECT  0.860 1.680 8.500 3.360 ;
        RECT  8.060 0.840 8.500 4.420 ;
        RECT  0.860 0.790 1.300 4.420 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.760 0.480 2.160 ;
        RECT  0.170 1.630 0.450 2.270 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 1.130 ;
        RECT  3.040 -0.380 3.440 1.130 ;
        RECT  4.480 -0.380 4.880 1.130 ;
        RECT  5.920 -0.380 6.320 1.130 ;
        RECT  7.360 -0.380 7.760 1.130 ;
        RECT  8.870 -0.380 9.270 1.130 ;
        RECT  0.000 -0.380 9.920 0.380 ;
        RECT  0.160 -0.380 0.560 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 3.910 2.000 5.420 ;
        RECT  3.040 3.910 3.440 5.420 ;
        RECT  4.480 3.910 4.880 5.420 ;
        RECT  5.920 3.910 6.320 5.420 ;
        RECT  7.360 3.910 7.760 5.420 ;
        RECT  8.870 3.910 9.270 5.420 ;
        RECT  0.000 4.660 9.920 5.420 ;
        RECT  0.160 3.910 0.560 5.420 ;
        END
    END VCC
END INV12CK

MACRO INV1CK
    CLASS CORE ;
    FOREIGN INV1CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.860 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 0.870 0.480 1.270 ;
        RECT  0.170 2.950 0.480 4.010 ;
        RECT  0.170 0.790 0.450 4.330 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.070 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.860 0.380 ;
        RECT  0.880 -0.380 1.280 1.130 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 1.860 5.420 ;
        RECT  1.160 3.910 1.560 5.420 ;
        END
    END VCC
END INV1CK

MACRO INV1S
    CLASS CORE ;
    FOREIGN INV1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.240 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.290 1.070 3.190 ;
        RECT  0.760 2.790 1.070 3.190 ;
        RECT  0.430 1.290 1.070 1.770 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.150 2.120 0.480 2.800 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.240 0.380 ;
        RECT  0.440 -0.380 0.840 1.030 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 1.240 5.420 ;
        RECT  0.160 3.540 0.560 5.420 ;
        END
    END VCC
END INV1S

MACRO INV2
    CLASS CORE ;
    FOREIGN INV2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.860 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.180 1.070 3.300 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.550 2.740 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 -0.380 1.700 0.560 ;
        RECT  0.000 -0.380 1.860 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 4.480 1.700 5.420 ;
        RECT  0.000 4.660 1.860 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
END INV2

MACRO INV2CK
    CLASS CORE ;
    FOREIGN INV2CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 0.860 1.200 1.260 ;
        RECT  0.790 2.950 1.200 4.010 ;
        RECT  0.790 0.790 1.070 4.330 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.760 0.480 2.160 ;
        RECT  0.170 1.630 0.450 2.270 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 1.130 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.160 -0.380 0.480 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 3.910 2.000 5.420 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.160 3.910 0.480 5.420 ;
        END
    END VCC
END INV2CK

MACRO INV3
    CLASS CORE ;
    FOREIGN INV3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.260 1.690 3.220 ;
        RECT  0.750 1.260 2.320 1.890 ;
        RECT  0.750 2.940 2.320 3.220 ;
        RECT  0.750 2.880 0.990 3.280 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.220 0.480 2.620 ;
        RECT  0.170 2.180 0.450 2.790 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 -0.380 1.700 0.560 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.340 4.480 1.740 5.420 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
END INV3

MACRO INV3CK
    CLASS CORE ;
    FOREIGN INV3CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.100 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.860 2.230 2.740 2.810 ;
        RECT  2.300 0.840 2.740 3.940 ;
        RECT  0.860 0.860 1.300 4.420 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.760 0.480 2.160 ;
        RECT  0.170 1.630 0.450 2.270 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 1.130 ;
        RECT  0.000 -0.380 3.100 0.380 ;
        RECT  0.160 -0.380 0.480 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 3.910 2.000 5.420 ;
        RECT  0.000 4.660 3.100 5.420 ;
        RECT  0.160 3.910 0.480 5.420 ;
        END
    END VCC
END INV3CK

MACRO INV4
    CLASS CORE ;
    FOREIGN INV4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.100 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.000 1.520 2.390 3.240 ;
        RECT  0.690 2.920 2.390 3.240 ;
        RECT  0.760 1.280 2.320 1.910 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.760 2.650 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.230 -0.380 1.630 0.560 ;
        RECT  2.540 -0.380 2.940 1.160 ;
        RECT  0.000 -0.380 3.100 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.230 4.480 1.630 5.420 ;
        RECT  2.540 4.180 2.940 5.420 ;
        RECT  0.000 4.660 3.100 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
END INV4

MACRO INV4CK
    CLASS CORE ;
    FOREIGN INV4CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 0.860 1.200 1.260 ;
        RECT  0.790 3.520 1.200 4.420 ;
        RECT  0.790 2.230 2.740 2.810 ;
        RECT  2.300 0.840 2.740 3.940 ;
        RECT  0.790 0.790 1.070 4.420 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.760 0.480 2.160 ;
        RECT  0.170 1.630 0.450 2.270 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 1.130 ;
        RECT  3.040 -0.380 3.440 1.130 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.160 -0.380 0.480 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 3.910 2.000 5.420 ;
        RECT  3.040 3.910 3.440 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.160 3.910 0.480 5.420 ;
        END
    END VCC
END INV4CK

MACRO INV6
    CLASS CORE ;
    FOREIGN INV6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.780 1.260 4.250 3.220 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.870 0.480 2.270 ;
        RECT  0.170 1.740 0.450 2.380 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.550 -0.380 1.950 1.000 ;
        RECT  2.280 -0.380 2.680 0.390 ;
        RECT  3.010 -0.380 3.410 1.000 ;
        RECT  4.400 -0.380 4.800 1.000 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.160 -0.380 0.560 1.000 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.390 3.870 1.790 5.420 ;
        RECT  2.280 4.650 2.680 5.420 ;
        RECT  3.170 3.870 3.570 5.420 ;
        RECT  4.410 3.870 4.800 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.160 3.870 0.550 5.420 ;
        END
    END VCC
END INV6

MACRO INV6CK
    CLASS CORE ;
    FOREIGN INV6CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 0.860 1.200 1.260 ;
        RECT  0.790 3.520 1.200 4.420 ;
        RECT  2.300 0.840 2.740 4.420 ;
        RECT  0.790 2.100 4.180 2.940 ;
        RECT  3.740 0.840 4.180 4.420 ;
        RECT  0.790 0.790 1.070 4.420 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.760 0.480 2.160 ;
        RECT  0.170 1.630 0.450 2.270 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 1.130 ;
        RECT  3.040 -0.380 3.440 1.130 ;
        RECT  4.550 -0.380 4.950 1.130 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.160 -0.380 0.480 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 3.910 2.000 5.420 ;
        RECT  3.040 3.910 3.440 5.420 ;
        RECT  4.550 3.910 4.950 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.160 3.910 0.480 5.420 ;
        END
    END VCC
END INV6CK

MACRO INV8
    CLASS CORE ;
    FOREIGN INV8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.190 1.360 5.410 3.740 ;
        RECT  0.770 3.040 5.410 3.740 ;
        RECT  0.850 1.360 5.410 1.880 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 2.240 2.940 2.800 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.530 -0.380 1.930 1.060 ;
        RECT  2.910 -0.380 3.310 0.560 ;
        RECT  4.270 -0.380 4.670 1.060 ;
        RECT  5.640 -0.380 6.040 1.010 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.140 -0.380 0.580 0.960 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.460 4.020 1.860 5.420 ;
        RECT  2.760 4.020 3.160 5.420 ;
        RECT  4.240 4.000 4.660 5.420 ;
        RECT  5.640 4.020 6.040 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.160 4.020 0.560 5.420 ;
        END
    END VCC
END INV8

MACRO INV8CK
    CLASS CORE ;
    FOREIGN INV8CK 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.300 0.840 2.740 4.420 ;
        RECT  3.740 0.840 4.180 4.420 ;
        RECT  0.860 2.100 5.620 2.940 ;
        RECT  5.180 0.840 5.620 4.420 ;
        RECT  0.860 0.790 1.300 4.420 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.760 0.480 2.160 ;
        RECT  0.170 1.630 0.450 2.270 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 1.130 ;
        RECT  3.040 -0.380 3.440 1.130 ;
        RECT  4.480 -0.380 4.880 1.130 ;
        RECT  5.990 -0.380 6.390 1.130 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  0.160 -0.380 0.480 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 3.910 2.000 5.420 ;
        RECT  3.040 3.910 3.440 5.420 ;
        RECT  4.480 3.910 4.880 5.420 ;
        RECT  5.990 3.910 6.390 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  0.160 3.910 0.480 5.420 ;
        END
    END VCC
END INV8CK

MACRO INVT1
    CLASS CORE ;
    FOREIGN INVT1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.100 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.620 2.980 2.930 3.380 ;
        RECT  2.650 0.620 2.930 3.860 ;
        RECT  2.620 1.220 2.930 1.620 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.370 2.440 1.690 2.840 ;
        RECT  1.410 2.200 1.690 2.840 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.180 1.070 2.380 ;
        RECT  0.790 1.260 2.310 1.500 ;
        RECT  2.030 1.180 2.310 2.160 ;
        RECT  0.730 1.830 1.070 2.230 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.380 1.540 0.860 ;
        RECT  0.000 -0.380 3.100 0.380 ;
        RECT  0.300 -0.380 0.700 0.390 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.200 4.180 1.600 5.420 ;
        RECT  0.000 4.660 3.100 5.420 ;
        RECT  0.300 4.650 0.700 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.190 3.540 2.290 3.780 ;
        RECT  2.050 2.440 2.290 3.780 ;
        RECT  0.190 2.980 0.480 3.780 ;
        RECT  0.190 1.220 0.430 3.780 ;
        RECT  0.190 1.220 0.480 1.620 ;
    END
END INVT1

MACRO INVT2
    CLASS CORE ;
    FOREIGN INVT2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 0.620 3.550 3.260 ;
        RECT  2.600 2.980 3.550 3.260 ;
        RECT  2.450 0.620 3.550 0.900 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.260 1.820 2.660 ;
        RECT  1.410 2.940 2.310 3.220 ;
        RECT  2.030 2.940 2.310 4.340 ;
        RECT  3.150 3.510 3.430 4.340 ;
        RECT  2.030 4.060 3.430 4.340 ;
        RECT  3.800 2.330 4.170 2.730 ;
        RECT  3.890 2.330 4.170 3.790 ;
        RECT  3.150 3.510 4.170 3.790 ;
        RECT  1.410 2.260 1.690 3.220 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.470 1.090 1.580 1.330 ;
        RECT  1.340 1.240 2.930 1.480 ;
        RECT  2.650 1.240 2.930 2.180 ;
        RECT  0.470 0.880 0.870 1.330 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.790 -0.380 4.130 1.890 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  1.260 -0.380 1.660 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.690 4.120 4.090 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  1.180 3.850 1.500 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.500 2.820 0.790 3.220 ;
        RECT  0.500 1.570 0.740 3.220 ;
        RECT  2.170 2.460 2.770 2.700 ;
        RECT  2.170 1.770 2.410 2.700 ;
        RECT  0.500 1.770 2.410 2.010 ;
        RECT  0.470 1.570 0.870 1.810 ;
    END
END INVT2

MACRO INVT4
    CLASS CORE ;
    FOREIGN INVT4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.760 1.260 7.890 1.540 ;
        RECT  7.610 1.230 7.890 3.220 ;
        RECT  5.750 2.940 7.890 3.220 ;
        RECT  5.750 2.960 7.950 3.200 ;
        RECT  7.560 1.230 7.960 1.470 ;
        RECT  5.930 1.230 6.330 1.540 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.230 2.240 3.570 2.800 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.490 2.140 ;
        RECT  0.170 1.640 0.450 2.280 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.380 2.940 0.730 ;
        RECT  5.310 -0.380 5.710 0.800 ;
        RECT  6.860 -0.380 7.260 0.800 ;
        RECT  8.110 -0.380 8.510 0.800 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  0.980 -0.380 1.380 0.610 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.720 3.720 4.120 5.420 ;
        RECT  5.040 4.100 5.440 5.420 ;
        RECT  6.630 4.100 7.030 5.420 ;
        RECT  8.060 4.100 8.460 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  1.180 4.180 1.420 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.430 2.990 4.770 3.390 ;
        RECT  4.530 1.840 4.770 3.390 ;
        RECT  4.530 2.400 6.690 2.640 ;
        RECT  6.290 2.320 6.690 2.640 ;
        RECT  4.350 1.100 4.590 2.080 ;
        RECT  3.880 1.100 4.590 1.340 ;
        RECT  2.160 2.880 2.430 3.280 ;
        RECT  1.750 2.880 2.430 3.200 ;
        RECT  1.750 0.970 1.990 3.200 ;
        RECT  5.150 1.780 6.000 2.080 ;
        RECT  5.150 1.280 5.390 2.080 ;
        RECT  4.830 1.280 5.390 1.520 ;
        RECT  4.830 0.620 5.070 1.520 ;
        RECT  1.750 0.970 3.530 1.210 ;
        RECT  3.290 0.620 3.530 1.210 ;
        RECT  3.290 0.620 5.070 0.860 ;
        RECT  2.670 3.060 3.130 3.460 ;
        RECT  2.670 1.660 2.910 3.460 ;
        RECT  2.230 2.050 2.910 2.640 ;
        RECT  3.860 1.660 4.100 2.070 ;
        RECT  2.670 1.660 4.100 1.960 ;
        RECT  3.130 1.570 3.530 1.960 ;
        RECT  3.040 4.080 3.440 4.420 ;
        RECT  2.050 4.080 3.440 4.320 ;
        RECT  2.050 3.520 2.290 4.320 ;
        RECT  0.160 3.790 0.970 4.030 ;
        RECT  0.730 3.520 0.970 4.030 ;
        RECT  0.730 3.520 2.290 3.760 ;
        RECT  0.160 2.980 0.560 3.310 ;
        RECT  0.160 2.980 1.290 3.220 ;
        RECT  1.050 1.050 1.290 3.220 ;
        RECT  0.160 1.050 1.290 1.290 ;
    END
END INVT4

MACRO JKFN
    CLASS CORE ;
    FOREIGN JKFN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.760 2.310 3.100 ;
        RECT  1.850 2.120 2.310 2.520 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.210 0.690 2.610 ;
        RECT  0.170 1.920 0.450 3.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.120 4.790 2.840 ;
        RECT  4.390 2.230 4.790 2.630 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 1.480 14.710 3.200 ;
        RECT  14.400 2.800 14.710 3.200 ;
        RECT  14.400 1.480 14.710 1.880 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.080 0.620 13.360 1.540 ;
        RECT  13.190 1.260 13.470 3.190 ;
        RECT  12.960 2.790 13.470 3.190 ;
        RECT  12.960 0.620 13.360 1.020 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.410 -0.380 1.810 0.560 ;
        RECT  2.590 -0.380 2.990 0.560 ;
        RECT  4.800 -0.380 5.940 0.560 ;
        RECT  8.690 -0.380 9.090 0.840 ;
        RECT  11.580 -0.380 11.980 0.560 ;
        RECT  13.600 -0.380 14.000 0.940 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  0.670 -0.380 1.070 0.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 4.480 2.070 5.420 ;
        RECT  3.360 4.480 3.760 5.420 ;
        RECT  4.710 4.480 5.110 5.420 ;
        RECT  8.850 4.200 9.250 5.420 ;
        RECT  11.780 4.480 12.180 5.420 ;
        RECT  13.600 4.260 14.000 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  12.450 3.780 14.140 4.020 ;
        RECT  13.900 2.160 14.140 4.020 ;
        RECT  12.450 1.490 12.690 4.020 ;
        RECT  11.400 2.980 12.690 3.220 ;
        RECT  11.400 2.820 11.640 3.220 ;
        RECT  7.290 3.700 7.690 3.940 ;
        RECT  7.290 0.620 7.530 3.940 ;
        RECT  10.440 0.800 10.680 3.200 ;
        RECT  11.970 0.800 12.210 2.430 ;
        RECT  8.210 1.080 10.680 1.320 ;
        RECT  10.440 0.800 11.060 1.090 ;
        RECT  8.210 0.620 8.450 1.320 ;
        RECT  10.440 0.800 12.210 1.040 ;
        RECT  7.290 0.620 8.450 0.860 ;
        RECT  6.810 4.180 8.170 4.420 ;
        RECT  7.930 3.620 8.170 4.420 ;
        RECT  6.360 3.700 7.050 4.240 ;
        RECT  1.110 4.000 7.050 4.240 ;
        RECT  7.930 3.620 10.310 3.860 ;
        RECT  10.070 3.600 11.270 3.840 ;
        RECT  6.810 0.620 7.050 4.420 ;
        RECT  10.920 1.490 11.160 3.840 ;
        RECT  10.920 1.490 11.270 1.890 ;
        RECT  6.300 0.620 7.050 0.860 ;
        RECT  8.680 2.880 10.200 3.120 ;
        RECT  9.960 1.580 10.200 3.120 ;
        RECT  8.680 2.260 8.920 3.120 ;
        RECT  9.640 1.580 10.200 1.820 ;
        RECT  7.770 1.500 8.010 3.200 ;
        RECT  9.160 2.340 9.680 2.580 ;
        RECT  9.160 1.730 9.400 2.580 ;
        RECT  7.770 1.730 9.400 1.970 ;
        RECT  2.750 3.030 3.150 3.270 ;
        RECT  6.330 1.100 6.570 3.200 ;
        RECT  2.830 1.570 3.070 3.270 ;
        RECT  2.830 1.570 4.290 1.810 ;
        RECT  4.050 0.800 4.290 1.810 ;
        RECT  5.740 1.100 6.570 1.340 ;
        RECT  5.740 0.800 5.980 1.340 ;
        RECT  4.050 0.800 5.980 1.040 ;
        RECT  5.500 3.520 5.910 3.760 ;
        RECT  5.670 1.580 5.910 3.760 ;
        RECT  5.670 2.460 6.010 2.860 ;
        RECT  5.530 1.580 5.930 1.820 ;
        RECT  4.080 3.520 5.240 3.760 ;
        RECT  5.000 3.060 5.240 3.760 ;
        RECT  5.040 2.900 5.330 3.300 ;
        RECT  5.040 1.580 5.280 3.300 ;
        RECT  4.750 1.580 5.280 1.820 ;
        RECT  2.000 1.280 2.400 1.520 ;
        RECT  2.160 0.850 2.400 1.520 ;
        RECT  2.160 0.850 3.810 1.090 ;
        RECT  0.960 3.520 3.650 3.760 ;
        RECT  3.410 2.360 3.650 3.760 ;
        RECT  0.960 1.440 1.200 3.760 ;
        RECT  3.330 2.360 3.730 2.600 ;
        RECT  0.160 1.440 1.200 1.680 ;
    END
END JKFN

MACRO JKFRBN
    CLASS CORE ;
    FOREIGN JKFRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.740 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 3.300 12.850 3.940 ;
        RECT  12.460 3.300 12.850 3.700 ;
        END
    END RB
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.990 2.500 ;
        RECT  1.410 1.740 1.690 2.740 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.050 0.490 2.450 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.080 2.380 4.790 2.660 ;
        RECT  4.510 2.380 4.790 3.240 ;
        RECT  4.080 1.460 4.360 2.660 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 1.480 16.570 3.280 ;
        RECT  16.260 2.880 16.570 3.280 ;
        RECT  16.260 1.480 16.570 1.880 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.050 1.480 15.330 3.370 ;
        RECT  14.820 2.970 15.330 3.370 ;
        RECT  14.820 1.480 15.330 1.880 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.480 -0.380 6.060 0.560 ;
        RECT  12.560 -0.380 13.500 0.570 ;
        RECT  15.460 -0.380 15.860 1.030 ;
        RECT  0.000 -0.380 16.740 0.380 ;
        RECT  1.320 -0.380 2.720 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.480 4.480 1.880 5.420 ;
        RECT  3.300 4.480 3.700 5.420 ;
        RECT  4.900 4.480 5.300 5.420 ;
        RECT  9.930 4.480 10.330 5.420 ;
        RECT  13.380 4.180 14.320 5.420 ;
        RECT  15.460 4.260 15.860 5.420 ;
        RECT  0.000 4.660 16.740 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.780 3.700 15.890 3.940 ;
        RECT  15.650 2.120 15.890 3.940 ;
        RECT  14.340 0.780 14.580 3.940 ;
        RECT  13.780 2.940 14.020 3.940 ;
        RECT  13.130 2.940 14.020 3.180 ;
        RECT  15.650 2.120 15.970 2.520 ;
        RECT  14.020 0.780 14.580 1.020 ;
        RECT  7.550 3.700 7.950 3.940 ;
        RECT  7.550 0.620 7.790 3.940 ;
        RECT  13.860 1.290 14.100 2.580 ;
        RECT  13.010 1.290 14.100 1.530 ;
        RECT  7.550 1.100 10.170 1.340 ;
        RECT  9.930 0.620 10.170 1.340 ;
        RECT  13.010 0.810 13.250 1.530 ;
        RECT  12.040 0.810 13.250 1.050 ;
        RECT  9.930 0.620 12.280 0.860 ;
        RECT  10.570 4.180 12.860 4.420 ;
        RECT  7.070 4.180 8.430 4.420 ;
        RECT  8.190 3.700 8.430 4.420 ;
        RECT  9.900 4.000 10.810 4.240 ;
        RECT  3.290 4.000 6.730 4.240 ;
        RECT  6.490 3.620 6.730 4.240 ;
        RECT  11.980 2.680 12.220 4.420 ;
        RECT  7.070 0.620 7.310 4.420 ;
        RECT  9.900 3.700 10.140 4.240 ;
        RECT  3.290 3.680 3.530 4.240 ;
        RECT  8.190 3.700 10.140 3.940 ;
        RECT  0.990 3.680 3.530 3.920 ;
        RECT  6.490 3.620 7.310 3.860 ;
        RECT  12.220 1.640 12.460 2.920 ;
        RECT  6.650 0.620 7.310 0.860 ;
        RECT  10.380 3.520 11.740 3.760 ;
        RECT  11.500 2.200 11.740 3.760 ;
        RECT  10.380 3.180 10.620 3.760 ;
        RECT  8.830 3.180 10.620 3.420 ;
        RECT  11.560 1.100 11.800 2.440 ;
        RECT  8.790 1.580 9.190 1.860 ;
        RECT  8.790 1.580 10.650 1.820 ;
        RECT  10.410 1.100 10.650 1.820 ;
        RECT  10.410 1.100 11.800 1.340 ;
        RECT  10.860 3.040 11.260 3.280 ;
        RECT  10.940 1.720 11.180 3.280 ;
        RECT  9.210 2.160 9.670 2.400 ;
        RECT  10.890 1.720 11.180 2.300 ;
        RECT  9.430 2.060 11.180 2.300 ;
        RECT  10.890 1.720 11.320 1.960 ;
        RECT  8.030 1.620 8.270 3.300 ;
        RECT  8.030 2.640 10.290 2.880 ;
        RECT  9.890 2.540 10.290 2.880 ;
        RECT  8.030 1.620 8.430 1.860 ;
        RECT  8.750 0.620 9.690 0.860 ;
        RECT  8.670 4.180 9.660 4.420 ;
        RECT  6.590 1.100 6.830 3.300 ;
        RECT  2.820 2.920 3.840 3.160 ;
        RECT  3.600 0.800 3.840 3.160 ;
        RECT  5.760 1.100 6.830 1.340 ;
        RECT  5.760 0.800 6.000 1.340 ;
        RECT  3.600 0.800 6.000 1.040 ;
        RECT  3.760 0.740 4.160 1.040 ;
        RECT  5.690 3.480 6.090 3.720 ;
        RECT  5.850 1.580 6.090 3.720 ;
        RECT  5.850 2.500 6.200 2.900 ;
        RECT  5.690 1.580 6.090 1.820 ;
        RECT  4.260 3.480 5.310 3.720 ;
        RECT  5.070 1.540 5.310 3.720 ;
        RECT  5.070 2.720 5.490 3.120 ;
        RECT  5.010 1.540 5.310 1.940 ;
        RECT  2.180 1.260 3.360 1.500 ;
        RECT  3.120 0.660 3.360 1.500 ;
        RECT  0.810 3.000 2.470 3.240 ;
        RECT  2.230 2.440 2.470 3.240 ;
        RECT  0.810 2.840 1.080 3.240 ;
        RECT  0.810 1.260 1.050 3.240 ;
        RECT  2.230 2.440 3.330 2.680 ;
        RECT  3.090 2.280 3.330 2.680 ;
        RECT  0.160 1.260 1.050 1.500 ;
    END
END JKFRBN

MACRO JKFRBP
    CLASS CORE ;
    FOREIGN JKFRBP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.980 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 3.300 12.850 3.940 ;
        RECT  12.460 3.300 12.850 3.700 ;
        END
    END RB
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.990 2.500 ;
        RECT  1.410 1.740 1.690 2.740 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.050 0.490 2.450 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.080 2.380 4.790 2.660 ;
        RECT  4.510 2.380 4.790 3.240 ;
        RECT  4.080 1.460 4.360 2.660 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.530 1.300 17.810 3.220 ;
        RECT  16.700 2.940 17.810 3.220 ;
        RECT  16.700 1.300 17.810 1.580 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.990 1.460 15.660 1.700 ;
        RECT  14.990 2.960 15.660 3.200 ;
        RECT  14.990 1.460 15.390 3.200 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.480 -0.380 6.060 0.560 ;
        RECT  12.690 -0.380 13.630 0.570 ;
        RECT  14.540 -0.380 14.940 0.840 ;
        RECT  15.980 -0.380 16.380 0.840 ;
        RECT  17.420 -0.380 17.820 0.840 ;
        RECT  0.000 -0.380 17.980 0.380 ;
        RECT  1.320 -0.380 2.720 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.480 4.480 1.880 5.420 ;
        RECT  3.300 4.480 3.700 5.420 ;
        RECT  4.900 4.480 5.300 5.420 ;
        RECT  9.930 4.480 10.330 5.420 ;
        RECT  13.380 4.180 13.780 5.420 ;
        RECT  14.540 4.260 14.940 5.420 ;
        RECT  15.980 4.260 16.380 5.420 ;
        RECT  17.420 4.260 17.820 5.420 ;
        RECT  0.000 4.660 17.980 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.780 3.700 16.410 3.940 ;
        RECT  16.170 2.160 16.410 3.940 ;
        RECT  14.340 1.360 14.580 3.940 ;
        RECT  13.780 2.820 14.020 3.940 ;
        RECT  13.130 2.820 14.020 3.060 ;
        RECT  16.170 2.160 16.490 2.560 ;
        RECT  14.020 1.360 14.580 1.600 ;
        RECT  7.550 3.700 7.950 3.940 ;
        RECT  7.550 0.620 7.790 3.940 ;
        RECT  13.860 2.180 14.100 2.580 ;
        RECT  13.010 2.180 14.100 2.420 ;
        RECT  13.010 0.810 13.250 2.420 ;
        RECT  7.550 1.100 10.170 1.340 ;
        RECT  9.930 0.620 10.170 1.340 ;
        RECT  12.040 0.810 13.250 1.050 ;
        RECT  9.930 0.620 12.280 0.860 ;
        RECT  10.570 4.180 12.860 4.420 ;
        RECT  7.070 4.180 8.430 4.420 ;
        RECT  8.190 3.700 8.430 4.420 ;
        RECT  9.900 4.000 10.810 4.240 ;
        RECT  3.290 4.000 6.730 4.240 ;
        RECT  6.490 3.620 6.730 4.240 ;
        RECT  11.980 2.680 12.220 4.420 ;
        RECT  7.070 0.620 7.310 4.420 ;
        RECT  9.900 3.700 10.140 4.240 ;
        RECT  3.290 3.680 3.530 4.240 ;
        RECT  8.190 3.700 10.140 3.940 ;
        RECT  0.990 3.680 3.530 3.920 ;
        RECT  6.490 3.620 7.310 3.860 ;
        RECT  12.220 1.640 12.460 2.920 ;
        RECT  6.650 0.620 7.310 0.860 ;
        RECT  10.380 3.520 11.740 3.760 ;
        RECT  11.500 2.200 11.740 3.760 ;
        RECT  10.380 3.180 10.620 3.760 ;
        RECT  8.830 3.180 10.620 3.420 ;
        RECT  11.560 1.100 11.800 2.440 ;
        RECT  8.790 1.580 9.190 1.860 ;
        RECT  8.790 1.580 10.650 1.820 ;
        RECT  10.410 1.100 10.650 1.820 ;
        RECT  10.410 1.100 11.800 1.340 ;
        RECT  10.860 3.040 11.260 3.280 ;
        RECT  10.940 1.720 11.180 3.280 ;
        RECT  9.210 2.160 9.670 2.400 ;
        RECT  10.890 1.720 11.180 2.300 ;
        RECT  9.430 2.060 11.180 2.300 ;
        RECT  10.890 1.720 11.320 1.960 ;
        RECT  8.030 1.620 8.270 3.300 ;
        RECT  8.030 2.640 10.290 2.880 ;
        RECT  9.890 2.540 10.290 2.880 ;
        RECT  8.030 1.620 8.430 1.860 ;
        RECT  8.750 0.620 9.690 0.860 ;
        RECT  8.670 4.180 9.660 4.420 ;
        RECT  6.590 1.100 6.830 3.300 ;
        RECT  2.820 2.920 3.840 3.160 ;
        RECT  3.600 0.800 3.840 3.160 ;
        RECT  5.760 1.100 6.830 1.340 ;
        RECT  5.760 0.800 6.000 1.340 ;
        RECT  3.600 0.800 6.000 1.040 ;
        RECT  3.760 0.740 4.160 1.040 ;
        RECT  5.690 3.480 6.090 3.720 ;
        RECT  5.850 1.580 6.090 3.720 ;
        RECT  5.850 2.500 6.200 2.900 ;
        RECT  5.690 1.580 6.090 1.820 ;
        RECT  4.260 3.480 5.310 3.720 ;
        RECT  5.070 1.540 5.310 3.720 ;
        RECT  5.070 2.720 5.490 3.120 ;
        RECT  5.010 1.540 5.310 1.940 ;
        RECT  2.180 1.260 3.360 1.500 ;
        RECT  3.120 0.660 3.360 1.500 ;
        RECT  0.810 3.000 2.470 3.240 ;
        RECT  2.230 2.440 2.470 3.240 ;
        RECT  0.810 2.840 1.080 3.240 ;
        RECT  0.810 1.260 1.050 3.240 ;
        RECT  2.230 2.440 3.330 2.680 ;
        RECT  3.090 2.280 3.330 2.680 ;
        RECT  0.160 1.260 1.050 1.500 ;
    END
END JKFRBP

MACRO JKZN
    CLASS CORE ;
    FOREIGN JKZN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.980 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.760 2.310 3.100 ;
        RECT  1.880 2.120 2.310 2.520 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.400 0.690 2.800 ;
        RECT  0.170 1.920 0.450 3.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.230 8.750 2.630 ;
        RECT  8.230 2.230 8.510 2.800 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.270 6.790 2.670 ;
        RECT  6.370 2.120 6.650 2.800 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.530 1.480 17.810 3.200 ;
        RECT  17.500 2.800 17.810 3.200 ;
        RECT  17.500 1.480 17.810 1.880 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.180 0.620 16.460 1.540 ;
        RECT  16.290 1.260 16.570 3.200 ;
        RECT  16.060 2.800 16.570 3.200 ;
        RECT  16.060 0.620 16.460 1.020 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.610 2.120 7.890 2.800 ;
        RECT  7.340 2.120 7.890 2.570 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.410 -0.380 1.810 0.560 ;
        RECT  2.590 -0.380 2.990 0.560 ;
        RECT  3.330 -0.380 4.250 0.460 ;
        RECT  6.460 -0.380 6.860 0.560 ;
        RECT  8.950 -0.380 9.350 0.560 ;
        RECT  15.130 -0.380 15.530 0.560 ;
        RECT  16.700 -0.380 17.100 0.940 ;
        RECT  0.000 -0.380 17.980 0.380 ;
        RECT  0.670 -0.380 1.070 0.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 4.480 2.070 5.420 ;
        RECT  3.550 4.480 3.950 5.420 ;
        RECT  6.700 4.480 7.100 5.420 ;
        RECT  8.870 4.480 9.270 5.420 ;
        RECT  12.670 4.480 13.070 5.420 ;
        RECT  14.500 4.480 14.900 5.420 ;
        RECT  16.700 4.260 17.100 5.420 ;
        RECT  0.000 4.660 17.980 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  15.470 3.850 15.870 4.090 ;
        RECT  17.010 2.160 17.250 4.020 ;
        RECT  15.550 3.780 17.250 4.020 ;
        RECT  15.550 1.480 15.790 4.090 ;
        RECT  14.710 2.560 15.790 2.800 ;
        RECT  14.710 2.400 14.950 2.800 ;
        RECT  15.240 0.800 15.640 1.100 ;
        RECT  14.650 0.800 15.640 1.040 ;
        RECT  11.420 0.620 14.890 0.860 ;
        RECT  11.420 3.520 11.820 3.920 ;
        RECT  11.420 3.520 15.200 3.760 ;
        RECT  14.960 3.080 15.200 3.760 ;
        RECT  9.890 4.160 11.180 4.400 ;
        RECT  10.940 0.620 11.180 4.400 ;
        RECT  8.200 4.000 10.130 4.240 ;
        RECT  1.110 4.000 4.920 4.240 ;
        RECT  4.680 3.520 4.920 4.240 ;
        RECT  10.540 3.680 11.180 4.400 ;
        RECT  8.200 3.520 8.440 4.240 ;
        RECT  4.680 3.520 8.440 3.760 ;
        RECT  14.170 3.040 14.600 3.280 ;
        RECT  14.170 1.100 14.410 3.280 ;
        RECT  10.940 1.100 14.410 1.340 ;
        RECT  10.430 0.620 11.180 0.860 ;
        RECT  12.410 3.040 13.920 3.280 ;
        RECT  13.680 1.580 13.920 3.280 ;
        RECT  12.410 2.260 12.650 3.280 ;
        RECT  13.370 1.580 13.920 1.820 ;
        RECT  11.500 1.580 11.740 3.200 ;
        RECT  12.890 2.260 13.330 2.660 ;
        RECT  12.890 1.580 13.130 2.660 ;
        RECT  11.420 1.580 13.130 1.820 ;
        RECT  10.460 1.100 10.700 3.200 ;
        RECT  5.490 2.560 5.890 2.800 ;
        RECT  5.570 1.280 5.810 2.800 ;
        RECT  4.930 1.280 7.960 1.520 ;
        RECT  7.720 1.100 10.700 1.340 ;
        RECT  7.560 1.260 10.700 1.340 ;
        RECT  4.930 0.700 5.170 1.520 ;
        RECT  4.770 0.700 5.170 0.940 ;
        RECT  9.660 3.040 10.060 3.280 ;
        RECT  9.800 1.580 10.040 3.280 ;
        RECT  9.800 2.260 10.220 2.660 ;
        RECT  9.660 1.580 10.060 1.820 ;
        RECT  8.280 3.040 9.420 3.280 ;
        RECT  9.180 1.680 9.420 3.280 ;
        RECT  9.180 2.420 9.520 2.820 ;
        RECT  8.280 1.680 9.420 1.920 ;
        RECT  8.280 1.580 8.680 1.920 ;
        RECT  5.820 0.800 7.340 1.040 ;
        RECT  7.100 0.620 8.620 0.860 ;
        RECT  5.820 0.620 6.220 1.040 ;
        RECT  4.700 3.040 7.890 3.280 ;
        RECT  7.490 4.000 7.890 4.420 ;
        RECT  5.840 4.000 7.890 4.240 ;
        RECT  2.750 3.040 3.150 3.280 ;
        RECT  2.830 2.000 3.070 3.280 ;
        RECT  2.830 2.000 5.240 2.240 ;
        RECT  5.000 1.840 5.240 2.240 ;
        RECT  4.110 1.360 4.350 2.240 ;
        RECT  0.960 3.520 3.650 3.760 ;
        RECT  3.410 2.480 3.650 3.760 ;
        RECT  0.960 1.440 1.200 3.760 ;
        RECT  3.330 2.480 3.730 2.720 ;
        RECT  0.160 1.440 1.200 1.680 ;
        RECT  2.000 1.280 3.710 1.520 ;
    END
END JKZN

MACRO JKZRBN
    CLASS CORE ;
    FOREIGN JKZRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.080 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.230 2.080 16.630 2.320 ;
        RECT  16.290 1.180 16.570 2.320 ;
        END
    END RB
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.740 2.310 2.760 ;
        RECT  1.880 2.300 2.310 2.700 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.610 0.490 3.010 ;
        RECT  0.170 2.570 0.450 3.350 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.310 8.510 3.150 ;
        RECT  8.230 2.750 8.720 3.150 ;
        RECT  8.120 1.310 8.510 1.710 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 1.640 7.270 2.840 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  20.630 0.630 20.910 3.200 ;
        RECT  20.520 2.960 20.920 3.200 ;
        RECT  20.600 1.490 20.910 1.890 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  19.120 2.880 19.670 3.280 ;
        RECT  19.390 1.570 19.670 3.860 ;
        RECT  18.940 1.570 19.670 1.810 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.960 6.150 2.360 ;
        RECT  5.750 1.860 6.030 3.100 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 -0.380 1.780 1.810 ;
        RECT  4.310 -0.380 4.550 1.700 ;
        RECT  6.730 -0.380 7.130 0.840 ;
        RECT  15.190 -0.380 16.760 0.840 ;
        RECT  16.520 -0.380 16.760 0.920 ;
        RECT  19.730 -0.380 20.130 0.850 ;
        RECT  0.000 -0.380 21.080 0.380 ;
        RECT  0.840 -0.380 1.780 0.570 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.550 4.200 1.950 5.420 ;
        RECT  3.300 4.480 3.700 5.420 ;
        RECT  4.920 4.480 5.320 5.420 ;
        RECT  8.460 4.400 8.860 5.420 ;
        RECT  16.010 4.480 16.410 5.420 ;
        RECT  18.030 4.480 18.430 5.420 ;
        RECT  19.800 4.260 20.200 5.420 ;
        RECT  0.000 4.660 21.080 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.640 4.180 15.770 4.420 ;
        RECT  15.530 3.520 15.770 4.420 ;
        RECT  11.190 0.700 11.430 4.420 ;
        RECT  15.530 3.520 18.210 3.760 ;
        RECT  17.970 2.020 18.210 3.760 ;
        RECT  20.030 2.120 20.370 2.520 ;
        RECT  17.000 2.020 18.210 2.260 ;
        RECT  20.030 1.090 20.270 2.520 ;
        RECT  17.000 0.620 17.240 2.260 ;
        RECT  19.120 1.090 20.270 1.330 ;
        RECT  19.120 0.620 19.360 1.330 ;
        RECT  10.850 0.700 11.430 0.940 ;
        RECT  17.000 0.620 19.360 0.860 ;
        RECT  16.970 4.000 18.690 4.240 ;
        RECT  18.450 1.540 18.690 4.240 ;
        RECT  18.450 2.220 18.830 2.620 ;
        RECT  17.480 1.540 18.690 1.780 ;
        RECT  11.670 3.700 12.070 3.940 ;
        RECT  11.750 0.620 11.990 3.940 ;
        RECT  15.750 2.560 17.490 2.800 ;
        RECT  17.090 2.500 17.490 2.800 ;
        RECT  15.750 1.090 15.990 2.800 ;
        RECT  14.710 1.090 15.990 1.330 ;
        RECT  11.750 0.620 12.050 1.190 ;
        RECT  14.710 0.620 14.950 1.330 ;
        RECT  11.750 0.620 14.950 0.860 ;
        RECT  13.930 3.220 14.650 3.460 ;
        RECT  13.930 3.220 15.390 3.320 ;
        RECT  15.070 3.040 17.390 3.280 ;
        RECT  14.410 3.080 17.390 3.280 ;
        RECT  15.070 1.700 15.310 3.320 ;
        RECT  14.370 1.700 14.610 2.100 ;
        RECT  14.370 1.700 15.310 1.940 ;
        RECT  15.110 1.660 15.510 1.900 ;
        RECT  13.090 3.700 15.290 3.940 ;
        RECT  13.160 2.740 13.400 3.940 ;
        RECT  13.160 2.740 14.090 2.980 ;
        RECT  13.850 1.100 14.090 2.980 ;
        RECT  13.540 1.100 14.090 1.340 ;
        RECT  12.230 2.980 12.630 3.220 ;
        RECT  12.230 1.680 12.470 3.220 ;
        RECT  13.210 2.220 13.610 2.500 ;
        RECT  12.230 2.220 13.610 2.460 ;
        RECT  12.230 1.680 12.630 1.920 ;
        RECT  10.710 1.260 10.950 3.300 ;
        RECT  6.390 1.140 6.630 3.100 ;
        RECT  5.510 1.380 6.630 1.620 ;
        RECT  10.370 1.260 10.950 1.500 ;
        RECT  7.380 0.620 7.620 1.380 ;
        RECT  6.390 1.140 7.620 1.380 ;
        RECT  10.370 0.620 10.610 1.500 ;
        RECT  7.380 0.620 10.610 0.860 ;
        RECT  9.990 1.840 10.230 4.170 ;
        RECT  9.990 3.560 10.850 3.800 ;
        RECT  9.890 1.540 10.130 2.080 ;
        RECT  7.750 3.770 8.180 4.170 ;
        RECT  7.750 3.770 9.410 4.010 ;
        RECT  9.170 2.120 9.410 4.010 ;
        RECT  9.160 2.810 9.410 3.210 ;
        RECT  9.020 2.120 9.410 2.520 ;
        RECT  4.130 3.340 7.530 3.580 ;
        RECT  7.130 3.100 7.530 3.580 ;
        RECT  5.770 4.180 6.700 4.420 ;
        RECT  4.280 4.000 6.010 4.240 ;
        RECT  2.820 3.180 3.220 3.420 ;
        RECT  2.870 2.860 3.220 3.420 ;
        RECT  2.870 2.860 5.470 3.100 ;
        RECT  5.230 1.960 5.470 3.100 ;
        RECT  2.870 1.490 3.110 3.420 ;
        RECT  3.590 2.370 4.870 2.610 ;
        RECT  3.590 1.300 3.830 2.610 ;
        RECT  0.810 3.720 3.450 3.960 ;
        RECT  0.810 3.560 1.080 3.960 ;
        RECT  0.810 1.570 1.050 3.960 ;
        RECT  0.160 1.570 1.050 1.810 ;
    END
END JKZRBN

MACRO JKZRBP
    CLASS CORE ;
    FOREIGN JKZRBP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.320 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.210 2.080 16.610 2.320 ;
        RECT  16.290 1.180 16.570 2.320 ;
        END
    END RB
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.740 2.310 2.760 ;
        RECT  1.880 2.300 2.310 2.700 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.610 0.490 3.010 ;
        RECT  0.170 2.570 0.450 3.350 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.310 8.510 3.150 ;
        RECT  8.230 2.750 8.720 3.150 ;
        RECT  8.120 1.310 8.510 1.710 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 1.640 7.270 2.840 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  21.870 1.530 22.150 3.220 ;
        RECT  21.040 2.940 22.150 3.220 ;
        RECT  21.040 1.530 22.150 1.810 ;
        END
    END QB
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  20.010 1.570 20.290 3.200 ;
        RECT  19.600 2.960 20.290 3.200 ;
        RECT  19.600 1.570 20.290 1.810 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.960 6.150 2.360 ;
        RECT  5.750 1.860 6.030 3.100 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 -0.380 1.780 1.810 ;
        RECT  4.310 -0.380 4.550 1.700 ;
        RECT  6.730 -0.380 7.130 0.840 ;
        RECT  15.170 -0.380 16.740 0.840 ;
        RECT  16.500 -0.380 16.740 0.920 ;
        RECT  18.760 -0.380 19.160 0.580 ;
        RECT  20.320 -0.380 20.720 0.950 ;
        RECT  21.760 -0.380 22.160 0.950 ;
        RECT  0.000 -0.380 22.320 0.380 ;
        RECT  0.840 -0.380 1.780 0.570 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.550 4.200 1.950 5.420 ;
        RECT  3.300 4.480 3.700 5.420 ;
        RECT  4.920 4.480 5.320 5.420 ;
        RECT  8.460 4.400 8.860 5.420 ;
        RECT  15.990 4.480 16.390 5.420 ;
        RECT  18.010 4.480 18.950 5.420 ;
        RECT  20.320 4.260 20.720 5.420 ;
        RECT  21.760 4.260 22.160 5.420 ;
        RECT  0.000 4.660 22.320 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.640 4.180 15.750 4.420 ;
        RECT  15.510 3.520 15.750 4.420 ;
        RECT  11.190 0.700 11.430 4.420 ;
        RECT  15.510 3.520 18.190 3.760 ;
        RECT  17.950 2.020 18.190 3.760 ;
        RECT  19.010 3.440 20.800 3.680 ;
        RECT  20.560 2.240 20.800 3.680 ;
        RECT  19.010 1.060 19.250 3.680 ;
        RECT  20.560 2.240 20.960 2.480 ;
        RECT  16.980 2.020 18.190 2.260 ;
        RECT  16.980 1.060 17.220 2.260 ;
        RECT  16.980 1.060 19.250 1.300 ;
        RECT  10.850 0.700 11.430 0.940 ;
        RECT  16.950 4.000 18.670 4.240 ;
        RECT  18.430 1.540 18.670 4.240 ;
        RECT  17.460 1.540 18.670 1.780 ;
        RECT  11.670 3.700 12.070 3.940 ;
        RECT  11.750 0.620 11.990 3.940 ;
        RECT  15.730 2.560 17.470 2.800 ;
        RECT  17.070 2.500 17.470 2.800 ;
        RECT  15.730 1.090 15.970 2.800 ;
        RECT  14.690 1.090 15.970 1.330 ;
        RECT  11.750 0.620 12.050 1.190 ;
        RECT  14.690 0.620 14.930 1.330 ;
        RECT  11.750 0.620 14.930 0.860 ;
        RECT  13.910 3.220 14.630 3.460 ;
        RECT  13.910 3.220 15.370 3.320 ;
        RECT  15.050 3.040 17.370 3.280 ;
        RECT  14.390 3.080 17.370 3.280 ;
        RECT  15.050 1.700 15.290 3.320 ;
        RECT  14.350 1.700 14.590 2.100 ;
        RECT  14.350 1.700 15.290 1.940 ;
        RECT  15.090 1.660 15.490 1.900 ;
        RECT  13.090 3.700 15.270 3.940 ;
        RECT  13.160 2.740 13.400 3.940 ;
        RECT  13.160 2.740 14.090 2.980 ;
        RECT  13.850 1.100 14.090 2.980 ;
        RECT  13.540 1.100 14.090 1.340 ;
        RECT  12.230 2.980 12.630 3.220 ;
        RECT  12.230 1.680 12.470 3.220 ;
        RECT  13.210 2.220 13.610 2.500 ;
        RECT  12.230 2.220 13.610 2.460 ;
        RECT  12.230 1.680 12.630 1.920 ;
        RECT  10.710 1.260 10.950 3.300 ;
        RECT  6.390 1.140 6.630 3.100 ;
        RECT  5.510 1.380 6.630 1.620 ;
        RECT  10.370 1.260 10.950 1.500 ;
        RECT  7.380 0.620 7.620 1.380 ;
        RECT  6.390 1.140 7.620 1.380 ;
        RECT  10.370 0.620 10.610 1.500 ;
        RECT  7.380 0.620 10.610 0.860 ;
        RECT  9.990 1.840 10.230 4.170 ;
        RECT  9.990 3.560 10.850 3.800 ;
        RECT  9.890 1.540 10.130 2.080 ;
        RECT  7.750 3.770 8.180 4.170 ;
        RECT  7.750 3.770 9.410 4.010 ;
        RECT  9.170 2.120 9.410 4.010 ;
        RECT  9.160 2.810 9.410 3.210 ;
        RECT  9.020 2.120 9.410 2.520 ;
        RECT  4.130 3.340 7.530 3.580 ;
        RECT  7.130 3.100 7.530 3.580 ;
        RECT  5.770 4.180 6.700 4.420 ;
        RECT  4.280 4.000 6.010 4.240 ;
        RECT  2.820 3.180 3.220 3.420 ;
        RECT  2.870 2.860 3.220 3.420 ;
        RECT  2.870 2.860 5.470 3.100 ;
        RECT  5.230 1.960 5.470 3.100 ;
        RECT  2.870 1.490 3.110 3.420 ;
        RECT  3.590 2.370 4.870 2.610 ;
        RECT  3.590 1.300 3.830 2.610 ;
        RECT  0.810 3.720 3.450 3.960 ;
        RECT  0.810 3.560 1.080 3.960 ;
        RECT  0.810 1.570 1.050 3.960 ;
        RECT  0.160 1.570 1.050 1.810 ;
    END
END JKZRBP

MACRO MAO222
    CLASS CORE ;
    FOREIGN MAO222 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.330 4.790 3.280 ;
        RECT  4.340 2.880 4.790 3.280 ;
        RECT  4.340 1.330 4.790 1.730 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.730 1.690 2.180 ;
        RECT  1.190 1.730 2.950 1.970 ;
        RECT  1.190 1.730 1.690 2.130 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.210 2.310 2.740 ;
        RECT  1.950 2.210 2.310 2.610 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.540 2.650 ;
        RECT  0.170 3.020 3.550 3.260 ;
        RECT  3.270 2.250 3.550 3.300 ;
        RECT  0.170 2.250 0.450 3.300 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.270 -0.380 3.670 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.980 -0.380 1.380 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.370 4.480 3.770 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.320 3.540 4.030 3.780 ;
        RECT  3.790 1.130 4.030 3.780 ;
        RECT  3.790 2.130 4.270 2.530 ;
        RECT  2.320 1.130 4.030 1.370 ;
        RECT  0.160 1.130 2.000 1.370 ;
        RECT  0.160 3.540 2.000 3.780 ;
    END
END MAO222

MACRO MAO222P
    CLASS CORE ;
    FOREIGN MAO222P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.400 1.260 5.410 1.540 ;
        RECT  5.130 1.260 5.410 3.220 ;
        RECT  4.500 2.940 5.410 3.220 ;
        RECT  4.500 2.790 4.740 3.220 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.730 1.690 2.180 ;
        RECT  1.290 1.730 3.090 1.970 ;
        RECT  2.690 1.730 3.090 2.030 ;
        RECT  1.290 1.730 1.690 2.030 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.210 2.430 2.740 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.070 3.300 ;
        RECT  0.790 3.020 3.550 3.260 ;
        RECT  3.270 2.250 3.550 3.300 ;
        RECT  3.270 2.250 3.730 2.650 ;
        RECT  0.710 2.250 1.070 2.650 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 -0.380 4.180 0.780 ;
        RECT  5.020 -0.380 5.420 0.780 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.950 -0.380 1.350 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 4.210 4.180 5.420 ;
        RECT  5.020 4.210 5.420 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.460 3.540 4.260 3.780 ;
        RECT  4.020 1.760 4.260 3.780 ;
        RECT  4.020 2.130 4.460 2.530 ;
        RECT  3.600 1.760 4.260 2.000 ;
        RECT  3.600 1.190 3.840 2.000 ;
        RECT  2.460 1.190 3.840 1.430 ;
        RECT  0.160 1.190 2.140 1.430 ;
        RECT  0.160 3.540 2.140 3.780 ;
    END
END MAO222P

MACRO MAO222S
    CLASS CORE ;
    FOREIGN MAO222S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.330 4.790 3.280 ;
        RECT  4.480 2.880 4.790 3.280 ;
        RECT  4.480 1.330 4.790 1.730 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.580 3.090 2.820 ;
        RECT  0.790 2.300 1.070 2.820 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.600 2.310 2.340 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.880 0.510 3.300 ;
        RECT  3.450 2.340 3.690 3.300 ;
        RECT  0.170 3.060 3.690 3.300 ;
        RECT  0.170 2.570 0.450 3.300 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 -0.380 4.010 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.430 -0.380 1.830 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 4.480 4.010 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  1.060 4.480 1.460 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.930 3.540 4.590 4.040 ;
        RECT  2.460 3.540 4.590 3.780 ;
        RECT  3.930 1.410 4.170 4.040 ;
        RECT  2.560 1.410 4.170 1.650 ;
        RECT  0.160 3.540 2.140 3.780 ;
        RECT  1.510 1.330 1.750 1.730 ;
        RECT  0.160 1.410 1.750 1.650 ;
    END
END MAO222S

MACRO MAO222T
    CLASS CORE ;
    FOREIGN MAO222T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 1.300 5.410 3.180 ;
        RECT  4.380 1.300 6.040 1.540 ;
        RECT  4.450 2.940 6.040 3.180 ;
        RECT  4.450 2.940 4.690 3.340 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.730 1.690 2.180 ;
        RECT  1.290 1.730 3.090 1.970 ;
        RECT  2.690 1.730 3.090 2.030 ;
        RECT  1.290 1.730 1.690 2.030 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.210 2.430 2.740 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.070 3.300 ;
        RECT  3.270 2.250 3.550 3.260 ;
        RECT  0.790 3.020 3.550 3.260 ;
        RECT  3.270 2.250 3.730 2.650 ;
        RECT  0.710 2.250 1.070 2.650 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.710 -0.380 4.110 0.880 ;
        RECT  5.020 -0.380 5.420 0.880 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.950 -0.380 1.350 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.760 4.210 4.160 5.420 ;
        RECT  5.020 4.210 5.420 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.460 3.540 4.210 3.780 ;
        RECT  3.970 1.770 4.210 3.780 ;
        RECT  3.970 2.130 4.440 2.530 ;
        RECT  3.600 1.770 4.210 2.010 ;
        RECT  3.600 1.190 3.840 2.010 ;
        RECT  2.460 1.190 3.840 1.430 ;
        RECT  0.160 1.190 2.140 1.430 ;
        RECT  0.160 3.540 2.140 3.780 ;
    END
END MAO222T

MACRO MAOI1
    CLASS CORE ;
    FOREIGN MAOI1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 1.200 4.790 1.600 ;
        RECT  4.480 2.790 4.790 3.190 ;
        RECT  4.510 1.180 4.790 3.300 ;
        RECT  2.330 1.220 4.790 1.500 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 2.300 1.740 2.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.300 0.580 2.760 ;
        RECT  0.170 1.740 0.450 2.760 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.250 3.700 2.740 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 2.250 2.930 2.740 ;
        RECT  2.650 1.740 2.930 2.740 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.610 -0.380 2.010 0.560 ;
        RECT  3.580 -0.380 3.980 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.960 4.260 3.360 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.260 4.480 0.660 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.820 2.980 4.240 3.220 ;
        RECT  4.000 2.250 4.240 3.220 ;
        RECT  0.820 1.490 1.060 3.220 ;
        RECT  4.000 2.250 4.270 2.650 ;
        RECT  0.820 1.490 1.170 1.890 ;
        RECT  2.240 3.520 4.100 3.760 ;
    END
END MAOI1

MACRO MAOI1H
    CLASS CORE ;
    FOREIGN MAOI1H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.440 0.710 5.680 1.630 ;
        RECT  6.240 2.790 6.650 3.190 ;
        RECT  6.370 1.390 6.650 3.300 ;
        RECT  5.440 1.390 7.280 1.630 ;
        RECT  4.000 0.710 5.680 0.950 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 2.190 1.740 2.630 ;
        RECT  1.410 2.190 1.690 3.060 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.580 2.650 ;
        RECT  0.170 1.740 0.450 2.650 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.250 3.550 3.060 ;
        RECT  3.130 2.250 3.550 2.650 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.250 4.810 2.650 ;
        RECT  4.510 2.250 4.790 3.060 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 1.250 ;
        RECT  3.130 -0.380 3.530 0.950 ;
        RECT  6.160 -0.380 6.560 1.150 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.160 -0.380 0.560 1.250 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.280 4.260 3.680 5.420 ;
        RECT  4.720 4.260 5.120 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.560 3.780 7.280 4.020 ;
        RECT  0.820 3.300 6.000 3.540 ;
        RECT  5.760 2.250 6.000 3.540 ;
        RECT  0.820 1.490 1.060 3.540 ;
        RECT  5.760 2.250 6.030 2.650 ;
        RECT  0.820 1.490 1.200 1.890 ;
        RECT  2.320 1.190 5.120 1.430 ;
    END
END MAOI1H

MACRO MAOI1HP
    CLASS CORE ;
    FOREIGN MAOI1HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.580 0.710 9.980 1.150 ;
        RECT  9.740 0.710 9.980 1.810 ;
        RECT  11.950 1.570 12.230 3.940 ;
        RECT  10.300 3.700 12.230 3.940 ;
        RECT  9.740 1.570 12.860 1.810 ;
        RECT  6.700 0.710 9.980 0.950 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.250 2.310 2.900 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.070 3.160 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.250 4.810 2.650 ;
        RECT  4.510 1.830 4.790 2.650 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.830 8.510 2.650 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 1.250 ;
        RECT  3.040 -0.380 3.440 1.250 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  5.920 -0.380 6.320 0.950 ;
        RECT  10.300 -0.380 10.700 1.150 ;
        RECT  11.740 -0.380 12.140 1.150 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  0.160 -0.380 0.560 1.250 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.540 3.930 4.940 5.420 ;
        RECT  5.980 4.260 6.380 5.420 ;
        RECT  7.420 4.180 7.820 5.420 ;
        RECT  8.860 4.180 9.260 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.580 4.180 12.860 4.420 ;
        RECT  9.580 3.450 9.860 4.420 ;
        RECT  3.820 3.450 9.860 3.690 ;
        RECT  2.320 3.140 2.790 3.380 ;
        RECT  2.550 1.570 2.790 3.380 ;
        RECT  9.260 2.330 9.500 3.210 ;
        RECT  2.550 2.970 9.500 3.210 ;
        RECT  9.260 2.330 10.970 2.570 ;
        RECT  0.880 1.570 2.790 1.810 ;
        RECT  3.760 1.190 9.260 1.430 ;
        RECT  0.160 3.780 3.440 4.020 ;
    END
END MAOI1HP

MACRO MAOI1HT
    CLASS CORE ;
    FOREIGN MAOI1HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.600 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.720 0.710 14.120 1.150 ;
        RECT  13.880 0.710 14.120 1.810 ;
        RECT  16.290 1.570 16.570 3.940 ;
        RECT  14.440 3.700 17.720 3.940 ;
        RECT  13.880 1.570 18.440 1.810 ;
        RECT  9.400 0.710 14.120 0.950 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.250 4.170 2.900 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 1.690 3.160 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.250 6.670 2.650 ;
        RECT  6.370 1.830 6.650 2.650 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 1.830 12.230 2.650 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.560 -0.380 2.000 1.250 ;
        RECT  3.040 -0.380 3.440 1.250 ;
        RECT  4.480 -0.380 4.880 1.250 ;
        RECT  5.920 -0.380 6.320 0.950 ;
        RECT  7.360 -0.380 7.760 0.950 ;
        RECT  8.800 -0.380 9.140 1.790 ;
        RECT  14.440 -0.380 14.840 1.150 ;
        RECT  15.880 -0.380 16.280 1.150 ;
        RECT  17.320 -0.380 17.720 1.150 ;
        RECT  0.000 -0.380 18.600 0.380 ;
        RECT  0.160 -0.380 0.560 1.250 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  5.800 3.930 6.200 5.420 ;
        RECT  7.240 3.930 7.640 5.420 ;
        RECT  8.680 4.260 9.080 5.420 ;
        RECT  10.120 4.180 10.520 5.420 ;
        RECT  11.560 4.180 11.960 5.420 ;
        RECT  13.000 3.910 13.400 5.420 ;
        RECT  0.000 4.660 18.600 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.720 4.180 18.440 4.420 ;
        RECT  13.720 3.430 14.000 4.420 ;
        RECT  5.160 3.430 5.400 3.990 ;
        RECT  5.160 3.430 14.120 3.670 ;
        RECT  2.920 3.300 4.720 3.540 ;
        RECT  4.480 2.950 4.720 3.540 ;
        RECT  2.920 1.570 3.160 3.540 ;
        RECT  4.480 2.950 13.640 3.190 ;
        RECT  13.400 2.330 13.640 3.190 ;
        RECT  13.400 2.330 15.110 2.570 ;
        RECT  0.880 1.570 4.160 1.810 ;
        RECT  8.160 2.030 10.440 2.270 ;
        RECT  10.200 1.190 10.440 2.270 ;
        RECT  8.160 1.190 8.400 2.270 ;
        RECT  10.200 1.190 13.400 1.430 ;
        RECT  5.200 1.190 8.400 1.430 ;
        RECT  0.880 3.780 4.160 4.020 ;
    END
END MAOI1HT

MACRO MAOI1S
    CLASS CORE ;
    FOREIGN MAOI1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 1.170 4.790 1.570 ;
        RECT  4.510 0.620 4.790 3.860 ;
        RECT  4.480 3.460 4.790 3.860 ;
        RECT  2.330 1.210 4.790 1.490 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 2.300 1.740 2.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.300 0.580 2.760 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.250 3.700 2.740 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.740 2.930 2.200 ;
        RECT  2.500 1.740 2.930 2.140 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.610 -0.380 2.010 0.560 ;
        RECT  3.580 -0.380 3.980 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.960 4.480 3.360 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.260 4.480 0.660 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.820 2.980 4.240 3.220 ;
        RECT  4.000 2.250 4.240 3.220 ;
        RECT  0.820 1.490 1.060 3.220 ;
        RECT  4.000 2.250 4.270 2.650 ;
        RECT  0.820 1.490 1.070 1.890 ;
        RECT  2.240 3.480 4.100 3.720 ;
    END
END MAOI1S

MACRO MOAI1
    CLASS CORE ;
    FOREIGN MOAI1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.180 3.550 3.260 ;
        RECT  2.530 2.980 3.550 3.260 ;
        RECT  3.180 1.180 3.550 1.580 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.250 1.740 1.690 2.180 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.600 3.420 1.090 3.870 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.130 4.170 2.740 ;
        RECT  3.850 2.130 4.170 2.530 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.490 1.740 2.930 2.240 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  1.440 -0.380 1.840 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.980 3.820 2.300 5.420 ;
        RECT  3.780 4.080 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.160 4.160 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.220 0.620 4.130 0.860 ;
        RECT  1.020 2.420 1.420 3.030 ;
        RECT  0.240 2.420 2.250 2.660 ;
        RECT  2.010 2.090 2.250 2.660 ;
        RECT  0.240 1.300 0.480 2.660 ;
    END
END MOAI1

MACRO MOAI1H
    CLASS CORE ;
    FOREIGN MOAI1H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.320 3.300 6.030 3.540 ;
        RECT  4.720 1.190 6.560 1.430 ;
        RECT  5.750 1.190 6.030 3.540 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 2.170 1.690 2.570 ;
        RECT  1.410 1.660 1.690 2.570 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.620 2.170 1.070 2.570 ;
        RECT  0.790 1.660 1.070 2.570 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.250 6.650 2.900 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.250 4.810 2.650 ;
        RECT  4.510 2.250 4.790 2.900 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.040 -0.380 3.440 1.330 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  1.600 -0.380 2.000 1.130 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 3.910 2.000 5.420 ;
        RECT  3.040 3.780 3.440 5.420 ;
        RECT  6.160 4.260 6.560 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.160 3.910 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.320 1.570 4.400 1.810 ;
        RECT  4.160 0.710 4.400 1.810 ;
        RECT  4.160 0.710 7.280 0.950 ;
        RECT  4.000 3.780 7.280 4.020 ;
        RECT  0.880 2.820 1.280 3.300 ;
        RECT  0.140 2.820 2.410 3.060 ;
        RECT  2.170 2.250 2.410 3.060 ;
        RECT  0.140 1.300 0.380 3.060 ;
        RECT  0.140 1.300 0.480 1.700 ;
    END
END MOAI1H

MACRO MOAI1HP
    CLASS CORE ;
    FOREIGN MOAI1HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.760 3.300 9.750 3.540 ;
        RECT  7.420 1.190 12.140 1.430 ;
        RECT  9.470 1.190 9.750 3.540 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.070 3.160 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.250 2.310 3.160 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.250 11.610 2.900 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.250 8.530 2.650 ;
        RECT  8.230 2.250 8.510 2.900 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.540 -0.380 4.940 1.130 ;
        RECT  5.980 -0.380 6.380 0.950 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  5.920 3.780 6.320 5.420 ;
        RECT  10.300 4.260 10.700 5.420 ;
        RECT  11.740 4.260 12.140 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.820 1.570 7.100 1.810 ;
        RECT  6.860 0.710 7.100 1.810 ;
        RECT  6.860 0.710 12.860 0.950 ;
        RECT  6.700 3.780 12.860 4.020 ;
        RECT  0.880 3.780 3.520 4.020 ;
        RECT  3.280 2.820 3.520 4.020 ;
        RECT  2.550 1.570 2.790 4.020 ;
        RECT  3.280 2.820 3.850 3.060 ;
        RECT  3.610 2.250 3.850 3.060 ;
        RECT  2.320 1.570 2.790 1.810 ;
        RECT  0.160 1.570 1.840 1.810 ;
        RECT  1.600 1.090 1.840 1.810 ;
        RECT  1.600 1.090 3.440 1.330 ;
    END
END MOAI1HP

MACRO MOAI1HT
    CLASS CORE ;
    FOREIGN MOAI1HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.600 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.190 13.470 3.300 ;
        RECT  5.200 3.060 13.470 3.300 ;
        RECT  13.190 1.570 17.720 1.810 ;
        RECT  10.120 1.190 13.470 1.430 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.250 3.550 3.160 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 1.690 3.160 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 2.250 16.570 2.900 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.150 11.630 2.550 ;
        RECT  11.330 2.150 11.610 2.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.480 -0.380 4.880 1.230 ;
        RECT  5.920 -0.380 6.320 1.230 ;
        RECT  7.360 -0.380 7.760 1.130 ;
        RECT  8.800 -0.380 9.200 0.950 ;
        RECT  0.000 -0.380 18.600 0.380 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 3.910 4.880 5.420 ;
        RECT  5.920 3.910 6.320 5.420 ;
        RECT  7.360 4.260 7.760 5.420 ;
        RECT  8.800 4.260 9.200 5.420 ;
        RECT  14.440 3.910 14.840 5.420 ;
        RECT  15.880 4.260 16.280 5.420 ;
        RECT  17.320 4.260 17.720 5.420 ;
        RECT  0.000 4.660 18.600 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.200 1.570 9.800 1.810 ;
        RECT  9.560 0.710 9.800 1.810 ;
        RECT  13.720 1.090 18.440 1.330 ;
        RECT  13.720 0.710 13.960 1.330 ;
        RECT  9.560 0.710 13.960 0.950 ;
        RECT  9.400 3.780 14.120 4.020 ;
        RECT  13.880 3.430 14.120 4.020 ;
        RECT  9.400 3.540 9.800 4.020 ;
        RECT  13.880 3.430 18.440 3.670 ;
        RECT  0.160 3.780 4.160 4.020 ;
        RECT  3.920 2.330 4.160 4.020 ;
        RECT  0.160 1.570 0.400 4.020 ;
        RECT  3.920 2.330 5.870 2.570 ;
        RECT  0.160 1.570 2.000 1.810 ;
        RECT  2.480 1.570 4.160 1.810 ;
        RECT  2.480 1.090 2.720 1.810 ;
        RECT  0.880 1.090 2.720 1.330 ;
    END
END MOAI1HT

MACRO MOAI1S
    CLASS CORE ;
    FOREIGN MOAI1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.230 0.620 3.600 1.020 ;
        RECT  3.240 1.490 3.600 1.890 ;
        RECT  3.270 0.620 3.600 2.200 ;
        RECT  3.360 0.620 3.600 3.760 ;
        RECT  1.970 3.520 3.600 3.760 ;
        RECT  1.970 3.360 2.210 3.760 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.420 1.160 2.820 ;
        RECT  0.790 2.200 1.070 2.860 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.210 0.480 2.610 ;
        RECT  0.170 2.210 0.450 3.010 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 0.880 2.930 3.020 ;
        RECT  2.650 2.620 3.120 3.020 ;
        RECT  2.630 0.880 2.930 1.280 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.440 2.400 2.840 ;
        RECT  2.030 2.200 2.310 2.860 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  1.080 -0.380 1.480 0.960 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.150 4.480 3.550 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.300 4.480 1.390 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.430 4.000 2.060 4.240 ;
        RECT  1.430 1.260 1.670 4.240 ;
        RECT  0.440 3.540 0.840 3.880 ;
        RECT  0.440 3.540 1.670 3.780 ;
        RECT  0.240 1.260 1.670 1.500 ;
        RECT  0.240 0.720 0.480 1.500 ;
    END
END MOAI1S

MACRO MULBE
    CLASS CORE ;
    FOREIGN MULBE 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN M
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 1.280 7.270 3.640 ;
        RECT  6.990 2.880 7.330 3.280 ;
        RECT  6.440 1.280 7.270 1.520 ;
        END
    END M
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.110 2.880 10.350 4.010 ;
        RECT  10.480 1.280 10.970 1.520 ;
        RECT  10.730 1.280 10.970 3.120 ;
        RECT  9.990 2.880 10.970 3.120 ;
        RECT  9.990 2.880 10.350 3.280 ;
        END
    END Z
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.870 2.130 9.110 3.150 ;
        RECT  8.870 2.250 9.730 2.650 ;
        RECT  8.700 2.130 9.110 2.530 ;
        END
    END M2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 1.280 5.410 3.640 ;
        RECT  5.130 2.880 5.470 3.280 ;
        RECT  4.580 1.280 5.410 1.520 ;
        END
    END S
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 2.250 0.510 2.650 ;
        RECT  0.190 3.750 2.650 3.990 ;
        RECT  2.250 3.750 2.650 4.260 ;
        RECT  0.190 2.250 0.430 3.990 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.710 2.190 3.110 2.640 ;
        RECT  1.310 2.400 3.110 2.640 ;
        RECT  1.310 2.250 1.550 2.650 ;
        END
    END M0
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.990 -0.380 3.390 0.560 ;
        RECT  5.720 -0.380 6.120 0.560 ;
        RECT  7.580 -0.380 7.980 0.560 ;
        RECT  8.340 -0.380 8.740 0.560 ;
        RECT  9.340 -0.380 9.740 0.560 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 4.230 1.700 5.420 ;
        RECT  2.890 4.260 3.290 5.420 ;
        RECT  3.920 4.480 4.860 5.420 ;
        RECT  6.080 4.480 6.480 5.420 ;
        RECT  8.340 3.980 8.740 5.420 ;
        RECT  7.940 4.480 8.740 5.420 ;
        RECT  9.220 4.480 9.620 5.420 ;
        RECT  10.600 4.480 11.000 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.170 4.230 0.570 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.810 0.800 1.050 3.260 ;
        RECT  5.770 0.800 6.010 2.650 ;
        RECT  10.230 1.760 10.470 2.640 ;
        RECT  9.890 1.760 10.470 2.000 ;
        RECT  9.890 0.800 10.130 2.000 ;
        RECT  1.300 0.800 1.700 1.400 ;
        RECT  0.810 0.800 1.700 1.280 ;
        RECT  0.810 0.800 10.130 1.040 ;
        RECT  8.220 2.790 8.630 3.190 ;
        RECT  8.220 1.490 8.460 3.190 ;
        RECT  7.630 2.250 8.460 2.650 ;
        RECT  8.220 1.490 8.620 1.890 ;
        RECT  4.650 4.000 6.750 4.240 ;
        RECT  6.510 2.250 6.750 4.240 ;
        RECT  4.650 2.250 4.890 4.240 ;
        RECT  3.940 2.790 4.190 3.190 ;
        RECT  3.950 1.490 4.190 3.190 ;
        RECT  3.950 2.410 4.890 2.650 ;
        RECT  3.940 1.490 4.190 1.890 ;
        RECT  2.020 3.170 3.620 3.410 ;
        RECT  3.380 1.710 3.620 3.410 ;
        RECT  3.380 2.130 3.710 2.530 ;
        RECT  2.300 1.710 3.620 1.950 ;
        RECT  2.300 1.570 2.700 1.950 ;
    END
END MULBE

MACRO MULBEP
    CLASS CORE ;
    FOREIGN MULBEP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN M
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.710 2.960 10.510 3.200 ;
        RECT  7.920 1.370 11.020 1.610 ;
        RECT  8.850 1.370 9.130 3.200 ;
        END
    END M
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.240 1.330 15.340 1.570 ;
        RECT  15.070 1.330 15.310 3.540 ;
        RECT  12.950 3.300 15.310 3.540 ;
        RECT  14.940 1.330 15.340 1.600 ;
        RECT  12.950 3.300 13.190 3.700 ;
        END
    END Z
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 1.820 12.230 3.430 ;
        RECT  13.190 1.820 13.470 2.580 ;
        RECT  13.190 1.820 13.820 2.350 ;
        RECT  11.780 1.820 14.250 2.100 ;
        RECT  11.780 1.820 12.230 2.450 ;
        END
    END M2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.050 2.960 6.850 3.200 ;
        RECT  4.500 1.370 7.600 1.610 ;
        RECT  5.130 1.370 5.410 3.200 ;
        END
    END S
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 2.250 0.480 2.650 ;
        RECT  0.190 0.930 2.120 1.170 ;
        RECT  0.190 0.930 0.430 3.640 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.630 2.190 3.030 2.660 ;
        RECT  1.250 2.380 3.030 2.660 ;
        RECT  1.250 2.240 1.490 2.660 ;
        END
    END M0
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.750 -0.380 4.230 0.560 ;
        RECT  5.850 -0.380 6.250 0.560 ;
        RECT  9.270 -0.380 9.670 0.560 ;
        RECT  11.340 -0.380 11.740 0.560 ;
        RECT  13.590 -0.380 13.990 0.560 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 4.400 1.620 5.420 ;
        RECT  2.750 4.480 4.780 5.420 ;
        RECT  5.760 4.480 6.160 5.420 ;
        RECT  7.140 4.480 8.420 5.420 ;
        RECT  9.400 4.480 9.800 5.420 ;
        RECT  10.800 4.480 11.200 5.420 ;
        RECT  11.460 4.400 11.860 5.420 ;
        RECT  12.180 4.480 12.580 5.420 ;
        RECT  13.560 4.480 13.960 5.420 ;
        RECT  14.940 4.480 15.340 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.160 4.230 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  12.800 0.800 14.780 1.040 ;
        RECT  14.380 0.670 14.780 1.040 ;
        RECT  12.800 0.670 13.200 1.040 ;
        RECT  1.200 3.920 12.710 4.160 ;
        RECT  12.470 2.340 12.710 4.160 ;
        RECT  1.200 3.650 1.440 4.160 ;
        RECT  0.770 3.650 1.440 3.890 ;
        RECT  0.770 1.570 1.010 3.890 ;
        RECT  12.470 2.820 14.730 3.060 ;
        RECT  14.490 2.030 14.730 3.060 ;
        RECT  12.470 2.340 12.870 2.580 ;
        RECT  0.770 1.570 1.700 1.810 ;
        RECT  11.300 2.790 11.700 3.190 ;
        RECT  11.300 1.290 11.540 3.190 ;
        RECT  9.370 1.850 9.770 2.350 ;
        RECT  9.370 1.850 11.540 2.090 ;
        RECT  11.300 1.290 11.740 1.530 ;
        RECT  4.420 3.440 11.060 3.680 ;
        RECT  10.820 2.330 11.060 3.680 ;
        RECT  8.140 2.250 8.380 3.680 ;
        RECT  7.090 2.330 7.330 3.680 ;
        RECT  4.420 2.250 4.660 3.680 ;
        RECT  3.860 2.950 4.810 3.190 ;
        RECT  3.860 2.790 4.110 3.190 ;
        RECT  3.870 1.490 4.110 3.190 ;
        RECT  8.140 2.250 8.610 2.650 ;
        RECT  4.420 2.250 4.810 2.650 ;
        RECT  10.580 2.330 11.060 2.570 ;
        RECT  6.910 2.330 7.330 2.570 ;
        RECT  3.860 1.490 4.110 1.890 ;
        RECT  8.480 0.800 10.460 1.040 ;
        RECT  10.060 0.670 10.460 1.040 ;
        RECT  8.480 0.670 8.880 1.040 ;
        RECT  7.660 1.850 7.900 3.200 ;
        RECT  5.760 1.850 6.160 2.350 ;
        RECT  5.760 1.850 7.900 2.090 ;
        RECT  5.060 0.800 7.040 1.040 ;
        RECT  6.640 0.670 7.040 1.040 ;
        RECT  5.060 0.670 5.460 1.040 ;
        RECT  1.940 3.170 3.540 3.410 ;
        RECT  3.300 1.570 3.540 3.410 ;
        RECT  3.300 2.130 3.630 2.530 ;
        RECT  2.220 1.570 3.540 1.810 ;
    END
END MULBEP

MACRO MULBET
    CLASS CORE ;
    FOREIGN MULBET 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 23.560 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN M
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.240 1.370 12.940 1.610 ;
        RECT  11.250 2.870 15.790 3.110 ;
        RECT  11.950 1.370 12.230 3.110 ;
        END
    END M
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  18.170 3.070 22.710 3.310 ;
        RECT  21.080 1.440 22.780 1.680 ;
        RECT  21.870 1.440 22.150 3.310 ;
        END
    END Z
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.530 2.110 17.930 2.350 ;
        RECT  17.530 2.110 17.810 3.410 ;
        END
    END M2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.120 1.370 6.820 1.610 ;
        RECT  5.010 2.870 9.490 3.110 ;
        RECT  5.750 1.370 6.030 3.110 ;
        END
    END S
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 2.250 0.480 2.650 ;
        RECT  0.190 0.930 2.120 1.170 ;
        RECT  0.190 0.930 0.430 3.640 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.630 2.190 3.030 2.660 ;
        RECT  1.250 2.380 3.030 2.660 ;
        RECT  1.250 2.240 1.490 2.660 ;
        END
    END M0
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.700 -0.380 4.180 0.560 ;
        RECT  7.890 -0.380 8.290 0.560 ;
        RECT  9.270 -0.380 9.670 0.560 ;
        RECT  14.010 -0.380 14.410 0.560 ;
        RECT  15.390 -0.380 15.790 0.560 ;
        RECT  16.740 -0.380 17.140 0.910 ;
        RECT  18.230 -0.380 18.630 0.560 ;
        RECT  19.610 -0.380 20.010 0.560 ;
        RECT  0.000 -0.380 23.560 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 4.400 1.620 5.420 ;
        RECT  2.700 4.480 3.100 5.420 ;
        RECT  4.320 4.480 4.720 5.420 ;
        RECT  5.700 4.480 6.100 5.420 ;
        RECT  7.080 4.480 7.480 5.420 ;
        RECT  8.460 4.480 8.860 5.420 ;
        RECT  9.840 4.480 10.240 5.420 ;
        RECT  10.560 4.480 10.960 5.420 ;
        RECT  11.940 4.480 12.340 5.420 ;
        RECT  13.320 4.480 13.720 5.420 ;
        RECT  14.700 4.480 15.100 5.420 ;
        RECT  16.080 4.400 17.140 5.420 ;
        RECT  17.480 4.480 17.880 5.420 ;
        RECT  18.860 4.480 19.260 5.420 ;
        RECT  20.240 4.480 20.640 5.420 ;
        RECT  21.620 4.480 22.020 5.420 ;
        RECT  23.000 4.480 23.400 5.420 ;
        RECT  0.000 4.660 23.560 5.420 ;
        RECT  0.160 4.230 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  17.580 1.570 20.640 1.810 ;
        RECT  20.400 0.620 20.640 1.810 ;
        RECT  20.400 0.620 23.400 0.860 ;
        RECT  0.770 3.650 23.190 3.890 ;
        RECT  22.950 2.110 23.190 3.890 ;
        RECT  9.730 2.330 10.010 3.890 ;
        RECT  0.770 1.570 1.010 3.890 ;
        RECT  9.440 2.330 10.010 2.570 ;
        RECT  22.790 2.110 23.190 2.350 ;
        RECT  0.770 1.570 1.700 1.810 ;
        RECT  16.790 1.490 17.030 3.190 ;
        RECT  15.970 2.330 17.030 2.570 ;
        RECT  16.790 1.490 17.060 1.890 ;
        RECT  13.380 1.570 16.420 1.810 ;
        RECT  13.380 0.620 13.620 1.810 ;
        RECT  10.620 0.620 13.620 0.860 ;
        RECT  10.880 1.850 11.280 2.570 ;
        RECT  6.760 1.850 7.000 2.430 ;
        RECT  6.760 1.850 11.280 2.090 ;
        RECT  7.260 1.370 10.300 1.610 ;
        RECT  7.260 0.620 7.500 1.610 ;
        RECT  4.500 0.620 7.500 0.860 ;
        RECT  3.860 2.790 4.110 3.190 ;
        RECT  3.870 1.490 4.110 3.190 ;
        RECT  3.870 2.030 4.660 2.430 ;
        RECT  3.860 1.490 4.110 1.890 ;
        RECT  1.940 3.170 3.540 3.410 ;
        RECT  3.300 1.570 3.540 3.410 ;
        RECT  3.300 2.130 3.630 2.530 ;
        RECT  2.220 1.570 3.540 1.810 ;
    END
END MULBET

MACRO MULPA
    CLASS CORE ;
    FOREIGN MULPA 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN M
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END M
    PIN Z
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.400 13.470 3.080 ;
        END
    END S
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.250 2.260 8.620 2.660 ;
        RECT  8.250 2.400 9.060 2.640 ;
        RECT  8.250 2.010 8.490 2.830 ;
        END
    END M0
    PIN P
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 1.180 14.710 3.310 ;
        RECT  14.400 2.910 14.710 3.310 ;
        RECT  14.400 1.490 14.710 1.890 ;
        END
    END P
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.060 -0.380 2.460 0.640 ;
        RECT  7.890 -0.380 9.910 0.560 ;
        RECT  13.610 -0.380 14.010 0.560 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.060 4.480 2.460 5.420 ;
        RECT  8.170 4.480 9.110 5.420 ;
        RECT  9.600 4.280 10.000 5.420 ;
        RECT  13.610 4.480 14.010 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.270 4.180 13.370 4.420 ;
        RECT  13.130 3.920 13.370 4.420 ;
        RECT  11.270 1.370 11.510 4.420 ;
        RECT  13.130 3.920 14.030 4.160 ;
        RECT  13.790 2.100 14.030 4.160 ;
        RECT  13.790 2.100 14.160 2.500 ;
        RECT  12.100 3.700 12.890 3.940 ;
        RECT  12.650 0.730 12.890 3.940 ;
        RECT  12.650 2.900 12.950 3.300 ;
        RECT  12.650 1.370 12.950 1.770 ;
        RECT  11.990 0.890 12.230 3.320 ;
        RECT  8.830 2.910 9.750 3.310 ;
        RECT  9.510 0.890 9.750 3.310 ;
        RECT  8.830 1.370 9.750 1.770 ;
        RECT  9.510 0.890 12.230 1.130 ;
        RECT  10.550 1.370 10.790 3.310 ;
        RECT  4.370 4.070 7.950 4.310 ;
        RECT  7.710 3.710 7.950 4.310 ;
        RECT  4.370 1.370 4.610 4.310 ;
        RECT  7.710 3.710 10.640 3.950 ;
        RECT  6.530 0.890 6.770 3.310 ;
        RECT  6.530 0.890 9.270 1.130 ;
        RECT  7.730 3.070 8.210 3.470 ;
        RECT  7.730 1.370 7.970 3.470 ;
        RECT  7.680 2.010 7.970 2.410 ;
        RECT  7.730 1.370 8.210 1.770 ;
        RECT  5.270 3.550 5.670 3.830 ;
        RECT  5.090 3.550 7.440 3.790 ;
        RECT  7.200 1.370 7.440 3.790 ;
        RECT  5.090 1.370 5.330 3.790 ;
        RECT  7.200 2.910 7.490 3.310 ;
        RECT  7.200 1.370 7.490 1.770 ;
        RECT  0.900 0.890 1.140 3.330 ;
        RECT  5.810 0.890 6.050 3.310 ;
        RECT  3.650 2.910 4.130 3.310 ;
        RECT  3.890 0.890 4.130 3.310 ;
        RECT  0.830 2.910 1.140 3.310 ;
        RECT  3.650 1.370 4.130 1.770 ;
        RECT  0.830 1.370 1.140 1.770 ;
        RECT  0.900 0.890 6.050 1.130 ;
        RECT  3.730 4.000 4.130 4.350 ;
        RECT  1.550 4.000 4.130 4.240 ;
        RECT  1.550 2.910 1.790 4.240 ;
        RECT  1.530 1.370 1.770 3.150 ;
        RECT  1.530 1.370 1.790 1.770 ;
        RECT  2.850 2.990 3.410 3.230 ;
        RECT  3.170 1.370 3.410 3.230 ;
        RECT  3.170 2.100 3.610 2.500 ;
        RECT  2.930 1.370 3.410 1.770 ;
    END
END MULPA

MACRO MULPAP
    CLASS CORE ;
    FOREIGN MULPAP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN M
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END M
    PIN Z
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.400 13.470 3.080 ;
        RECT  13.160 2.030 13.470 2.430 ;
        END
    END S
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.250 2.260 8.620 2.660 ;
        RECT  8.250 2.400 9.060 2.640 ;
        RECT  8.250 2.010 8.490 2.830 ;
        END
    END M0
    PIN P
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 1.180 14.710 3.310 ;
        RECT  14.350 2.910 14.710 3.310 ;
        RECT  14.350 1.490 14.710 1.890 ;
        END
    END P
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.060 -0.380 2.460 0.640 ;
        RECT  7.890 -0.380 9.910 0.560 ;
        RECT  13.560 -0.380 13.960 0.560 ;
        RECT  14.940 -0.380 15.340 0.560 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.060 4.480 2.460 5.420 ;
        RECT  8.170 4.480 9.110 5.420 ;
        RECT  9.600 4.280 10.000 5.420 ;
        RECT  13.560 4.480 13.960 5.420 ;
        RECT  14.940 4.480 15.340 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.270 4.180 13.320 4.420 ;
        RECT  13.080 3.920 13.320 4.420 ;
        RECT  11.270 1.370 11.510 4.420 ;
        RECT  13.080 3.920 13.980 4.160 ;
        RECT  13.740 2.100 13.980 4.160 ;
        RECT  13.740 2.100 14.080 2.500 ;
        RECT  12.100 3.700 12.840 3.940 ;
        RECT  12.600 0.730 12.840 3.940 ;
        RECT  12.600 2.900 12.950 3.300 ;
        RECT  12.600 1.370 12.950 1.770 ;
        RECT  12.520 0.730 12.840 1.130 ;
        RECT  11.990 0.890 12.230 3.320 ;
        RECT  8.830 2.910 9.750 3.310 ;
        RECT  9.510 0.890 9.750 3.310 ;
        RECT  8.830 1.370 9.750 1.770 ;
        RECT  9.510 0.890 12.230 1.130 ;
        RECT  10.550 1.370 10.790 3.310 ;
        RECT  4.370 4.070 7.950 4.310 ;
        RECT  7.710 3.710 7.950 4.310 ;
        RECT  4.370 1.370 4.610 4.310 ;
        RECT  7.710 3.710 10.640 3.950 ;
        RECT  6.530 0.890 6.770 3.310 ;
        RECT  6.530 0.890 9.270 1.130 ;
        RECT  7.730 3.070 8.210 3.470 ;
        RECT  7.730 1.370 7.970 3.470 ;
        RECT  7.680 2.010 7.970 2.410 ;
        RECT  7.730 1.370 8.210 1.770 ;
        RECT  5.270 3.550 5.670 3.830 ;
        RECT  5.090 3.550 7.440 3.790 ;
        RECT  7.200 1.370 7.440 3.790 ;
        RECT  5.090 1.370 5.330 3.790 ;
        RECT  7.200 2.910 7.490 3.310 ;
        RECT  7.200 1.370 7.490 1.770 ;
        RECT  0.900 0.890 1.140 3.330 ;
        RECT  5.810 0.890 6.050 3.310 ;
        RECT  3.650 2.910 4.130 3.310 ;
        RECT  3.890 0.890 4.130 3.310 ;
        RECT  0.830 2.910 1.140 3.310 ;
        RECT  3.650 1.370 4.130 1.770 ;
        RECT  0.830 1.370 1.140 1.770 ;
        RECT  0.900 0.890 6.050 1.130 ;
        RECT  3.730 4.000 4.130 4.350 ;
        RECT  1.550 4.000 4.130 4.240 ;
        RECT  1.550 2.910 1.790 4.240 ;
        RECT  1.530 1.370 1.770 3.150 ;
        RECT  1.530 1.370 1.790 1.770 ;
        RECT  2.850 2.990 3.410 3.230 ;
        RECT  3.170 1.370 3.410 3.230 ;
        RECT  3.170 2.100 3.610 2.500 ;
        RECT  2.930 1.370 3.410 1.770 ;
    END
END MULPAP

MACRO MULPAT
    CLASS CORE ;
    FOREIGN MULPAT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.740 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN M
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END M
    PIN Z
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.400 13.470 3.080 ;
        RECT  13.020 2.030 13.470 2.430 ;
        END
    END S
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.250 2.260 8.620 2.660 ;
        RECT  8.250 2.400 9.060 2.640 ;
        RECT  8.250 2.010 8.490 2.830 ;
        END
    END M0
    PIN P
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.290 1.180 14.570 3.310 ;
        RECT  14.210 2.910 14.570 3.310 ;
        RECT  15.590 1.490 15.950 1.890 ;
        RECT  14.290 2.410 15.950 2.650 ;
        RECT  15.670 1.180 15.950 3.310 ;
        RECT  15.590 2.910 15.950 3.310 ;
        RECT  14.210 1.490 14.570 1.890 ;
        END
    END P
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.060 -0.380 2.460 0.640 ;
        RECT  7.780 -0.380 9.800 0.560 ;
        RECT  13.420 -0.380 13.820 0.560 ;
        RECT  14.800 -0.380 15.200 0.560 ;
        RECT  16.180 -0.380 16.580 0.560 ;
        RECT  0.000 -0.380 16.740 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.060 4.480 2.460 5.420 ;
        RECT  8.170 4.480 9.110 5.420 ;
        RECT  9.540 4.280 9.940 5.420 ;
        RECT  13.420 4.480 13.820 5.420 ;
        RECT  14.800 4.480 15.200 5.420 ;
        RECT  16.180 4.480 16.580 5.420 ;
        RECT  0.000 4.660 16.740 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.130 4.180 13.180 4.420 ;
        RECT  12.940 3.920 13.180 4.420 ;
        RECT  11.130 1.370 11.370 4.420 ;
        RECT  12.940 3.920 13.950 4.160 ;
        RECT  13.710 2.100 13.950 4.160 ;
        RECT  13.710 2.100 14.050 2.500 ;
        RECT  11.960 3.700 12.700 3.940 ;
        RECT  12.460 0.730 12.700 3.940 ;
        RECT  12.460 2.900 12.810 3.300 ;
        RECT  12.460 1.370 12.810 1.770 ;
        RECT  12.380 0.730 12.700 1.130 ;
        RECT  11.850 0.890 12.090 3.320 ;
        RECT  8.830 2.910 9.750 3.310 ;
        RECT  9.510 0.890 9.750 3.310 ;
        RECT  8.830 1.370 9.750 1.770 ;
        RECT  9.510 0.890 12.090 1.130 ;
        RECT  10.410 1.370 10.650 3.310 ;
        RECT  4.370 4.070 7.950 4.310 ;
        RECT  7.710 3.710 7.950 4.310 ;
        RECT  4.370 1.370 4.610 4.310 ;
        RECT  7.710 3.710 10.500 3.950 ;
        RECT  6.530 0.890 6.770 3.310 ;
        RECT  6.530 0.890 9.270 1.130 ;
        RECT  7.730 3.070 8.210 3.470 ;
        RECT  7.730 1.370 7.970 3.470 ;
        RECT  7.680 2.010 7.970 2.410 ;
        RECT  7.730 1.370 8.210 1.770 ;
        RECT  5.270 3.550 5.670 3.830 ;
        RECT  5.090 3.550 7.440 3.790 ;
        RECT  7.200 1.370 7.440 3.790 ;
        RECT  5.090 1.370 5.330 3.790 ;
        RECT  7.200 2.910 7.490 3.310 ;
        RECT  7.200 1.370 7.490 1.770 ;
        RECT  0.900 0.890 1.140 3.330 ;
        RECT  5.810 0.890 6.050 3.310 ;
        RECT  3.650 2.910 4.130 3.310 ;
        RECT  3.890 0.890 4.130 3.310 ;
        RECT  0.830 2.910 1.140 3.310 ;
        RECT  3.650 1.370 4.130 1.770 ;
        RECT  0.830 1.370 1.140 1.770 ;
        RECT  0.900 0.890 6.050 1.130 ;
        RECT  3.730 4.000 4.130 4.350 ;
        RECT  1.550 4.000 4.130 4.240 ;
        RECT  1.550 2.910 1.790 4.240 ;
        RECT  1.530 1.370 1.770 3.150 ;
        RECT  1.530 1.370 1.790 1.770 ;
        RECT  2.850 2.990 3.410 3.230 ;
        RECT  3.170 1.370 3.410 3.230 ;
        RECT  3.170 2.100 3.610 2.500 ;
        RECT  2.930 1.370 3.410 1.770 ;
    END
END MULPAT

MACRO MUX2
    CLASS CORE ;
    FOREIGN MUX2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.130 4.180 2.020 ;
        RECT  3.900 1.130 4.180 3.110 ;
        RECT  3.780 2.870 4.180 3.110 ;
        RECT  3.860 1.490 4.180 1.890 ;
        END
    END O
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.500 1.070 3.780 ;
        RECT  0.830 3.500 1.070 4.420 ;
        RECT  0.170 3.420 0.450 3.780 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.200 0.490 2.600 ;
        RECT  0.170 1.640 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.700 3.830 4.170 4.110 ;
        RECT  3.890 3.420 4.170 4.110 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.080 -0.380 3.480 0.720 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.430 -0.380 0.830 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.460 4.470 3.370 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.140 4.050 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.790 3.350 3.520 3.590 ;
        RECT  3.280 2.230 3.520 3.590 ;
        RECT  1.790 1.490 2.030 3.590 ;
        RECT  3.280 2.230 3.660 2.630 ;
        RECT  2.430 2.870 2.910 3.110 ;
        RECT  2.670 1.570 2.910 3.110 ;
        RECT  2.430 1.570 2.910 1.810 ;
        RECT  1.310 4.170 1.790 4.410 ;
        RECT  1.310 0.640 1.550 4.410 ;
        RECT  1.290 0.750 1.690 0.990 ;
        RECT  1.860 0.620 2.260 0.880 ;
        RECT  1.310 0.640 2.260 0.880 ;
        RECT  0.830 1.490 1.070 3.190 ;
    END
END MUX2

MACRO MUX2F
    CLASS CORE ;
    FOREIGN MUX2F 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.220 4.790 3.190 ;
        RECT  4.440 2.790 4.790 3.190 ;
        RECT  5.720 1.220 6.030 1.900 ;
        RECT  4.510 1.620 6.030 1.900 ;
        RECT  5.750 1.220 6.030 3.190 ;
        RECT  5.720 2.790 6.030 3.190 ;
        RECT  4.480 1.220 4.790 1.620 ;
        END
    END O
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 3.900 1.530 4.300 ;
        RECT  0.790 3.430 1.070 4.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.200 0.530 2.600 ;
        RECT  0.170 2.200 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.520 4.170 2.610 ;
        RECT  3.380 2.030 4.170 2.430 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.100 -0.380 1.500 0.570 ;
        RECT  3.780 -0.380 4.180 0.860 ;
        RECT  5.000 -0.380 5.420 0.940 ;
        RECT  6.240 -0.380 6.660 0.940 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  0.160 -0.380 0.560 0.570 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.010 4.470 2.410 5.420 ;
        RECT  3.700 4.100 4.100 5.420 ;
        RECT  4.980 4.100 5.380 5.420 ;
        RECT  6.260 4.100 6.660 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  0.160 3.800 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.920 3.430 5.320 3.670 ;
        RECT  5.080 2.230 5.320 3.670 ;
        RECT  2.250 3.250 4.160 3.490 ;
        RECT  2.250 1.360 2.490 3.490 ;
        RECT  5.080 2.230 5.370 2.630 ;
        RECT  2.790 2.770 3.290 3.010 ;
        RECT  2.790 1.260 3.030 3.010 ;
        RECT  2.790 1.260 3.390 1.500 ;
        RECT  1.770 3.750 2.410 3.990 ;
        RECT  1.770 0.780 2.010 3.990 ;
        RECT  1.290 1.970 2.010 2.370 ;
        RECT  1.770 0.780 2.830 1.020 ;
        RECT  1.890 0.620 2.290 1.020 ;
        RECT  0.810 2.770 1.430 3.010 ;
        RECT  0.810 1.360 1.050 3.010 ;
        RECT  0.810 1.360 1.090 1.760 ;
    END
END MUX2F

MACRO MUX2P
    CLASS CORE ;
    FOREIGN MUX2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.830 1.260 4.790 1.540 ;
        RECT  4.510 1.260 4.790 3.220 ;
        RECT  3.780 2.940 4.790 3.220 ;
        RECT  3.830 1.260 4.150 1.750 ;
        END
    END O
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.730 4.130 1.150 4.420 ;
        RECT  0.790 3.430 1.070 4.420 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.200 0.490 2.600 ;
        RECT  0.170 2.200 0.450 3.300 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 3.460 4.170 4.110 ;
        RECT  2.030 3.830 4.170 4.110 ;
        RECT  2.030 3.830 2.310 4.420 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 -0.380 2.940 1.030 ;
        RECT  2.520 -0.380 3.500 0.790 ;
        RECT  4.380 -0.380 4.800 1.020 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.430 -0.380 0.830 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.970 4.470 3.370 5.420 ;
        RECT  4.430 4.100 4.820 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.140 3.910 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.990 3.350 3.530 3.590 ;
        RECT  3.290 2.310 3.530 3.590 ;
        RECT  1.990 1.490 2.230 3.590 ;
        RECT  1.830 2.870 2.230 3.270 ;
        RECT  3.290 2.310 4.120 2.640 ;
        RECT  1.830 1.490 2.230 1.890 ;
        RECT  2.470 2.870 2.910 3.110 ;
        RECT  2.670 1.490 2.910 3.110 ;
        RECT  2.550 1.490 2.910 1.890 ;
        RECT  1.390 4.170 1.790 4.420 ;
        RECT  1.390 3.520 1.750 4.420 ;
        RECT  1.350 0.720 1.590 3.760 ;
        RECT  1.290 1.010 2.260 1.250 ;
        RECT  1.290 0.720 1.690 1.250 ;
        RECT  0.810 2.790 1.110 3.190 ;
        RECT  0.810 1.490 1.050 3.190 ;
        RECT  0.810 1.490 1.110 1.890 ;
    END
END MUX2P

MACRO MUX2S
    CLASS CORE ;
    FOREIGN MUX2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 0.650 4.170 3.700 ;
        RECT  3.860 3.300 4.170 3.700 ;
        RECT  3.860 0.650 4.170 1.050 ;
        END
    END O
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.880 1.040 4.120 ;
        RECT  0.800 3.880 1.040 4.420 ;
        RECT  0.800 4.180 2.320 4.420 ;
        RECT  0.170 3.420 0.450 4.120 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.830 0.480 2.230 ;
        RECT  0.170 1.640 0.450 2.280 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.190 3.550 2.840 ;
        RECT  3.130 2.190 3.550 2.590 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.060 0.690 3.500 0.930 ;
        RECT  3.260 -0.380 3.500 1.890 ;
        RECT  3.260 1.490 3.640 1.890 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.700 4.480 3.100 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.550 4.180 3.950 4.420 ;
        RECT  2.660 4.000 3.940 4.240 ;
        RECT  2.660 3.520 2.900 4.240 ;
        RECT  1.920 3.520 2.900 3.760 ;
        RECT  1.920 1.290 2.160 3.760 ;
        RECT  1.760 2.790 2.160 3.190 ;
        RECT  1.840 1.290 2.160 1.690 ;
        RECT  2.480 2.790 2.890 3.190 ;
        RECT  2.650 1.490 2.890 3.190 ;
        RECT  2.650 1.490 2.920 1.890 ;
        RECT  1.280 3.640 1.680 3.880 ;
        RECT  1.280 2.250 1.520 3.880 ;
        RECT  1.360 0.620 1.600 2.490 ;
        RECT  1.360 0.620 2.700 0.860 ;
        RECT  0.790 1.290 1.030 3.190 ;
        RECT  0.790 1.290 1.120 1.690 ;
    END
END MUX2S

MACRO MUX2T
    CLASS CORE ;
    FOREIGN MUX2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.360 4.790 3.190 ;
        RECT  4.480 2.790 4.790 3.190 ;
        RECT  5.720 1.360 6.030 1.760 ;
        RECT  5.750 1.360 6.030 3.190 ;
        RECT  5.720 2.790 6.030 3.190 ;
        RECT  4.480 1.480 6.040 1.760 ;
        RECT  4.480 1.360 4.790 1.760 ;
        END
    END O
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 3.900 1.530 4.300 ;
        RECT  0.790 3.420 1.070 4.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.200 0.530 2.600 ;
        RECT  0.170 2.200 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.520 4.170 2.610 ;
        RECT  3.430 2.030 4.170 2.430 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.100 -0.380 1.500 0.570 ;
        RECT  3.780 -0.380 4.180 0.860 ;
        RECT  5.000 -0.380 5.420 0.940 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.160 -0.380 0.560 0.570 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.010 4.470 2.410 5.420 ;
        RECT  3.880 4.100 4.280 5.420 ;
        RECT  5.130 4.100 5.530 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.240 3.800 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.960 3.550 5.300 3.790 ;
        RECT  5.060 2.230 5.300 3.790 ;
        RECT  3.960 3.250 4.200 3.790 ;
        RECT  2.250 3.250 4.200 3.490 ;
        RECT  2.250 1.360 2.490 3.490 ;
        RECT  2.790 2.770 3.290 3.010 ;
        RECT  2.790 1.260 3.030 3.010 ;
        RECT  2.790 1.260 3.390 1.500 ;
        RECT  1.770 3.750 2.410 3.990 ;
        RECT  1.770 0.780 2.010 3.990 ;
        RECT  1.320 1.960 2.010 2.360 ;
        RECT  1.770 0.780 2.830 1.020 ;
        RECT  1.890 0.620 2.290 1.020 ;
        RECT  0.840 2.770 1.350 3.010 ;
        RECT  0.840 1.440 1.080 3.010 ;
        RECT  0.840 1.440 1.280 1.680 ;
    END
END MUX2T

MACRO MUX3
    CLASS CORE ;
    FOREIGN MUX3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 2.790 7.270 3.860 ;
        RECT  7.050 1.490 7.290 3.310 ;
        RECT  6.960 2.910 7.290 3.310 ;
        RECT  6.960 1.490 7.290 1.890 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.440 1.070 3.720 ;
        RECT  0.780 3.440 1.070 4.420 ;
        RECT  0.750 4.180 1.150 4.420 ;
        RECT  0.170 3.210 0.450 3.720 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 3.430 6.650 4.010 ;
        RECT  5.810 3.630 6.650 3.870 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.050 0.490 2.450 ;
        RECT  0.170 1.830 0.450 2.620 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.000 2.040 3.550 2.440 ;
        RECT  3.270 1.610 3.550 2.440 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 3.630 4.170 3.910 ;
        RECT  3.930 3.630 4.170 4.180 ;
        RECT  3.270 3.420 3.550 3.910 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.030 -0.380 3.430 0.560 ;
        RECT  6.040 -0.380 6.600 0.770 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.430 -0.380 0.830 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.260 4.150 3.660 5.420 ;
        RECT  5.910 4.480 6.310 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.140 4.110 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.940 2.790 5.320 3.190 ;
        RECT  5.080 1.010 5.320 3.190 ;
        RECT  6.390 2.150 6.810 2.550 ;
        RECT  6.390 1.010 6.630 2.550 ;
        RECT  4.940 1.490 5.320 1.890 ;
        RECT  5.080 1.010 6.630 1.250 ;
        RECT  5.660 2.790 6.010 3.190 ;
        RECT  5.770 1.490 6.010 3.190 ;
        RECT  5.660 1.490 6.010 1.890 ;
        RECT  4.490 4.170 4.890 4.420 ;
        RECT  4.490 3.520 4.730 4.420 ;
        RECT  4.460 0.700 4.700 3.760 ;
        RECT  4.460 2.030 4.740 2.430 ;
        RECT  4.270 0.700 4.700 1.140 ;
        RECT  3.970 1.380 4.210 3.390 ;
        RECT  1.790 1.100 2.030 3.200 ;
        RECT  3.790 0.800 4.030 1.620 ;
        RECT  1.790 1.100 2.890 1.340 ;
        RECT  2.650 0.800 2.890 1.340 ;
        RECT  2.650 0.800 4.030 1.040 ;
        RECT  2.510 1.580 2.750 3.200 ;
        RECT  2.430 1.580 2.830 1.820 ;
        RECT  1.390 4.170 1.790 4.410 ;
        RECT  1.390 3.430 1.630 4.410 ;
        RECT  1.310 0.620 1.550 3.740 ;
        RECT  1.310 0.620 2.340 0.860 ;
        RECT  0.810 1.490 1.050 3.200 ;
        RECT  0.810 1.490 1.070 1.890 ;
    END
END MUX3

MACRO MUX3P
    CLASS CORE ;
    FOREIGN MUX3P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.060 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.960 1.260 7.890 1.540 ;
        RECT  7.610 1.260 7.890 3.220 ;
        RECT  6.920 2.940 7.890 3.220 ;
        RECT  6.960 1.260 7.200 1.890 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.440 1.070 3.720 ;
        RECT  0.780 3.440 1.070 4.420 ;
        RECT  0.730 4.130 1.150 4.420 ;
        RECT  0.170 3.230 0.450 3.720 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 3.290 6.650 4.100 ;
        RECT  5.810 3.630 6.650 3.870 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.030 0.490 2.430 ;
        RECT  0.170 1.620 0.450 2.430 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.000 2.040 3.550 2.440 ;
        RECT  3.270 1.610 3.550 2.440 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 3.630 4.170 3.910 ;
        RECT  3.930 3.630 4.170 4.180 ;
        RECT  3.270 3.420 3.550 3.910 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.030 -0.380 3.430 0.560 ;
        RECT  6.040 -0.380 6.600 0.770 ;
        RECT  7.500 -0.380 7.900 0.990 ;
        RECT  0.000 -0.380 8.060 0.380 ;
        RECT  0.430 -0.380 0.830 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.260 4.150 3.660 5.420 ;
        RECT  5.480 4.480 6.380 5.420 ;
        RECT  7.500 4.210 7.900 5.420 ;
        RECT  0.000 4.660 8.060 5.420 ;
        RECT  0.160 4.110 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.940 2.790 5.320 3.190 ;
        RECT  5.080 1.010 5.320 3.190 ;
        RECT  6.390 2.150 6.810 2.550 ;
        RECT  6.390 1.010 6.630 2.550 ;
        RECT  4.940 1.490 5.320 1.890 ;
        RECT  5.080 1.010 6.630 1.250 ;
        RECT  5.660 2.790 6.010 3.190 ;
        RECT  5.770 1.490 6.010 3.190 ;
        RECT  5.660 1.490 6.010 1.890 ;
        RECT  4.490 4.170 4.890 4.420 ;
        RECT  4.490 3.520 4.730 4.420 ;
        RECT  4.460 0.700 4.700 3.760 ;
        RECT  4.460 2.030 4.740 2.430 ;
        RECT  4.270 0.700 4.700 1.140 ;
        RECT  3.970 1.380 4.210 3.390 ;
        RECT  1.790 2.800 2.110 3.200 ;
        RECT  1.870 1.100 2.110 3.200 ;
        RECT  1.790 1.500 2.110 1.900 ;
        RECT  3.790 0.800 4.030 1.620 ;
        RECT  1.870 1.100 2.890 1.340 ;
        RECT  2.650 0.800 2.890 1.340 ;
        RECT  2.650 0.800 4.030 1.040 ;
        RECT  2.510 1.580 2.750 3.200 ;
        RECT  2.430 1.580 2.830 1.820 ;
        RECT  1.390 4.170 1.790 4.410 ;
        RECT  1.390 3.430 1.630 4.410 ;
        RECT  1.310 0.620 1.550 3.740 ;
        RECT  1.310 0.620 2.340 0.860 ;
        RECT  0.810 1.490 1.050 3.200 ;
        RECT  0.810 1.490 1.070 1.890 ;
    END
END MUX3P

MACRO MUX3S
    CLASS CORE ;
    FOREIGN MUX3S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.680 3.660 7.270 4.060 ;
        RECT  6.990 0.630 7.270 2.660 ;
        RECT  6.990 3.500 7.270 4.080 ;
        RECT  7.040 2.380 7.320 3.780 ;
        RECT  6.960 0.630 7.270 1.030 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.960 1.070 4.240 ;
        RECT  0.830 3.960 1.070 4.420 ;
        RECT  0.170 3.380 0.450 4.240 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.350 2.130 6.670 2.740 ;
        RECT  6.320 2.170 6.670 2.570 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.160 0.480 2.560 ;
        RECT  0.170 1.980 0.450 2.620 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.640 3.750 2.960 4.150 ;
        RECT  2.640 3.420 2.930 4.310 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.260 3.730 2.660 ;
        RECT  3.270 2.130 3.550 2.840 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.900 -0.380 3.300 0.560 ;
        RECT  6.240 0.630 6.610 1.030 ;
        RECT  6.330 -0.380 6.610 1.890 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.500 -0.380 0.900 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.530 4.070 3.930 5.420 ;
        RECT  6.180 3.020 6.440 5.420 ;
        RECT  6.180 3.020 6.760 3.260 ;
        RECT  6.180 4.480 7.000 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.700 3.820 5.940 4.220 ;
        RECT  5.090 3.820 5.940 4.060 ;
        RECT  5.090 3.350 5.330 4.060 ;
        RECT  4.930 1.480 5.170 3.590 ;
        RECT  5.650 1.490 5.890 3.190 ;
        RECT  4.450 4.160 4.850 4.400 ;
        RECT  4.450 0.620 4.690 4.400 ;
        RECT  3.840 0.620 4.690 0.860 ;
        RECT  3.860 3.170 4.210 3.570 ;
        RECT  3.970 1.100 4.210 3.570 ;
        RECT  1.810 1.100 2.050 3.200 ;
        RECT  1.810 1.100 4.210 1.340 ;
        RECT  2.460 2.880 2.860 3.120 ;
        RECT  2.540 1.580 2.780 3.120 ;
        RECT  2.460 1.580 2.860 1.820 ;
        RECT  1.390 4.170 1.790 4.410 ;
        RECT  1.390 3.490 1.630 4.410 ;
        RECT  1.330 0.620 1.570 3.740 ;
        RECT  1.330 0.620 2.550 0.860 ;
        RECT  0.840 1.490 1.080 3.200 ;
    END
END MUX3S

MACRO MUX3T
    CLASS CORE ;
    FOREIGN MUX3T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.920 1.490 7.230 1.890 ;
        RECT  7.610 1.530 7.890 3.220 ;
        RECT  6.920 1.530 8.520 1.810 ;
        RECT  6.960 2.940 8.520 3.220 ;
        RECT  6.960 2.800 7.200 3.220 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.880 1.070 4.160 ;
        RECT  0.730 4.130 1.150 4.420 ;
        RECT  0.170 3.420 0.450 4.160 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 3.420 6.650 4.110 ;
        RECT  5.770 3.630 6.650 3.870 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.160 0.490 2.560 ;
        RECT  0.170 1.980 0.450 2.620 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.970 2.040 3.550 2.440 ;
        RECT  3.270 1.610 3.550 2.440 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 3.630 4.170 3.910 ;
        RECT  3.930 3.630 4.170 4.180 ;
        RECT  3.270 3.420 3.550 3.910 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.030 -0.380 3.430 0.560 ;
        RECT  6.000 -0.380 6.560 0.770 ;
        RECT  7.460 -0.380 7.860 0.990 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  0.430 -0.380 0.830 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.260 4.150 3.660 5.420 ;
        RECT  5.340 4.480 6.290 5.420 ;
        RECT  7.460 4.140 7.860 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.240 4.400 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.900 2.790 5.280 3.190 ;
        RECT  5.040 1.010 5.280 3.190 ;
        RECT  6.350 2.220 6.770 2.620 ;
        RECT  6.350 1.010 6.590 2.620 ;
        RECT  4.900 1.490 5.280 1.890 ;
        RECT  5.040 1.010 6.590 1.250 ;
        RECT  5.620 2.790 5.970 3.190 ;
        RECT  5.730 1.490 5.970 3.190 ;
        RECT  5.620 1.490 5.970 1.890 ;
        RECT  4.450 4.170 4.850 4.420 ;
        RECT  4.450 3.520 4.690 4.420 ;
        RECT  4.420 0.670 4.660 3.760 ;
        RECT  4.420 2.030 4.700 2.430 ;
        RECT  4.310 0.670 4.660 1.070 ;
        RECT  3.930 1.380 4.170 3.390 ;
        RECT  1.790 2.800 2.110 3.200 ;
        RECT  1.870 1.100 2.110 3.200 ;
        RECT  1.790 1.500 2.110 1.900 ;
        RECT  3.830 0.800 4.070 1.620 ;
        RECT  1.870 1.100 2.890 1.340 ;
        RECT  2.650 0.800 2.890 1.340 ;
        RECT  2.650 0.800 4.070 1.040 ;
        RECT  2.430 2.800 2.750 3.200 ;
        RECT  2.430 1.580 2.670 3.200 ;
        RECT  2.430 1.580 2.830 1.820 ;
        RECT  1.390 4.170 1.790 4.410 ;
        RECT  1.390 3.430 1.630 4.410 ;
        RECT  1.310 0.620 1.550 3.740 ;
        RECT  1.310 0.620 2.340 0.860 ;
        RECT  0.810 1.490 1.050 3.200 ;
        RECT  0.810 1.490 1.070 1.890 ;
    END
END MUX3T

MACRO MUX4
    CLASS CORE ;
    FOREIGN MUX4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.640 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.180 13.470 3.310 ;
        RECT  13.160 2.910 13.470 3.310 ;
        RECT  13.160 1.490 13.470 1.890 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.610 2.100 7.890 2.740 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.270 8.570 2.670 ;
        RECT  8.230 2.270 8.510 2.950 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.100 12.230 2.740 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.060 -0.380 2.460 0.640 ;
        RECT  7.930 -0.380 8.330 0.640 ;
        RECT  12.370 -0.380 12.770 0.560 ;
        RECT  0.000 -0.380 13.640 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.060 4.480 2.460 5.420 ;
        RECT  7.940 4.480 8.340 5.420 ;
        RECT  12.370 4.480 12.770 5.420 ;
        RECT  0.000 4.660 13.640 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.220 3.550 12.920 3.790 ;
        RECT  12.680 2.100 12.920 3.790 ;
        RECT  10.220 1.370 10.460 3.790 ;
        RECT  11.470 2.990 11.980 3.230 ;
        RECT  11.470 1.100 11.710 3.230 ;
        RECT  11.310 2.100 11.710 2.500 ;
        RECT  11.470 1.100 11.900 1.500 ;
        RECT  10.830 2.910 11.180 3.310 ;
        RECT  6.610 0.880 6.850 3.310 ;
        RECT  10.830 0.880 11.070 3.310 ;
        RECT  10.830 1.370 11.180 1.770 ;
        RECT  6.530 1.370 6.850 1.770 ;
        RECT  6.610 0.880 11.070 1.120 ;
        RECT  4.370 4.030 7.710 4.270 ;
        RECT  9.500 1.370 9.740 4.190 ;
        RECT  7.470 3.950 9.740 4.190 ;
        RECT  4.370 1.370 4.610 4.270 ;
        RECT  4.370 2.910 4.680 3.310 ;
        RECT  5.890 3.550 7.280 3.790 ;
        RECT  7.040 3.470 9.020 3.710 ;
        RECT  8.780 2.910 9.020 3.710 ;
        RECT  5.890 1.370 6.130 3.790 ;
        RECT  8.820 1.370 9.060 3.310 ;
        RECT  8.760 1.370 9.060 1.770 ;
        RECT  5.810 1.370 6.130 1.770 ;
        RECT  7.130 2.990 7.650 3.230 ;
        RECT  7.130 1.370 7.370 3.230 ;
        RECT  7.130 1.370 7.490 1.770 ;
        RECT  5.090 2.910 5.400 3.310 ;
        RECT  0.830 2.910 1.140 3.310 ;
        RECT  0.900 0.890 1.140 3.310 ;
        RECT  5.090 0.890 5.330 3.310 ;
        RECT  0.830 1.370 1.140 1.770 ;
        RECT  0.900 0.890 5.330 1.130 ;
        RECT  1.550 3.540 3.890 3.780 ;
        RECT  3.650 2.910 3.890 3.780 ;
        RECT  1.550 2.910 1.790 3.780 ;
        RECT  3.890 1.370 4.130 3.310 ;
        RECT  1.530 1.370 1.770 3.150 ;
        RECT  3.650 1.370 4.130 1.770 ;
        RECT  1.530 1.370 1.790 1.770 ;
        RECT  2.850 2.990 3.410 3.230 ;
        RECT  3.170 1.370 3.410 3.230 ;
        RECT  3.170 2.100 3.610 2.500 ;
        RECT  2.930 1.370 3.410 1.770 ;
    END
END MUX4

MACRO MUX4P
    CLASS CORE ;
    FOREIGN MUX4P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.300 2.790 14.710 3.190 ;
        RECT  14.430 1.180 14.710 3.300 ;
        RECT  14.300 1.490 14.710 1.890 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.100 8.510 2.740 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 2.100 9.270 2.500 ;
        RECT  8.850 2.100 9.130 2.740 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 2.100 13.470 2.740 ;
        RECT  13.160 2.100 13.470 2.500 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 -0.380 2.600 0.560 ;
        RECT  8.720 -0.380 9.120 0.560 ;
        RECT  13.500 -0.380 13.900 0.950 ;
        RECT  14.940 -0.380 15.340 1.030 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 4.480 2.600 5.420 ;
        RECT  8.720 4.480 9.120 5.420 ;
        RECT  13.500 4.260 13.900 5.420 ;
        RECT  14.940 4.180 15.340 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.000 3.780 14.060 4.020 ;
        RECT  13.820 2.100 14.060 4.020 ;
        RECT  11.000 1.370 11.240 4.020 ;
        RECT  13.820 2.100 14.080 2.500 ;
        RECT  12.440 1.490 12.680 3.310 ;
        RECT  11.720 0.800 11.960 3.310 ;
        RECT  6.680 2.990 7.080 3.230 ;
        RECT  6.760 0.800 7.000 3.230 ;
        RECT  6.760 0.800 11.960 1.040 ;
        RECT  4.600 4.000 10.520 4.240 ;
        RECT  10.280 1.370 10.520 4.240 ;
        RECT  4.600 1.370 4.840 4.240 ;
        RECT  6.040 3.520 9.800 3.760 ;
        RECT  9.560 1.490 9.800 3.760 ;
        RECT  6.040 1.370 6.280 3.760 ;
        RECT  7.550 1.490 7.790 3.190 ;
        RECT  0.830 0.800 1.070 3.380 ;
        RECT  5.320 0.800 5.560 3.310 ;
        RECT  0.830 0.800 5.560 1.040 ;
        RECT  1.530 4.000 4.120 4.240 ;
        RECT  3.880 1.370 4.120 4.240 ;
        RECT  1.530 1.490 1.770 4.240 ;
        RECT  1.530 2.980 1.790 3.380 ;
        RECT  1.530 1.490 1.790 1.890 ;
        RECT  3.160 2.880 3.530 3.280 ;
        RECT  3.290 1.490 3.530 3.280 ;
        RECT  3.290 2.100 3.610 2.500 ;
        RECT  3.160 1.490 3.530 1.890 ;
    END
END MUX4P

MACRO MUX4S
    CLASS CORE ;
    FOREIGN MUX4S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.640 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.180 13.470 3.310 ;
        RECT  13.160 2.910 13.470 3.310 ;
        RECT  13.160 1.490 13.470 1.890 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.610 2.100 7.890 2.740 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.370 8.570 2.770 ;
        RECT  8.230 2.300 8.510 2.950 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.100 12.230 2.740 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.060 -0.380 2.460 0.640 ;
        RECT  7.930 -0.380 8.330 0.640 ;
        RECT  12.370 -0.380 12.770 0.940 ;
        RECT  0.000 -0.380 13.640 0.380 ;
        RECT  0.160 -0.380 0.560 0.930 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.060 4.110 2.460 5.420 ;
        RECT  7.940 4.430 8.340 5.420 ;
        RECT  12.370 4.030 12.770 5.420 ;
        RECT  0.000 4.660 13.640 5.420 ;
        RECT  0.160 4.110 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.220 3.550 12.920 3.790 ;
        RECT  12.680 2.100 12.920 3.790 ;
        RECT  10.220 1.370 10.460 3.790 ;
        RECT  11.470 2.990 11.980 3.230 ;
        RECT  11.470 1.100 11.710 3.230 ;
        RECT  11.310 2.100 11.710 2.500 ;
        RECT  11.470 1.100 11.900 1.500 ;
        RECT  10.830 2.910 11.180 3.310 ;
        RECT  6.610 0.880 6.850 3.310 ;
        RECT  10.830 0.880 11.070 3.310 ;
        RECT  10.830 1.370 11.180 1.770 ;
        RECT  6.530 1.370 6.850 1.770 ;
        RECT  6.610 0.880 11.070 1.120 ;
        RECT  4.370 4.030 7.710 4.270 ;
        RECT  9.500 1.370 9.740 4.190 ;
        RECT  7.470 3.950 9.740 4.190 ;
        RECT  4.370 1.370 4.610 4.270 ;
        RECT  4.370 2.910 4.680 3.310 ;
        RECT  5.890 3.550 7.280 3.790 ;
        RECT  7.040 3.470 9.020 3.710 ;
        RECT  8.780 2.910 9.020 3.710 ;
        RECT  5.890 1.370 6.130 3.790 ;
        RECT  8.820 1.370 9.060 3.310 ;
        RECT  8.760 1.370 9.060 1.770 ;
        RECT  5.810 1.370 6.130 1.770 ;
        RECT  7.130 2.990 7.650 3.230 ;
        RECT  7.130 1.370 7.370 3.230 ;
        RECT  7.130 1.370 7.490 1.770 ;
        RECT  5.090 2.910 5.400 3.310 ;
        RECT  0.830 2.910 1.140 3.310 ;
        RECT  0.900 0.890 1.140 3.310 ;
        RECT  5.090 0.890 5.330 3.310 ;
        RECT  0.830 1.370 1.140 1.770 ;
        RECT  0.900 0.890 5.330 1.130 ;
        RECT  1.550 3.540 3.890 3.780 ;
        RECT  3.650 2.910 3.890 3.780 ;
        RECT  1.550 2.910 1.790 3.780 ;
        RECT  3.890 1.370 4.130 3.310 ;
        RECT  1.530 1.370 1.770 3.150 ;
        RECT  3.650 1.370 4.130 1.770 ;
        RECT  1.530 1.370 1.790 1.770 ;
        RECT  2.850 2.990 3.410 3.230 ;
        RECT  3.170 1.370 3.410 3.230 ;
        RECT  3.170 2.100 3.610 2.500 ;
        RECT  2.930 1.370 3.410 1.770 ;
    END
END MUX4S

MACRO MUX4T
    CLASS CORE ;
    FOREIGN MUX4T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.200 2.790 14.440 3.190 ;
        RECT  15.050 1.570 15.330 3.110 ;
        RECT  14.200 1.570 15.960 1.810 ;
        RECT  14.200 2.870 15.960 3.110 ;
        RECT  14.200 1.490 14.440 1.890 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.100 8.510 2.740 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 2.100 9.270 2.500 ;
        RECT  8.850 2.100 9.130 2.740 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 2.100 13.470 2.740 ;
        RECT  13.060 2.100 13.470 2.500 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 -0.380 2.600 0.560 ;
        RECT  8.720 -0.380 9.120 0.560 ;
        RECT  13.400 -0.380 13.800 1.110 ;
        RECT  14.840 -0.380 15.240 1.030 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 4.480 2.600 5.420 ;
        RECT  8.720 4.480 9.120 5.420 ;
        RECT  13.400 3.950 13.800 5.420 ;
        RECT  14.840 4.180 15.240 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.000 3.470 13.960 3.710 ;
        RECT  13.720 2.100 13.960 3.710 ;
        RECT  11.000 1.370 11.240 3.710 ;
        RECT  13.720 2.100 13.980 2.500 ;
        RECT  12.360 2.990 12.760 3.230 ;
        RECT  12.440 1.490 12.680 3.230 ;
        RECT  12.360 2.100 12.680 2.500 ;
        RECT  11.640 2.990 12.040 3.230 ;
        RECT  6.680 2.990 7.080 3.230 ;
        RECT  11.720 0.800 11.960 3.230 ;
        RECT  6.760 0.800 7.000 3.230 ;
        RECT  6.760 0.800 11.960 1.040 ;
        RECT  4.600 4.000 10.520 4.240 ;
        RECT  10.280 1.370 10.520 4.240 ;
        RECT  4.600 1.370 4.840 4.240 ;
        RECT  6.040 3.520 9.800 3.760 ;
        RECT  9.560 1.490 9.800 3.760 ;
        RECT  6.040 1.370 6.280 3.760 ;
        RECT  7.550 1.490 7.790 3.190 ;
        RECT  0.830 0.800 1.070 3.380 ;
        RECT  5.320 0.800 5.560 3.310 ;
        RECT  0.830 0.800 5.560 1.040 ;
        RECT  1.530 4.000 4.120 4.240 ;
        RECT  3.880 1.370 4.120 4.240 ;
        RECT  1.530 1.490 1.770 4.240 ;
        RECT  1.530 2.980 1.790 3.380 ;
        RECT  1.530 1.490 1.790 1.890 ;
        RECT  3.160 2.880 3.530 3.280 ;
        RECT  3.290 1.490 3.530 3.280 ;
        RECT  3.290 2.100 3.610 2.500 ;
        RECT  3.160 1.490 3.530 1.890 ;
    END
END MUX4T

MACRO MUXB2
    CLASS CORE ;
    FOREIGN MUXB2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.720 2.800 6.030 3.200 ;
        RECT  5.750 1.260 6.030 3.300 ;
        RECT  4.920 1.260 6.030 1.540 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.260 4.810 2.660 ;
        RECT  4.510 2.260 4.790 2.900 ;
        END
    END EB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.100 1.070 2.740 ;
        RECT  0.670 2.100 1.070 2.500 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.260 4.170 2.900 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.350 2.100 1.690 2.500 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.560 -0.380 6.040 0.560 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.640 -0.380 1.040 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.260 4.180 4.660 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  1.020 4.200 1.420 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.690 0.800 2.930 3.310 ;
        RECT  5.250 1.780 5.490 2.660 ;
        RECT  4.440 1.780 5.490 2.020 ;
        RECT  4.440 0.800 4.680 2.020 ;
        RECT  2.690 0.800 4.680 1.040 ;
        RECT  3.410 1.360 3.650 3.310 ;
        RECT  0.240 3.720 3.240 3.960 ;
        RECT  0.240 2.910 0.480 3.960 ;
        RECT  0.190 1.360 0.430 3.310 ;
        RECT  0.240 0.800 0.480 1.760 ;
        RECT  0.240 0.800 2.380 1.040 ;
        RECT  1.980 0.720 2.380 1.040 ;
        RECT  1.930 1.360 2.170 3.310 ;
    END
END MUXB2

MACRO MUXB2P
    CLASS CORE ;
    FOREIGN MUXB2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.060 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.830 1.290 7.180 1.530 ;
        RECT  6.060 3.220 7.900 3.460 ;
        RECT  6.370 1.290 6.650 3.460 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 2.250 5.410 2.900 ;
        END
    END EB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.100 1.070 2.740 ;
        RECT  0.670 2.100 1.070 2.500 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.250 4.170 2.900 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.350 2.100 1.690 2.500 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.120 -0.380 4.520 0.560 ;
        RECT  5.800 -0.380 6.200 0.560 ;
        RECT  7.500 -0.380 7.900 1.320 ;
        RECT  0.000 -0.380 8.060 0.380 ;
        RECT  0.640 -0.380 1.040 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.110 4.180 4.510 5.420 ;
        RECT  5.550 4.180 5.950 5.420 ;
        RECT  0.000 4.660 8.060 5.420 ;
        RECT  1.020 4.200 1.420 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.830 3.700 7.180 3.940 ;
        RECT  2.680 2.910 2.930 3.310 ;
        RECT  2.680 0.800 2.920 3.310 ;
        RECT  5.830 1.770 6.070 2.650 ;
        RECT  3.890 1.770 6.070 2.010 ;
        RECT  3.890 0.800 4.130 2.010 ;
        RECT  2.680 1.360 2.930 1.760 ;
        RECT  2.680 0.800 4.130 1.040 ;
        RECT  3.410 1.360 3.650 3.310 ;
        RECT  0.240 3.720 3.240 3.960 ;
        RECT  0.240 2.910 0.480 3.960 ;
        RECT  0.190 1.360 0.430 3.310 ;
        RECT  0.240 0.800 0.480 1.760 ;
        RECT  0.240 0.800 2.380 1.040 ;
        RECT  1.980 0.720 2.380 1.040 ;
        RECT  1.930 1.360 2.170 3.310 ;
    END
END MUXB2P

MACRO MUXB2S
    CLASS CORE ;
    FOREIGN MUXB2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.260 6.030 3.310 ;
        RECT  5.720 2.910 6.030 3.310 ;
        RECT  4.920 1.260 6.030 1.540 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.260 4.810 2.660 ;
        RECT  4.510 2.260 4.790 2.900 ;
        END
    END EB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.100 1.070 2.740 ;
        RECT  0.670 2.100 1.070 2.500 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.260 4.170 2.900 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.350 2.100 1.690 2.500 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.560 -0.380 6.040 0.560 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.640 -0.380 1.040 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.260 3.850 4.660 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  1.020 4.200 1.420 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.620 2.910 2.890 3.310 ;
        RECT  2.620 0.800 2.860 3.310 ;
        RECT  5.250 1.780 5.490 2.660 ;
        RECT  4.440 1.780 5.490 2.020 ;
        RECT  4.440 0.800 4.680 2.020 ;
        RECT  2.620 0.800 4.680 1.040 ;
        RECT  3.410 1.360 3.650 3.310 ;
        RECT  3.410 1.360 3.720 1.760 ;
        RECT  0.240 3.720 3.240 3.960 ;
        RECT  0.240 2.910 0.480 3.960 ;
        RECT  0.190 1.360 0.430 3.310 ;
        RECT  0.240 0.800 0.480 1.760 ;
        RECT  0.240 0.800 2.380 1.040 ;
        RECT  1.930 1.360 2.170 3.310 ;
        RECT  1.760 1.360 2.170 1.760 ;
    END
END MUXB2S

MACRO MUXB2T
    CLASS CORE ;
    FOREIGN MUXB2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.300 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.140 1.290 8.420 1.530 ;
        RECT  7.300 3.220 9.140 3.460 ;
        RECT  7.610 1.290 7.890 3.460 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 2.250 6.030 2.900 ;
        END
    END EB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.100 1.070 2.740 ;
        RECT  0.670 2.100 1.070 2.500 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.250 4.170 2.900 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.350 2.100 1.690 2.500 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.370 -0.380 4.770 0.560 ;
        RECT  5.930 -0.380 6.330 0.560 ;
        RECT  7.230 -0.380 7.630 0.560 ;
        RECT  8.740 -0.380 9.140 1.450 ;
        RECT  0.000 -0.380 9.300 0.380 ;
        RECT  0.640 -0.380 1.040 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.260 4.180 4.660 5.420 ;
        RECT  5.860 4.180 6.260 5.420 ;
        RECT  0.000 4.660 9.300 5.420 ;
        RECT  1.020 4.200 1.420 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.140 3.700 8.420 3.940 ;
        RECT  2.680 2.910 2.930 3.310 ;
        RECT  2.680 0.800 2.920 3.310 ;
        RECT  7.130 1.770 7.370 2.650 ;
        RECT  3.890 1.770 7.370 2.010 ;
        RECT  3.890 0.800 4.130 2.010 ;
        RECT  2.680 1.360 2.930 1.760 ;
        RECT  2.680 0.800 4.130 1.040 ;
        RECT  3.410 1.360 3.650 3.310 ;
        RECT  0.240 3.720 3.240 3.960 ;
        RECT  0.240 2.910 0.480 3.960 ;
        RECT  0.190 1.360 0.430 3.310 ;
        RECT  0.240 0.800 0.480 1.760 ;
        RECT  0.240 0.800 2.380 1.040 ;
        RECT  1.980 0.720 2.380 1.040 ;
        RECT  1.930 1.360 2.170 3.310 ;
    END
END MUXB2T

MACRO MUXB4
    CLASS CORE ;
    FOREIGN MUXB4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.020 2.790 15.330 3.190 ;
        RECT  15.050 0.850 15.330 3.300 ;
        RECT  14.070 0.850 15.330 1.130 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END S0
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 2.100 14.090 2.740 ;
        END
    END EB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.100 8.510 2.740 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 2.100 9.280 2.500 ;
        RECT  8.850 2.100 9.130 2.740 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 2.100 13.470 2.740 ;
        RECT  13.170 2.100 13.470 2.500 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 -0.380 2.600 0.560 ;
        RECT  8.730 -0.380 9.130 0.560 ;
        RECT  13.300 -0.380 13.700 1.130 ;
        RECT  14.940 -0.380 15.340 0.560 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 4.480 2.600 5.420 ;
        RECT  8.730 4.480 9.130 5.420 ;
        RECT  13.510 4.260 13.910 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.960 3.780 14.690 4.020 ;
        RECT  14.450 2.100 14.690 4.020 ;
        RECT  10.960 1.370 11.200 4.020 ;
        RECT  14.450 2.100 14.810 2.500 ;
        RECT  12.400 1.170 12.640 3.310 ;
        RECT  11.680 0.800 11.920 3.310 ;
        RECT  6.690 2.990 7.090 3.230 ;
        RECT  6.770 0.800 7.010 3.230 ;
        RECT  6.770 0.800 11.920 1.040 ;
        RECT  4.610 4.000 10.480 4.240 ;
        RECT  10.240 1.370 10.480 4.240 ;
        RECT  4.610 1.370 4.850 4.240 ;
        RECT  6.050 3.520 9.760 3.760 ;
        RECT  9.520 1.490 9.760 3.760 ;
        RECT  6.050 1.370 6.290 3.760 ;
        RECT  7.560 1.490 7.800 3.190 ;
        RECT  0.830 0.800 1.070 3.380 ;
        RECT  5.330 0.800 5.570 3.310 ;
        RECT  0.830 0.800 5.570 1.040 ;
        RECT  1.550 4.000 4.130 4.240 ;
        RECT  3.890 1.370 4.130 4.240 ;
        RECT  1.550 2.980 1.790 4.240 ;
        RECT  1.530 1.490 1.770 3.220 ;
        RECT  1.530 1.490 1.790 1.890 ;
        RECT  3.170 1.490 3.410 3.190 ;
        RECT  3.170 2.100 3.610 2.500 ;
    END
END MUXB4

MACRO MUXB4P
    CLASS CORE ;
    FOREIGN MUXB4P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 1.570 16.570 3.540 ;
        RECT  15.360 3.300 17.200 3.540 ;
        RECT  13.850 1.570 16.570 1.810 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END S0
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 2.100 14.090 2.740 ;
        END
    END EB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.100 8.510 2.740 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 2.100 9.280 2.500 ;
        RECT  8.850 2.100 9.130 2.740 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 2.100 13.470 2.740 ;
        RECT  12.980 2.100 13.470 2.500 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 -0.380 2.600 0.560 ;
        RECT  8.730 -0.380 9.130 0.560 ;
        RECT  13.060 -0.380 13.460 0.560 ;
        RECT  14.560 -0.380 14.960 0.560 ;
        RECT  15.280 -0.380 15.680 0.560 ;
        RECT  16.800 -0.380 17.200 1.450 ;
        RECT  0.000 -0.380 17.360 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 4.480 2.600 5.420 ;
        RECT  8.730 4.480 9.130 5.420 ;
        RECT  13.100 4.260 13.500 5.420 ;
        RECT  14.540 4.260 14.940 5.420 ;
        RECT  0.000 4.660 17.360 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.820 3.780 16.480 4.020 ;
        RECT  10.960 3.780 13.580 4.020 ;
        RECT  13.340 3.190 13.580 4.020 ;
        RECT  10.960 1.370 11.200 4.020 ;
        RECT  13.340 3.190 15.020 3.430 ;
        RECT  14.780 2.100 15.020 3.430 ;
        RECT  14.780 2.100 15.450 2.500 ;
        RECT  12.210 2.910 12.640 3.310 ;
        RECT  12.210 1.490 12.450 3.310 ;
        RECT  12.210 1.490 12.640 1.890 ;
        RECT  11.680 0.800 11.920 3.310 ;
        RECT  6.690 2.990 7.090 3.230 ;
        RECT  6.770 0.800 7.010 3.230 ;
        RECT  6.770 0.800 11.920 1.040 ;
        RECT  4.610 4.000 10.480 4.240 ;
        RECT  10.240 1.370 10.480 4.240 ;
        RECT  4.610 1.370 4.850 4.240 ;
        RECT  6.050 3.520 9.760 3.760 ;
        RECT  9.520 1.490 9.760 3.760 ;
        RECT  6.050 1.370 6.290 3.760 ;
        RECT  7.560 1.490 7.800 3.190 ;
        RECT  0.830 0.800 1.070 3.380 ;
        RECT  5.330 0.800 5.570 3.310 ;
        RECT  0.830 0.800 5.570 1.040 ;
        RECT  1.550 4.000 4.130 4.240 ;
        RECT  3.890 1.370 4.130 4.240 ;
        RECT  1.550 2.980 1.790 4.240 ;
        RECT  1.530 1.490 1.770 3.220 ;
        RECT  1.530 1.490 1.790 1.890 ;
        RECT  3.170 1.490 3.410 3.190 ;
        RECT  3.170 2.100 3.610 2.500 ;
    END
END MUXB4P

MACRO MUXB4S
    CLASS CORE ;
    FOREIGN MUXB4S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.020 2.790 15.330 3.190 ;
        RECT  15.050 1.050 15.330 3.300 ;
        RECT  14.070 1.050 15.330 1.330 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END S0
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 2.100 14.090 2.740 ;
        END
    END EB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.100 8.510 2.740 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 2.100 9.280 2.500 ;
        RECT  8.850 2.100 9.130 2.740 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 2.100 13.470 2.740 ;
        RECT  13.170 2.100 13.470 2.500 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 -0.380 2.600 0.560 ;
        RECT  8.730 -0.380 9.130 0.560 ;
        RECT  13.300 -0.380 13.700 1.330 ;
        RECT  14.940 -0.380 15.340 0.560 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 4.480 2.600 5.420 ;
        RECT  8.730 4.480 9.130 5.420 ;
        RECT  13.510 3.730 13.910 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.960 3.550 13.120 3.790 ;
        RECT  12.880 2.980 13.120 3.790 ;
        RECT  10.960 1.370 11.200 3.790 ;
        RECT  12.880 2.980 14.690 3.220 ;
        RECT  14.450 2.100 14.690 3.220 ;
        RECT  14.450 2.100 14.810 2.500 ;
        RECT  12.400 1.170 12.640 3.310 ;
        RECT  11.680 0.800 11.920 3.310 ;
        RECT  6.690 2.990 7.090 3.230 ;
        RECT  6.770 0.800 7.010 3.230 ;
        RECT  6.770 0.800 11.920 1.040 ;
        RECT  4.610 4.000 10.480 4.240 ;
        RECT  10.240 1.370 10.480 4.240 ;
        RECT  4.610 1.370 4.850 4.240 ;
        RECT  6.050 3.520 9.760 3.760 ;
        RECT  9.520 1.490 9.760 3.760 ;
        RECT  6.050 1.370 6.290 3.760 ;
        RECT  7.560 1.490 7.800 3.190 ;
        RECT  0.830 0.800 1.070 3.380 ;
        RECT  5.330 0.800 5.570 3.310 ;
        RECT  0.830 0.800 5.570 1.040 ;
        RECT  1.550 4.000 4.130 4.240 ;
        RECT  3.890 1.370 4.130 4.240 ;
        RECT  1.550 2.980 1.790 4.240 ;
        RECT  1.530 1.490 1.770 3.220 ;
        RECT  1.530 1.490 1.790 1.890 ;
        RECT  3.170 1.490 3.410 3.190 ;
        RECT  3.170 2.100 3.610 2.500 ;
    END
END MUXB4S

MACRO MUXB4T
    CLASS CORE ;
    FOREIGN MUXB4T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.980 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.910 1.570 17.190 3.540 ;
        RECT  15.980 3.300 17.820 3.540 ;
        RECT  13.850 1.570 17.190 1.810 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END S0
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 2.100 14.090 2.740 ;
        END
    END EB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.100 8.510 2.740 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 2.100 9.280 2.500 ;
        RECT  8.850 2.100 9.130 2.740 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 2.100 13.470 2.740 ;
        RECT  12.980 2.100 13.470 2.500 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 -0.380 2.600 0.560 ;
        RECT  8.730 -0.380 9.130 0.560 ;
        RECT  13.060 -0.380 13.460 0.560 ;
        RECT  14.640 -0.380 15.040 0.560 ;
        RECT  15.910 -0.380 16.310 0.560 ;
        RECT  17.420 -0.380 17.820 1.450 ;
        RECT  0.000 -0.380 17.980 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 4.480 2.600 5.420 ;
        RECT  8.730 4.480 9.130 5.420 ;
        RECT  13.100 4.260 13.500 5.420 ;
        RECT  14.540 4.260 14.940 5.420 ;
        RECT  0.000 4.660 17.980 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.820 3.780 17.100 4.020 ;
        RECT  10.960 3.780 13.580 4.020 ;
        RECT  13.340 3.190 13.580 4.020 ;
        RECT  10.960 1.370 11.200 4.020 ;
        RECT  13.340 3.190 15.740 3.430 ;
        RECT  15.500 2.100 15.740 3.430 ;
        RECT  15.500 2.100 16.070 2.500 ;
        RECT  12.210 2.910 12.640 3.310 ;
        RECT  12.210 1.490 12.450 3.310 ;
        RECT  12.210 1.490 12.640 1.890 ;
        RECT  11.680 0.800 11.920 3.310 ;
        RECT  6.690 2.990 7.090 3.230 ;
        RECT  6.770 0.800 7.010 3.230 ;
        RECT  6.770 0.800 11.920 1.040 ;
        RECT  4.610 4.000 10.480 4.240 ;
        RECT  10.240 1.370 10.480 4.240 ;
        RECT  4.610 1.370 4.850 4.240 ;
        RECT  6.050 3.520 9.760 3.760 ;
        RECT  9.520 1.490 9.760 3.760 ;
        RECT  6.050 1.370 6.290 3.760 ;
        RECT  7.560 1.490 7.800 3.190 ;
        RECT  0.830 0.800 1.070 3.380 ;
        RECT  5.330 0.800 5.570 3.310 ;
        RECT  0.830 0.800 5.570 1.040 ;
        RECT  1.550 4.000 4.130 4.240 ;
        RECT  3.890 1.370 4.130 4.240 ;
        RECT  1.550 2.980 1.790 4.240 ;
        RECT  1.530 1.490 1.770 3.220 ;
        RECT  1.530 1.490 1.790 1.890 ;
        RECT  3.170 1.490 3.410 3.190 ;
        RECT  3.170 2.100 3.610 2.500 ;
    END
END MUXB4T

MACRO MXL2H
    CLASS CORE ;
    FOREIGN MXL2H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.730 1.100 4.970 1.720 ;
        RECT  4.730 1.480 6.650 1.720 ;
        RECT  6.370 1.480 6.650 3.460 ;
        RECT  3.280 3.220 6.650 3.460 ;
        RECT  3.210 1.100 4.970 1.340 ;
        END
    END OB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.170 2.360 2.570 ;
        RECT  2.030 2.170 2.310 2.790 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.150 0.690 2.550 ;
        RECT  0.170 2.150 0.450 2.790 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.250 8.510 2.890 ;
        RECT  7.990 2.250 8.510 2.650 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 -0.380 2.070 0.770 ;
        RECT  6.610 -0.380 7.010 0.760 ;
        RECT  8.120 -0.380 8.520 0.950 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 4.480 2.170 5.420 ;
        RECT  6.680 4.260 7.080 5.420 ;
        RECT  8.120 4.260 8.520 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.000 3.700 7.720 3.940 ;
        RECT  7.480 1.000 7.720 3.940 ;
        RECT  5.370 1.000 7.720 1.240 ;
        RECT  2.620 4.180 5.840 4.420 ;
        RECT  0.960 4.000 2.860 4.240 ;
        RECT  0.960 1.010 1.200 4.240 ;
        RECT  0.960 1.010 2.550 1.250 ;
        RECT  2.310 0.620 2.550 1.250 ;
        RECT  2.310 0.620 4.330 0.860 ;
        RECT  2.640 1.490 2.880 3.190 ;
        RECT  2.640 2.330 5.310 2.570 ;
        RECT  2.570 1.490 2.880 1.890 ;
    END
END MXL2H

MACRO MXL2HF
    CLASS CORE ;
    FOREIGN MXL2HF 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 28.520 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.440 2.870 10.680 3.460 ;
        RECT  21.270 1.570 21.510 3.460 ;
        RECT  10.440 3.220 21.640 3.460 ;
        RECT  9.840 1.570 21.760 1.810 ;
        RECT  9.720 2.870 10.680 3.110 ;
        END
    END OB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.170 6.650 2.810 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.150 3.550 2.790 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  25.590 2.250 25.870 2.890 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  5.990 -0.380 6.390 0.850 ;
        RECT  7.710 -0.380 8.110 0.850 ;
        RECT  9.330 -0.380 9.730 0.850 ;
        RECT  22.200 -0.380 22.600 0.870 ;
        RECT  23.640 -0.380 24.040 0.850 ;
        RECT  25.080 -0.380 25.480 0.850 ;
        RECT  26.520 -0.380 26.920 0.850 ;
        RECT  27.960 -0.380 28.360 0.850 ;
        RECT  0.000 -0.380 28.520 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  5.930 4.260 6.330 5.420 ;
        RECT  7.580 3.930 7.980 5.420 ;
        RECT  9.180 3.930 9.580 5.420 ;
        RECT  22.200 4.190 22.600 5.420 ;
        RECT  23.640 4.260 24.040 5.420 ;
        RECT  25.080 4.260 25.480 5.420 ;
        RECT  26.520 4.260 26.920 5.420 ;
        RECT  27.960 4.260 28.360 5.420 ;
        RECT  0.000 4.660 28.520 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.440 3.700 27.640 3.940 ;
        RECT  23.000 3.660 27.640 3.940 ;
        RECT  23.000 1.110 23.240 3.940 ;
        RECT  23.000 1.390 27.640 1.670 ;
        RECT  21.860 1.110 23.240 1.350 ;
        RECT  16.320 1.090 22.100 1.330 ;
        RECT  9.960 4.180 20.920 4.420 ;
        RECT  9.960 3.420 10.200 4.420 ;
        RECT  0.880 3.420 10.200 3.660 ;
        RECT  5.280 1.090 5.520 3.660 ;
        RECT  0.880 1.210 5.520 1.450 ;
        RECT  10.560 0.710 10.800 1.330 ;
        RECT  5.280 1.090 10.800 1.330 ;
        RECT  10.560 0.710 15.280 0.950 ;
        RECT  6.860 2.940 8.860 3.180 ;
        RECT  8.540 1.570 8.780 3.180 ;
        RECT  8.540 2.330 16.690 2.570 ;
        RECT  6.890 1.570 8.940 1.810 ;
    END
END MXL2HF

MACRO MXL2HP
    CLASS CORE ;
    FOREIGN MXL2HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.340 3.220 11.500 3.460 ;
        RECT  5.290 1.570 11.530 1.810 ;
        RECT  10.090 1.570 10.370 3.460 ;
        END
    END OB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.170 3.790 2.570 ;
        RECT  3.270 2.170 3.550 2.810 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.150 1.690 2.810 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 2.250 14.090 2.910 ;
        RECT  13.690 2.250 14.090 2.650 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.110 -0.380 3.510 0.850 ;
        RECT  4.840 -0.380 5.240 0.850 ;
        RECT  11.990 -0.380 12.390 0.870 ;
        RECT  13.500 -0.380 13.900 0.950 ;
        RECT  14.940 -0.380 15.340 0.950 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.050 4.260 3.450 5.420 ;
        RECT  4.790 4.180 5.190 5.420 ;
        RECT  12.060 4.190 12.460 5.420 ;
        RECT  13.500 4.260 13.900 5.420 ;
        RECT  14.940 4.260 15.340 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.060 3.700 14.620 3.940 ;
        RECT  12.860 3.660 14.620 3.940 ;
        RECT  12.860 1.110 13.100 3.940 ;
        RECT  12.860 1.190 14.620 1.470 ;
        RECT  11.650 1.110 13.100 1.350 ;
        RECT  8.890 1.090 11.890 1.330 ;
        RECT  5.580 4.180 10.780 4.420 ;
        RECT  5.580 3.700 5.820 4.420 ;
        RECT  0.880 3.700 5.820 3.940 ;
        RECT  2.400 1.090 2.640 3.940 ;
        RECT  0.880 1.190 2.640 1.470 ;
        RECT  2.400 1.090 7.930 1.330 ;
        RECT  4.080 1.570 4.320 3.190 ;
        RECT  4.080 2.330 9.480 2.570 ;
        RECT  3.930 1.570 4.330 1.810 ;
    END
END MXL2HP

MACRO MXL2HS
    CLASS CORE ;
    FOREIGN MXL2HS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.910 1.480 4.150 3.110 ;
        RECT  2.860 2.870 4.150 3.110 ;
        RECT  2.880 1.480 4.150 1.720 ;
        END
    END OB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.170 1.720 2.570 ;
        RECT  1.410 2.170 1.690 2.790 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.150 1.070 2.790 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.250 4.790 2.890 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.230 -0.380 4.630 0.560 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.950 -0.380 1.350 0.840 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.120 4.480 4.520 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.930 4.130 1.330 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.140 4.000 2.540 4.320 ;
        RECT  2.140 4.000 5.340 4.240 ;
        RECT  5.100 1.000 5.340 4.240 ;
        RECT  3.600 1.000 5.340 1.240 ;
        RECT  0.240 3.510 3.980 3.750 ;
        RECT  0.240 1.080 0.480 3.750 ;
        RECT  0.240 1.080 1.830 1.320 ;
        RECT  1.590 0.620 1.830 1.320 ;
        RECT  1.590 0.620 2.560 0.860 ;
        RECT  1.630 3.030 2.340 3.270 ;
        RECT  2.100 1.560 2.340 3.270 ;
        RECT  2.100 2.330 3.470 2.570 ;
        RECT  1.630 1.560 2.340 1.800 ;
    END
END MXL2HS

MACRO MXL2HT
    CLASS CORE ;
    FOREIGN MXL2HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.700 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 1.570 16.570 3.460 ;
        RECT  7.670 1.570 16.710 1.810 ;
        RECT  7.750 3.220 16.710 3.460 ;
        RECT  7.750 3.220 7.990 3.890 ;
        END
    END OB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.170 5.030 2.570 ;
        RECT  4.510 2.170 4.790 2.810 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.310 2.840 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  19.390 2.250 19.670 2.890 ;
        RECT  19.270 2.250 19.670 2.650 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.550 -0.380 4.950 0.850 ;
        RECT  6.160 -0.380 6.560 0.850 ;
        RECT  16.820 -0.380 17.220 0.780 ;
        RECT  18.260 -0.380 18.660 0.780 ;
        RECT  19.700 -0.380 20.100 0.780 ;
        RECT  21.140 -0.380 21.540 0.780 ;
        RECT  0.000 -0.380 21.700 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  6.160 3.930 6.560 5.420 ;
        RECT  16.820 4.260 17.220 5.420 ;
        RECT  18.260 4.260 18.660 5.420 ;
        RECT  19.700 4.260 20.100 5.420 ;
        RECT  21.140 4.260 21.540 5.420 ;
        RECT  0.000 4.660 21.700 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.390 3.700 20.820 3.940 ;
        RECT  17.620 1.040 17.860 3.940 ;
        RECT  12.710 1.040 20.820 1.280 ;
        RECT  7.270 4.180 15.990 4.420 ;
        RECT  7.270 3.430 7.510 4.420 ;
        RECT  0.880 3.430 7.510 3.670 ;
        RECT  3.840 1.090 4.080 3.670 ;
        RECT  0.880 1.210 4.080 1.450 ;
        RECT  7.200 0.710 7.440 1.330 ;
        RECT  3.840 1.090 7.440 1.330 ;
        RECT  7.200 0.710 11.670 0.950 ;
        RECT  5.440 2.870 7.420 3.110 ;
        RECT  7.100 1.570 7.340 3.110 ;
        RECT  7.100 2.330 13.100 2.570 ;
        RECT  5.340 1.570 7.370 1.810 ;
    END
END MXL2HT

MACRO MXL3
    CLASS CORE ;
    FOREIGN MXL3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.880 1.090 4.160 ;
        RECT  0.750 3.920 1.150 4.420 ;
        RECT  0.170 3.420 0.450 4.160 ;
        END
    END S0
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.220 8.510 3.310 ;
        RECT  8.200 2.910 8.510 3.310 ;
        RECT  8.200 1.490 8.510 1.890 ;
        END
    END OB
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.350 2.130 6.670 2.740 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.160 0.480 2.560 ;
        RECT  0.170 1.980 0.450 2.620 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 3.750 2.960 4.150 ;
        RECT  2.650 3.500 2.930 4.420 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.100 3.730 2.500 ;
        RECT  3.270 2.100 3.550 2.850 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.470 -0.380 3.870 0.860 ;
        RECT  6.240 0.630 6.720 1.030 ;
        RECT  6.440 -0.380 6.720 1.890 ;
        RECT  6.440 1.490 6.780 1.890 ;
        RECT  7.650 -0.380 7.960 1.100 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  0.500 -0.380 0.900 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 4.160 4.010 5.420 ;
        RECT  5.640 4.480 6.040 5.420 ;
        RECT  6.360 2.980 6.620 5.420 ;
        RECT  6.360 2.980 6.760 3.220 ;
        RECT  7.580 4.160 7.990 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.140 4.400 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.860 3.680 7.100 4.370 ;
        RECT  6.860 3.680 7.870 3.920 ;
        RECT  7.630 1.340 7.870 3.920 ;
        RECT  7.090 1.340 7.870 1.580 ;
        RECT  7.090 0.630 7.330 1.580 ;
        RECT  6.960 0.630 7.330 1.030 ;
        RECT  5.650 0.620 5.890 3.190 ;
        RECT  5.650 1.490 6.060 1.890 ;
        RECT  5.020 0.620 5.890 0.860 ;
        RECT  5.050 3.770 6.040 4.010 ;
        RECT  5.050 2.950 5.290 4.010 ;
        RECT  4.930 1.480 5.170 3.190 ;
        RECT  4.450 4.180 4.870 4.420 ;
        RECT  4.450 0.620 4.690 4.420 ;
        RECT  4.190 0.620 4.690 0.860 ;
        RECT  3.970 1.100 4.210 3.570 ;
        RECT  1.810 1.100 2.050 3.200 ;
        RECT  1.810 1.100 4.210 1.340 ;
        RECT  2.460 2.880 2.860 3.120 ;
        RECT  2.540 1.580 2.780 3.120 ;
        RECT  2.450 1.580 2.850 1.820 ;
        RECT  1.390 4.170 1.790 4.410 ;
        RECT  1.390 3.490 1.630 4.410 ;
        RECT  1.330 0.620 1.570 3.740 ;
        RECT  1.330 0.620 2.550 0.860 ;
        RECT  0.840 1.490 1.080 3.200 ;
    END
END MXL3

MACRO MXL3P
    CLASS CORE ;
    FOREIGN MXL3P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.880 1.090 4.160 ;
        RECT  0.750 3.920 1.150 4.420 ;
        RECT  0.170 3.410 0.450 4.160 ;
        END
    END S0
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 1.490 9.130 3.190 ;
        RECT  8.720 2.790 9.130 3.190 ;
        RECT  8.720 1.490 9.130 1.890 ;
        END
    END OB
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.350 2.130 6.670 2.740 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.160 0.480 2.560 ;
        RECT  0.170 1.980 0.450 2.620 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 3.750 2.960 4.150 ;
        RECT  2.650 3.480 2.930 4.420 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.200 3.730 2.600 ;
        RECT  3.270 2.200 3.550 2.850 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.470 -0.380 3.870 0.860 ;
        RECT  6.520 -0.380 6.800 1.890 ;
        RECT  7.930 -0.380 8.310 1.030 ;
        RECT  9.370 -0.380 9.750 1.030 ;
        RECT  0.000 -0.380 9.920 0.380 ;
        RECT  0.500 -0.380 0.900 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 4.170 4.010 5.420 ;
        RECT  5.640 4.480 6.040 5.420 ;
        RECT  6.360 3.090 6.760 5.420 ;
        RECT  7.920 4.180 8.330 5.420 ;
        RECT  9.350 4.180 9.760 5.420 ;
        RECT  0.000 4.660 9.920 5.420 ;
        RECT  0.160 4.400 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.260 1.490 7.500 3.190 ;
        RECT  7.260 2.300 8.450 2.540 ;
        RECT  5.650 0.620 5.890 3.190 ;
        RECT  5.650 1.490 6.060 1.890 ;
        RECT  5.020 0.620 5.890 0.860 ;
        RECT  5.050 3.770 6.040 4.010 ;
        RECT  5.050 2.950 5.290 4.010 ;
        RECT  4.930 1.480 5.170 3.190 ;
        RECT  4.450 4.180 4.870 4.420 ;
        RECT  4.450 0.620 4.690 4.420 ;
        RECT  4.190 0.620 4.690 0.860 ;
        RECT  3.970 1.100 4.210 3.570 ;
        RECT  1.810 1.100 2.050 3.200 ;
        RECT  1.810 1.100 4.210 1.340 ;
        RECT  2.460 2.880 2.860 3.120 ;
        RECT  2.540 1.580 2.780 3.120 ;
        RECT  2.450 1.580 2.850 1.820 ;
        RECT  1.390 4.170 1.790 4.410 ;
        RECT  1.390 3.500 1.630 4.410 ;
        RECT  1.330 0.620 1.570 3.740 ;
        RECT  1.330 0.620 2.550 0.860 ;
        RECT  0.840 1.490 1.080 3.200 ;
    END
END MXL3P

MACRO MXL3S
    CLASS CORE ;
    FOREIGN MXL3S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.880 1.090 4.160 ;
        RECT  0.750 3.920 1.150 4.420 ;
        RECT  0.170 3.420 0.450 4.160 ;
        END
    END S0
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 0.770 8.510 4.100 ;
        RECT  8.200 3.700 8.510 4.100 ;
        RECT  8.200 0.770 8.510 1.170 ;
        END
    END OB
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.350 2.130 6.670 2.740 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.160 0.480 2.560 ;
        RECT  0.170 1.980 0.450 2.620 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 3.750 2.960 4.150 ;
        RECT  2.650 3.500 2.930 4.420 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.200 3.730 2.600 ;
        RECT  3.270 2.200 3.550 2.850 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.470 -0.380 3.870 0.860 ;
        RECT  6.520 -0.380 6.800 1.890 ;
        RECT  7.410 -0.380 7.720 1.170 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  0.500 -0.380 0.900 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 4.170 4.010 5.420 ;
        RECT  5.640 4.480 6.040 5.420 ;
        RECT  6.360 3.090 6.760 5.420 ;
        RECT  7.400 4.180 7.810 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.140 4.400 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.350 1.490 7.590 3.190 ;
        RECT  7.350 2.300 7.930 2.540 ;
        RECT  5.650 0.620 5.890 3.190 ;
        RECT  5.650 1.490 6.060 1.890 ;
        RECT  5.020 0.620 5.890 0.860 ;
        RECT  5.050 3.770 6.040 4.010 ;
        RECT  5.050 2.950 5.290 4.010 ;
        RECT  4.930 1.480 5.170 3.190 ;
        RECT  4.450 4.180 4.870 4.420 ;
        RECT  4.450 0.620 4.690 4.420 ;
        RECT  4.190 0.620 4.690 0.860 ;
        RECT  3.970 1.100 4.210 3.570 ;
        RECT  1.810 1.100 2.050 3.200 ;
        RECT  1.810 1.100 4.210 1.340 ;
        RECT  2.460 2.880 2.860 3.120 ;
        RECT  2.540 1.580 2.780 3.120 ;
        RECT  2.450 1.580 2.850 1.820 ;
        RECT  1.390 4.170 1.790 4.410 ;
        RECT  1.390 3.500 1.630 4.410 ;
        RECT  1.330 0.620 1.570 3.740 ;
        RECT  1.330 0.620 2.550 0.860 ;
        RECT  0.840 1.490 1.080 3.200 ;
    END
END MXL3S

MACRO MXL3T
    CLASS CORE ;
    FOREIGN MXL3T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.540 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.880 1.090 4.160 ;
        RECT  0.750 3.920 1.150 4.420 ;
        RECT  0.170 3.420 0.450 4.160 ;
        END
    END S0
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.540 1.570 10.380 1.810 ;
        RECT  8.540 2.870 10.380 3.110 ;
        RECT  9.470 1.570 9.750 3.110 ;
        END
    END OB
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.350 2.130 6.670 2.740 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.160 0.480 2.560 ;
        RECT  0.170 1.980 0.450 2.620 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.640 3.830 3.040 4.070 ;
        RECT  2.650 3.500 2.930 4.420 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.200 3.730 2.600 ;
        RECT  3.270 2.200 3.550 2.850 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.470 -0.380 3.870 0.860 ;
        RECT  6.520 -0.380 6.800 1.890 ;
        RECT  7.830 -0.380 8.210 1.030 ;
        RECT  9.270 -0.380 9.650 1.030 ;
        RECT  0.000 -0.380 10.540 0.380 ;
        RECT  0.500 -0.380 0.900 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 4.170 4.010 5.420 ;
        RECT  5.640 4.480 6.040 5.420 ;
        RECT  6.360 3.090 6.760 5.420 ;
        RECT  7.820 4.180 8.230 5.420 ;
        RECT  9.250 4.180 9.660 5.420 ;
        RECT  0.000 4.660 10.540 5.420 ;
        RECT  0.140 4.400 0.480 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.260 1.490 7.500 3.190 ;
        RECT  7.260 2.300 8.350 2.540 ;
        RECT  5.650 0.620 5.890 3.190 ;
        RECT  5.650 1.490 6.060 1.890 ;
        RECT  5.020 0.620 5.890 0.860 ;
        RECT  5.050 3.770 6.040 4.010 ;
        RECT  5.050 2.950 5.290 4.010 ;
        RECT  4.930 1.480 5.170 3.190 ;
        RECT  4.450 4.180 4.870 4.420 ;
        RECT  4.450 0.620 4.690 4.420 ;
        RECT  4.190 0.620 4.690 0.860 ;
        RECT  3.970 1.100 4.210 3.570 ;
        RECT  1.810 1.100 2.050 3.200 ;
        RECT  1.810 1.100 4.210 1.340 ;
        RECT  2.460 2.880 2.860 3.120 ;
        RECT  2.460 1.580 2.700 3.120 ;
        RECT  2.460 1.580 2.860 1.820 ;
        RECT  1.390 4.170 1.790 4.410 ;
        RECT  1.390 3.500 1.630 4.410 ;
        RECT  1.330 0.620 1.570 3.740 ;
        RECT  1.330 0.620 2.550 0.860 ;
        RECT  0.840 1.490 1.080 3.200 ;
    END
END MXL3T

MACRO ND2
    CLASS CORE ;
    FOREIGN ND2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.860 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.260 1.070 3.300 ;
        RECT  0.160 1.260 1.070 1.540 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.200 1.690 2.840 ;
        RECT  1.350 2.250 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.550 2.650 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.860 0.380 ;
        RECT  1.300 -0.380 1.700 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 4.480 1.700 5.420 ;
        RECT  0.000 4.660 1.860 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
END ND2

MACRO ND2F
    CLASS CORE ;
    FOREIGN ND2F 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 3.070 4.170 3.780 ;
        RECT  0.160 3.500 4.170 3.780 ;
        RECT  1.410 1.260 5.410 1.540 ;
        RECT  5.130 1.260 5.410 3.350 ;
        RECT  3.890 3.070 6.050 3.350 ;
        RECT  1.550 1.260 1.950 1.650 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.030 1.070 3.220 ;
        RECT  3.130 2.460 3.410 3.220 ;
        RECT  0.790 2.940 3.410 3.220 ;
        RECT  0.690 2.030 1.070 2.430 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.160 1.820 4.170 2.100 ;
        RECT  3.890 1.820 4.170 2.740 ;
        RECT  1.640 2.090 2.440 2.370 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.730 -0.380 3.130 0.870 ;
        RECT  5.460 -0.380 5.860 0.870 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.160 -0.380 0.560 0.840 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 4.260 2.640 5.420 ;
        RECT  3.550 4.260 3.950 5.420 ;
        RECT  4.940 3.890 5.340 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.860 4.260 1.260 5.420 ;
        END
    END VCC
END ND2F

MACRO ND2P
    CLASS CORE ;
    FOREIGN ND2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.450 1.200 2.930 1.600 ;
        RECT  2.400 3.480 2.930 3.760 ;
        RECT  0.790 3.520 2.930 3.760 ;
        RECT  2.650 1.200 2.930 3.860 ;
        RECT  0.970 3.380 1.370 3.760 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.110 1.070 2.840 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.110 2.350 2.510 ;
        RECT  2.030 2.110 2.310 2.840 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  1.040 -0.380 1.440 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.640 4.480 2.040 5.420 ;
        RECT  3.160 4.480 3.560 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 1.430 2.050 1.670 ;
        RECT  1.810 0.720 2.050 1.670 ;
        RECT  1.810 0.720 3.490 0.960 ;
    END
END ND2P

MACRO ND2S
    CLASS CORE ;
    FOREIGN ND2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.860 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.260 1.070 3.280 ;
        RECT  0.160 1.260 1.070 1.540 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.200 1.690 2.840 ;
        RECT  1.350 2.250 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.550 2.650 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.860 0.380 ;
        RECT  1.300 -0.380 1.700 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.290 4.230 1.690 5.420 ;
        RECT  0.000 4.660 1.860 5.420 ;
        RECT  0.160 4.230 0.560 5.420 ;
        END
    END VCC
END ND2S

MACRO ND2T
    CLASS CORE ;
    FOREIGN ND2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.710 3.500 3.940 3.780 ;
        RECT  4.280 1.280 4.790 1.580 ;
        RECT  1.410 1.340 4.790 1.580 ;
        RECT  3.660 3.350 4.790 3.630 ;
        RECT  4.510 1.180 4.790 3.630 ;
        RECT  1.410 1.190 1.730 1.840 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.460 2.930 3.220 ;
        RECT  0.170 2.940 2.930 3.220 ;
        RECT  2.650 2.460 3.170 2.860 ;
        RECT  0.170 2.030 1.070 3.220 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.820 4.170 2.100 ;
        RECT  3.890 1.820 4.170 2.740 ;
        RECT  1.640 2.100 2.310 2.340 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.830 -0.380 3.230 1.100 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.620 4.260 2.020 5.420 ;
        RECT  2.930 4.260 3.330 5.420 ;
        RECT  4.320 3.930 4.720 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.240 4.260 0.640 5.420 ;
        END
    END VCC
END ND2T

MACRO ND3
    CLASS CORE ;
    FOREIGN ND3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 0.890 1.690 1.950 ;
        RECT  1.410 0.890 2.320 1.130 ;
        RECT  0.670 3.040 2.320 3.280 ;
        RECT  1.430 0.890 1.670 3.280 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.220 1.180 2.620 ;
        RECT  0.790 2.200 1.070 2.800 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.200 2.310 2.800 ;
        RECT  1.950 2.250 2.310 2.650 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.490 2.650 ;
        RECT  0.170 2.200 0.450 2.800 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.520 4.480 1.920 5.420 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
END ND3

MACRO ND3HT
    CLASS CORE ;
    FOREIGN ND3HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.440 1.190 7.280 1.430 ;
        RECT  0.880 3.430 7.280 3.670 ;
        RECT  6.390 1.190 6.630 3.670 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.040 4.170 2.810 ;
        RECT  3.870 2.060 4.170 2.460 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.720 2.040 6.060 2.810 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 2.060 1.730 2.460 ;
        RECT  1.400 2.060 1.700 2.860 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 -0.380 2.240 1.110 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 3.910 2.240 5.420 ;
        RECT  3.280 3.910 3.680 5.420 ;
        RECT  4.720 3.910 5.120 5.420 ;
        RECT  6.160 3.910 6.560 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.160 3.910 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.280 0.710 6.560 0.950 ;
        RECT  0.880 1.350 4.400 1.590 ;
    END
END ND3HT

MACRO ND3P
    CLASS CORE ;
    FOREIGN ND3P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.150 4.790 3.960 ;
        RECT  0.850 3.720 4.790 3.960 ;
        RECT  2.140 1.150 4.790 1.390 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.250 3.550 3.480 ;
        RECT  1.410 3.240 3.550 3.480 ;
        RECT  1.410 2.250 1.690 3.480 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.450 2.740 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.630 4.170 2.840 ;
        RECT  0.530 1.630 4.180 1.870 ;
        RECT  3.890 1.820 4.270 2.220 ;
        RECT  0.530 1.630 0.770 2.210 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.260 -0.380 4.660 0.910 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.300 -0.380 0.700 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.440 4.480 1.840 5.420 ;
        RECT  2.900 4.480 3.300 5.420 ;
        RECT  4.400 4.480 4.800 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
END ND3P

MACRO ND3S
    CLASS CORE ;
    FOREIGN ND3S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.500 1.250 1.740 3.460 ;
        RECT  1.410 1.250 2.320 1.550 ;
        RECT  0.670 3.220 2.320 3.460 ;
        RECT  1.410 1.050 1.690 1.990 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.220 1.260 2.620 ;
        RECT  0.790 2.200 1.070 2.800 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.200 2.310 2.800 ;
        RECT  1.980 2.250 2.310 2.650 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.550 2.650 ;
        RECT  0.170 2.200 0.450 2.800 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 4.480 2.100 5.420 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
END ND3S

MACRO ND4
    CLASS CORE ;
    FOREIGN ND4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.720 2.930 6.030 3.330 ;
        RECT  5.750 1.180 6.030 3.860 ;
        RECT  5.720 1.350 6.030 1.750 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.800 1.850 2.200 ;
        RECT  1.410 1.560 1.690 2.200 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        RECT  2.590 2.100 2.930 2.500 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.300 1.070 2.940 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.560 0.500 1.960 ;
        RECT  0.170 1.560 0.450 2.200 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.550 -0.380 3.950 0.560 ;
        RECT  5.060 -0.380 5.460 0.900 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  1.250 -0.380 1.650 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.900 4.480 3.300 5.420 ;
        RECT  4.870 4.260 5.270 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.160 4.480 1.740 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.230 3.270 4.710 3.670 ;
        RECT  4.470 0.660 4.710 3.670 ;
        RECT  4.470 2.380 5.410 2.620 ;
        RECT  4.340 0.660 4.740 0.900 ;
        RECT  2.130 3.720 3.990 3.960 ;
        RECT  3.750 0.870 3.990 3.960 ;
        RECT  3.750 2.290 4.230 2.690 ;
        RECT  2.790 0.870 3.990 1.110 ;
        RECT  0.750 3.720 1.890 3.960 ;
        RECT  1.650 3.240 1.890 3.960 ;
        RECT  1.650 3.240 3.510 3.480 ;
        RECT  3.270 1.350 3.510 3.480 ;
        RECT  2.050 1.350 3.510 1.590 ;
        RECT  2.050 1.080 2.290 1.590 ;
        RECT  0.160 1.080 2.290 1.320 ;
    END
END ND4

MACRO ND4P
    CLASS CORE ;
    FOREIGN ND4P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 1.260 6.650 3.220 ;
        RECT  5.540 2.940 6.650 3.220 ;
        RECT  5.640 1.260 6.650 1.670 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.850 2.500 ;
        RECT  1.410 2.100 1.690 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        RECT  2.630 2.100 2.930 2.500 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.300 1.070 2.940 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.700 0.490 2.100 ;
        RECT  0.170 1.560 0.450 2.200 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.400 -0.380 3.800 0.560 ;
        RECT  5.050 -0.380 5.370 0.980 ;
        RECT  6.230 -0.380 6.630 0.900 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  1.210 -0.380 1.610 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.920 4.260 3.320 5.420 ;
        RECT  4.870 4.260 5.270 5.420 ;
        RECT  6.210 4.260 6.610 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  0.160 4.480 1.740 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.350 2.790 4.750 3.190 ;
        RECT  4.510 0.840 4.750 3.190 ;
        RECT  4.510 2.380 6.120 2.620 ;
        RECT  4.270 0.840 4.750 1.240 ;
        RECT  2.130 3.780 4.030 4.020 ;
        RECT  3.790 0.800 4.030 4.020 ;
        RECT  3.790 2.040 4.270 2.440 ;
        RECT  2.680 0.800 4.030 1.040 ;
        RECT  0.750 3.650 1.890 3.890 ;
        RECT  1.650 3.300 1.890 3.890 ;
        RECT  1.650 3.300 3.550 3.540 ;
        RECT  3.310 1.280 3.550 3.540 ;
        RECT  1.910 1.280 3.550 1.520 ;
        RECT  0.160 1.080 2.150 1.320 ;
    END
END ND4P

MACRO ND4S
    CLASS CORE ;
    FOREIGN ND4S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.720 3.340 6.030 3.740 ;
        RECT  5.750 0.880 6.030 3.860 ;
        RECT  5.720 1.030 6.030 1.430 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  1.940 2.100 2.310 2.500 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 2.930 2.740 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.100 1.070 2.740 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.540 0.500 1.940 ;
        RECT  0.170 1.540 0.450 2.180 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.530 -0.380 3.930 0.560 ;
        RECT  4.850 -0.380 5.250 0.560 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  1.480 -0.380 1.880 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.490 4.480 1.890 5.420 ;
        RECT  3.210 4.480 3.610 5.420 ;
        RECT  4.910 4.480 5.310 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.410 3.410 4.840 3.810 ;
        RECT  4.600 1.190 4.840 3.810 ;
        RECT  4.600 2.790 5.410 3.030 ;
        RECT  4.270 1.190 4.840 1.430 ;
        RECT  4.270 1.030 4.510 1.430 ;
        RECT  2.350 4.000 4.170 4.240 ;
        RECT  3.930 1.840 4.170 4.240 ;
        RECT  3.930 2.770 4.360 3.170 ;
        RECT  3.790 0.890 4.030 2.080 ;
        RECT  2.810 0.890 4.030 1.130 ;
        RECT  0.820 3.740 2.110 3.980 ;
        RECT  3.310 1.370 3.550 3.760 ;
        RECT  1.870 3.520 3.550 3.760 ;
        RECT  0.820 3.650 1.220 3.980 ;
        RECT  3.310 2.870 3.660 3.270 ;
        RECT  2.330 1.370 3.550 1.610 ;
        RECT  2.330 0.890 2.570 1.610 ;
        RECT  0.160 0.890 2.570 1.130 ;
    END
END ND4S

MACRO ND4T
    CLASS CORE ;
    FOREIGN ND4T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.060 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.210 1.260 7.900 1.540 ;
        RECT  6.220 2.940 7.900 3.220 ;
        RECT  6.990 1.260 7.270 3.220 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.340 1.790 2.740 ;
        RECT  1.410 2.150 1.690 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.910 2.930 2.740 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.300 1.070 2.940 ;
        RECT  0.750 2.340 1.070 2.740 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.560 0.490 1.960 ;
        RECT  0.170 1.500 0.450 2.180 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.470 -0.380 3.870 0.560 ;
        RECT  5.260 -0.380 5.660 0.860 ;
        RECT  6.870 -0.380 7.270 0.860 ;
        RECT  0.000 -0.380 8.060 0.380 ;
        RECT  1.340 -0.380 1.740 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.700 4.480 3.100 5.420 ;
        RECT  5.600 4.260 6.000 5.420 ;
        RECT  6.870 4.260 7.270 5.420 ;
        RECT  0.000 4.660 8.060 5.420 ;
        RECT  1.540 4.480 1.940 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.340 2.870 5.110 3.110 ;
        RECT  4.870 1.280 5.110 3.110 ;
        RECT  6.270 1.780 6.510 2.700 ;
        RECT  5.730 1.780 6.510 2.020 ;
        RECT  5.730 1.280 5.970 2.020 ;
        RECT  4.340 1.280 5.970 1.520 ;
        RECT  1.650 4.000 4.770 4.240 ;
        RECT  4.530 3.520 4.770 4.240 ;
        RECT  0.750 3.940 1.890 4.180 ;
        RECT  1.650 3.040 1.890 4.240 ;
        RECT  4.530 3.520 5.590 3.760 ;
        RECT  5.350 2.250 5.590 3.760 ;
        RECT  1.650 3.040 3.620 3.280 ;
        RECT  3.380 1.370 3.620 3.280 ;
        RECT  2.270 1.370 3.620 1.610 ;
        RECT  2.270 1.020 2.510 1.610 ;
        RECT  0.160 1.020 2.510 1.260 ;
        RECT  2.130 3.520 4.100 3.760 ;
        RECT  3.860 0.890 4.100 3.760 ;
        RECT  3.860 2.330 4.630 2.570 ;
        RECT  2.750 0.890 4.100 1.130 ;
    END
END ND4T

MACRO NR2
    CLASS CORE ;
    FOREIGN NR2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.860 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.960 1.700 3.200 ;
        RECT  0.790 1.180 1.070 3.200 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.380 2.030 1.690 2.430 ;
        RECT  1.410 1.740 1.690 2.430 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.180 0.480 2.580 ;
        RECT  0.170 2.180 0.450 2.840 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 -0.380 1.700 0.640 ;
        RECT  0.000 -0.380 1.860 0.380 ;
        RECT  0.160 -0.380 0.560 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 1.860 5.420 ;
        RECT  0.160 3.830 0.560 5.420 ;
        END
    END VCC
END NR2

MACRO NR2F
    CLASS CORE ;
    FOREIGN NR2F 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.350 2.980 1.880 3.780 ;
        RECT  1.570 1.160 1.970 1.500 ;
        RECT  3.880 2.980 4.280 3.780 ;
        RECT  0.160 1.220 6.650 1.500 ;
        RECT  6.270 2.790 6.650 3.780 ;
        RECT  6.370 0.620 6.650 3.780 ;
        RECT  1.350 3.500 6.650 3.780 ;
        RECT  0.160 1.160 0.560 1.500 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.300 4.170 2.740 ;
        RECT  3.890 2.310 4.300 2.660 ;
        RECT  1.410 2.380 4.300 2.660 ;
        RECT  1.410 2.420 4.770 2.660 ;
        RECT  4.530 2.420 4.770 3.220 ;
        RECT  5.770 2.230 6.010 3.220 ;
        RECT  4.530 2.980 6.010 3.220 ;
        RECT  5.770 2.230 6.090 2.630 ;
        RECT  1.580 2.330 1.980 2.660 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.740 1.070 2.740 ;
        RECT  3.190 1.760 3.590 2.130 ;
        RECT  0.790 1.760 5.410 2.000 ;
        RECT  5.130 1.760 5.410 2.740 ;
        RECT  0.630 2.230 1.070 2.630 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 -0.380 2.640 0.780 ;
        RECT  3.700 -0.380 4.100 0.780 ;
        RECT  5.330 -0.380 5.730 0.910 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  0.860 -0.380 1.260 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.700 4.110 3.100 5.420 ;
        RECT  4.860 4.120 5.260 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  0.240 4.220 0.640 5.420 ;
        END
    END VCC
END NR2F

MACRO NR2P
    CLASS CORE ;
    FOREIGN NR2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.240 1.370 1.800 1.610 ;
        RECT  1.560 0.870 1.970 1.420 ;
        RECT  1.560 1.180 3.550 1.420 ;
        RECT  3.240 0.870 3.550 1.420 ;
        RECT  0.160 3.540 3.550 3.820 ;
        RECT  3.270 0.620 3.550 3.940 ;
        RECT  3.160 3.520 3.560 3.760 ;
        RECT  0.240 0.810 0.480 1.610 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.530 2.650 ;
        RECT  2.670 1.740 2.910 3.220 ;
        RECT  0.170 2.980 2.910 3.220 ;
        RECT  0.170 2.250 0.450 3.300 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.740 2.310 2.740 ;
        RECT  1.980 2.250 2.310 2.650 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.440 -0.380 2.840 0.940 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.920 -0.380 1.320 1.130 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  1.660 4.060 2.060 5.420 ;
        END
    END VCC
END NR2P

MACRO NR2T
    CLASS CORE ;
    FOREIGN NR2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 3.180 0.480 3.780 ;
        RECT  0.170 3.500 1.690 3.780 ;
        RECT  3.260 3.260 3.660 3.820 ;
        RECT  1.410 3.540 3.660 3.820 ;
        RECT  0.170 1.260 4.380 1.500 ;
        RECT  0.170 1.180 0.450 3.860 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.740 1.070 2.180 ;
        RECT  0.710 1.840 1.670 2.080 ;
        RECT  1.430 1.820 4.170 2.060 ;
        RECT  3.290 1.820 4.170 2.080 ;
        RECT  0.710 1.740 1.070 2.140 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.330 2.710 2.740 ;
        RECT  4.360 2.330 4.790 2.740 ;
        RECT  4.510 2.300 4.790 2.740 ;
        RECT  2.030 2.500 4.790 2.740 ;
        RECT  2.030 2.300 2.310 2.940 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.260 -0.380 3.660 1.020 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.560 -0.380 1.960 1.020 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.400 4.130 4.800 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  1.710 4.130 2.110 5.420 ;
        END
    END VCC
END NR2T

MACRO NR3
    CLASS CORE ;
    FOREIGN NR3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.100 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.620 2.790 2.930 3.190 ;
        RECT  2.650 1.180 2.930 3.300 ;
        RECT  0.160 1.260 2.930 1.500 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.230 1.830 1.690 2.230 ;
        RECT  1.410 1.740 1.690 2.230 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.980 0.530 2.380 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.740 2.310 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.380 2.940 0.940 ;
        RECT  0.000 -0.380 3.100 0.380 ;
        RECT  0.950 -0.380 1.350 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.100 5.420 ;
        RECT  0.160 4.180 0.560 5.420 ;
        END
    END VCC
END NR3

MACRO NR3H
    CLASS CORE ;
    FOREIGN NR3H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.190 3.450 1.280 3.690 ;
        RECT  0.160 1.570 4.160 1.810 ;
        RECT  0.190 1.570 0.430 3.690 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.050 2.930 2.960 ;
        RECT  2.590 2.250 2.930 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.930 4.790 2.650 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.130 2.650 ;
        RECT  0.790 2.050 1.070 3.160 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.690 -0.380 3.090 1.290 ;
        RECT  4.480 -0.380 4.880 1.290 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.880 -0.380 1.280 1.290 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  4.300 3.910 4.700 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.320 3.200 5.420 3.440 ;
        RECT  0.160 3.930 3.440 4.170 ;
    END
END NR3H

MACRO NR3HP
    CLASS CORE ;
    FOREIGN NR3HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 3.450 2.000 3.690 ;
        RECT  0.810 1.570 6.390 1.810 ;
        RECT  0.810 1.570 1.050 3.690 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.050 3.550 2.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 2.250 6.030 2.960 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 1.840 2.650 ;
        RECT  1.410 2.050 1.690 3.160 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 -0.380 2.070 1.290 ;
        RECT  2.610 -0.380 3.010 1.290 ;
        RECT  4.190 -0.380 4.590 1.290 ;
        RECT  5.200 -0.380 5.600 1.290 ;
        RECT  6.780 -0.380 7.180 1.290 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.160 -0.380 0.560 1.530 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.880 4.260 7.280 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  5.440 3.910 5.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.040 3.200 6.560 3.440 ;
        RECT  0.880 3.930 4.160 4.170 ;
        RECT  3.760 3.910 4.160 4.170 ;
    END
END NR3HP

MACRO NR3HT
    CLASS CORE ;
    FOREIGN NR3HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.810 3.450 4.160 3.690 ;
        RECT  0.810 1.570 13.210 1.810 ;
        RECT  0.810 1.570 1.050 3.690 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.050 6.650 2.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.250 12.230 2.960 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.250 2.460 2.650 ;
        RECT  2.030 2.050 2.310 3.160 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 -0.380 2.640 1.290 ;
        RECT  3.830 -0.380 4.230 1.290 ;
        RECT  4.770 -0.380 5.170 1.290 ;
        RECT  6.350 -0.380 7.330 1.290 ;
        RECT  8.510 -0.380 8.910 1.290 ;
        RECT  9.860 -0.380 10.260 1.290 ;
        RECT  11.440 -0.380 12.420 1.290 ;
        RECT  13.600 -0.380 14.000 1.290 ;
        RECT  0.000 -0.380 14.260 0.380 ;
        RECT  0.160 -0.380 0.560 1.530 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  11.540 4.260 11.940 5.420 ;
        RECT  12.980 4.260 13.380 5.420 ;
        RECT  0.000 4.660 14.260 5.420 ;
        RECT  10.100 3.910 10.500 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.200 3.200 14.100 3.440 ;
        RECT  0.160 3.930 9.210 4.170 ;
        RECT  8.810 3.910 9.210 4.170 ;
        RECT  4.480 3.910 4.880 4.170 ;
    END
END NR3HT

MACRO NR4
    CLASS CORE ;
    FOREIGN NR4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.720 2.790 6.030 3.190 ;
        RECT  5.750 1.180 6.030 3.300 ;
        RECT  5.720 1.490 6.030 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.250 2.310 3.300 ;
        RECT  1.980 2.250 2.310 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.830 2.930 2.740 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.200 1.260 2.740 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.550 2.210 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.520 -0.380 1.920 0.560 ;
        RECT  2.880 -0.380 3.280 0.560 ;
        RECT  4.920 -0.380 5.320 1.030 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.160 -0.380 0.560 0.840 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 4.080 3.580 5.420 ;
        RECT  4.840 3.710 5.240 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.160 4.010 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.860 2.960 5.480 3.200 ;
        RECT  5.240 2.150 5.480 3.200 ;
        RECT  3.860 2.800 4.220 3.200 ;
        RECT  3.860 1.650 4.100 3.200 ;
        RECT  5.240 2.150 5.510 2.550 ;
        RECT  3.680 1.490 3.920 1.890 ;
        RECT  1.210 3.080 1.740 3.320 ;
        RECT  1.500 0.800 1.740 3.320 ;
        RECT  4.590 1.840 4.830 2.550 ;
        RECT  4.340 1.840 4.830 2.080 ;
        RECT  4.340 0.800 4.580 2.080 ;
        RECT  0.750 1.280 1.740 1.520 ;
        RECT  1.500 0.800 4.580 1.040 ;
        RECT  1.930 3.540 3.410 3.780 ;
        RECT  3.170 1.280 3.410 3.780 ;
        RECT  3.170 2.210 3.620 2.610 ;
        RECT  2.130 1.280 3.410 1.520 ;
    END
END NR4

MACRO NR4P
    CLASS CORE ;
    FOREIGN NR4P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.180 6.030 3.300 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 3.300 ;
        RECT  1.980 2.250 2.310 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.830 2.930 2.740 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.200 1.920 1.690 2.320 ;
        RECT  1.410 1.680 1.690 2.320 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.480 2.650 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.350 -0.380 3.250 0.560 ;
        RECT  5.020 -0.380 5.420 1.080 ;
        RECT  6.260 -0.380 6.660 1.080 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  0.160 -0.380 0.560 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.320 4.020 3.720 5.420 ;
        RECT  5.020 4.130 5.420 5.420 ;
        RECT  6.260 4.130 6.660 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  0.160 4.010 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.860 2.960 5.390 3.200 ;
        RECT  5.150 2.250 5.390 3.200 ;
        RECT  3.860 1.490 4.100 3.200 ;
        RECT  5.150 2.250 5.480 2.650 ;
        RECT  3.650 1.490 4.100 1.890 ;
        RECT  0.720 2.980 1.610 3.220 ;
        RECT  0.720 1.200 0.960 3.220 ;
        RECT  4.530 2.030 4.800 2.430 ;
        RECT  4.530 0.800 4.770 2.430 ;
        RECT  0.830 0.700 1.070 1.600 ;
        RECT  1.900 0.800 4.770 1.040 ;
        RECT  0.830 0.700 2.140 0.940 ;
        RECT  1.930 3.540 3.410 3.780 ;
        RECT  3.170 1.280 3.410 3.780 ;
        RECT  3.170 2.250 3.620 2.650 ;
        RECT  2.130 1.280 3.410 1.520 ;
    END
END NR4P

MACRO NR4S
    CLASS CORE ;
    FOREIGN NR4S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.720 2.790 6.030 3.190 ;
        RECT  5.750 1.180 6.030 3.300 ;
        RECT  5.720 1.490 6.030 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.090 2.930 2.740 ;
        RECT  2.630 2.250 2.930 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.180 2.310 1.820 ;
        RECT  1.930 1.270 2.310 1.670 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.180 0.480 1.580 ;
        RECT  0.170 1.180 0.450 1.820 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.380 ;
        RECT  1.230 1.830 1.690 2.230 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.160 0.700 0.560 0.940 ;
        RECT  1.600 -0.380 2.000 0.940 ;
        RECT  3.110 -0.380 3.510 1.370 ;
        RECT  5.010 -0.380 5.410 0.640 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.160 -0.380 0.510 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.780 4.100 3.180 5.420 ;
        RECT  4.220 4.100 4.620 5.420 ;
        RECT  4.920 3.050 5.320 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  1.340 3.250 1.740 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.500 4.180 3.900 4.420 ;
        RECT  3.660 3.620 3.900 4.420 ;
        RECT  3.660 3.620 4.680 3.860 ;
        RECT  4.440 1.050 4.680 3.860 ;
        RECT  4.440 2.330 5.370 2.570 ;
        RECT  4.290 1.050 4.690 1.290 ;
        RECT  3.960 1.610 4.200 3.380 ;
        RECT  2.520 2.980 4.200 3.220 ;
        RECT  2.550 1.610 4.200 1.850 ;
        RECT  2.550 0.700 2.790 1.850 ;
        RECT  2.320 0.700 2.790 0.940 ;
        RECT  2.040 3.620 3.380 3.860 ;
        RECT  3.140 3.460 3.380 3.860 ;
        RECT  2.040 2.770 2.280 3.860 ;
        RECT  0.240 2.770 0.480 3.190 ;
        RECT  0.240 2.770 2.280 3.010 ;
        RECT  0.750 1.280 0.990 3.010 ;
        RECT  0.930 0.620 1.170 1.520 ;
        RECT  0.930 0.620 1.200 1.020 ;
    END
END NR4S

MACRO NR4T
    CLASS CORE ;
    FOREIGN NR4T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.640 1.540 7.280 1.780 ;
        RECT  5.640 2.870 7.280 3.110 ;
        RECT  6.370 1.540 6.650 3.110 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 3.300 ;
        RECT  1.980 2.250 2.310 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.830 2.930 2.740 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.200 1.920 1.690 2.320 ;
        RECT  1.410 1.680 1.690 2.320 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.480 2.650 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 3.220 0.560 ;
        RECT  4.990 -0.380 5.390 1.080 ;
        RECT  6.230 -0.380 6.630 1.080 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.160 -0.380 0.560 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.290 4.020 3.690 5.420 ;
        RECT  4.990 4.130 5.390 5.420 ;
        RECT  6.230 4.130 6.630 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.160 4.010 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.860 2.960 5.360 3.200 ;
        RECT  5.120 2.250 5.360 3.200 ;
        RECT  3.860 1.490 4.100 3.200 ;
        RECT  5.120 2.250 5.480 2.650 ;
        RECT  3.650 1.490 4.100 1.890 ;
        RECT  0.720 2.980 1.610 3.220 ;
        RECT  0.720 1.200 0.960 3.220 ;
        RECT  4.500 2.030 4.800 2.430 ;
        RECT  4.500 0.800 4.740 2.430 ;
        RECT  0.830 0.700 1.070 1.600 ;
        RECT  1.840 0.800 4.740 1.040 ;
        RECT  0.830 0.700 2.080 0.940 ;
        RECT  1.930 3.540 3.410 3.780 ;
        RECT  3.170 1.280 3.410 3.780 ;
        RECT  3.170 2.250 3.620 2.650 ;
        RECT  2.130 1.280 3.410 1.520 ;
    END
END NR4T

MACRO OA112
    CLASS CORE ;
    FOREIGN OA112 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.380 3.340 4.790 3.740 ;
        RECT  4.510 0.620 4.790 3.860 ;
        RECT  4.480 1.490 4.790 1.890 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.880 ;
        RECT  1.310 2.270 1.690 2.670 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.270 0.550 2.670 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.230 3.550 3.300 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.270 2.410 2.670 ;
        RECT  2.030 1.740 2.310 2.880 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.820 -0.380 4.220 1.060 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  2.090 -0.380 2.510 0.980 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.400 4.260 3.800 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  1.100 3.740 1.500 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.120 3.540 4.080 3.780 ;
        RECT  3.840 2.270 4.080 3.780 ;
        RECT  2.120 3.230 2.360 3.780 ;
        RECT  0.170 3.230 2.360 3.470 ;
        RECT  0.810 1.260 1.050 3.470 ;
        RECT  0.170 3.000 0.570 3.470 ;
        RECT  3.840 2.270 4.260 2.670 ;
        RECT  0.160 1.260 1.050 1.500 ;
        RECT  1.370 1.260 3.310 1.500 ;
    END
END OA112

MACRO OA112P
    CLASS CORE ;
    FOREIGN OA112P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.380 3.340 4.790 3.740 ;
        RECT  4.510 1.350 4.790 3.860 ;
        RECT  4.380 1.490 4.790 1.890 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.780 1.690 2.880 ;
        RECT  1.310 2.270 1.690 2.670 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.270 0.550 2.670 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.210 3.550 3.300 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.270 2.410 2.670 ;
        RECT  2.030 1.780 2.310 2.880 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.580 -0.380 3.980 1.500 ;
        RECT  5.020 -0.380 5.420 0.950 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  2.040 -0.380 2.460 0.960 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.400 4.260 3.800 5.420 ;
        RECT  5.020 4.260 5.420 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  1.100 3.740 1.500 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.120 3.540 4.080 3.780 ;
        RECT  3.840 2.250 4.080 3.780 ;
        RECT  2.120 3.230 2.360 3.780 ;
        RECT  0.170 3.230 2.360 3.470 ;
        RECT  0.810 1.260 1.050 3.470 ;
        RECT  0.170 3.000 0.570 3.470 ;
        RECT  3.840 2.250 4.260 2.650 ;
        RECT  0.160 1.260 1.050 1.500 ;
        RECT  1.370 1.300 3.250 1.540 ;
    END
END OA112P

MACRO OA112S
    CLASS CORE ;
    FOREIGN OA112S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.380 3.150 4.790 3.550 ;
        RECT  4.510 1.170 4.790 3.860 ;
        RECT  4.480 1.490 4.790 1.890 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.880 ;
        RECT  1.310 2.270 1.690 2.670 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.270 0.550 2.670 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.100 3.550 2.750 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.270 2.410 2.670 ;
        RECT  2.030 1.740 2.310 2.880 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.820 -0.380 4.220 0.900 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  2.110 -0.380 2.510 1.020 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.350 3.490 3.790 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  1.100 3.740 1.500 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.170 3.230 2.800 3.470 ;
        RECT  3.840 2.420 4.080 3.230 ;
        RECT  2.560 2.990 4.080 3.230 ;
        RECT  0.810 1.260 1.050 3.470 ;
        RECT  0.170 3.060 0.570 3.470 ;
        RECT  3.840 2.420 4.260 2.820 ;
        RECT  0.160 1.260 1.050 1.500 ;
        RECT  1.370 1.260 3.310 1.500 ;
    END
END OA112S

MACRO OA112T
    CLASS CORE ;
    FOREIGN OA112T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 1.570 5.410 3.670 ;
        RECT  4.200 1.570 6.040 1.810 ;
        RECT  4.280 3.430 6.040 3.670 ;
        RECT  4.280 3.430 4.520 3.830 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.830 1.690 2.880 ;
        RECT  1.310 2.270 1.690 2.670 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.270 0.550 2.670 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.210 3.550 3.300 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.270 2.410 2.670 ;
        RECT  2.030 1.830 2.310 2.880 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.480 -0.380 3.880 1.500 ;
        RECT  4.920 -0.380 5.320 0.950 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  1.970 -0.380 2.370 0.910 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.400 4.260 3.800 5.420 ;
        RECT  4.920 4.260 5.320 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  1.100 3.740 1.500 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.120 3.540 4.030 3.780 ;
        RECT  3.790 2.250 4.030 3.780 ;
        RECT  2.120 3.230 2.360 3.780 ;
        RECT  0.170 3.230 2.360 3.470 ;
        RECT  0.810 1.260 1.050 3.470 ;
        RECT  0.170 3.000 0.570 3.470 ;
        RECT  3.790 2.250 4.260 2.650 ;
        RECT  0.160 1.260 1.050 1.500 ;
        RECT  1.370 1.350 3.160 1.590 ;
    END
END OA112T

MACRO OA12
    CLASS CORE ;
    FOREIGN OA12 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.180 3.550 3.300 ;
        RECT  3.170 2.900 3.550 3.300 ;
        RECT  3.210 1.270 3.550 1.670 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.600 1.070 3.860 ;
        RECT  0.600 2.770 1.070 3.170 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.600 1.690 3.310 ;
        RECT  1.310 2.600 1.690 3.000 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 3.310 ;
        RECT  2.020 2.600 2.310 3.000 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  2.390 -0.380 2.810 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.480 4.030 2.920 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.150 4.000 0.570 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.440 3.550 2.800 3.790 ;
        RECT  2.560 1.820 2.800 3.790 ;
        RECT  2.560 2.150 3.030 2.550 ;
        RECT  0.880 1.820 2.800 2.060 ;
        RECT  0.880 1.260 1.280 2.060 ;
        RECT  0.160 0.770 0.560 1.580 ;
        RECT  1.580 0.770 2.000 1.570 ;
        RECT  0.160 0.770 2.000 1.010 ;
    END
END OA12

MACRO OA12P
    CLASS CORE ;
    FOREIGN OA12P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.170 2.860 3.550 3.260 ;
        RECT  3.270 0.620 3.550 3.290 ;
        RECT  3.140 1.300 3.550 1.700 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.030 0.550 2.430 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 2.260 1.760 2.740 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.260 2.310 3.300 ;
        RECT  2.020 2.260 2.310 2.660 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.800 -0.380 4.180 1.070 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  2.410 -0.380 2.810 1.100 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.430 4.040 2.830 5.420 ;
        RECT  3.770 4.130 4.200 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.150 4.110 0.570 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.440 3.550 2.860 3.790 ;
        RECT  2.620 1.780 2.860 3.790 ;
        RECT  2.620 2.150 3.030 2.550 ;
        RECT  0.880 1.780 2.860 2.020 ;
        RECT  0.880 1.540 1.280 2.020 ;
        RECT  1.600 1.060 2.000 1.540 ;
        RECT  0.160 1.060 0.560 1.500 ;
        RECT  0.160 1.060 2.000 1.300 ;
    END
END OA12P

MACRO OA12S
    CLASS CORE ;
    FOREIGN OA12S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.240 3.470 3.550 3.870 ;
        RECT  3.270 1.180 3.550 4.420 ;
        RECT  3.240 1.490 3.550 1.890 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.670 1.070 3.310 ;
        RECT  0.550 2.670 1.070 3.070 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.300 1.690 3.310 ;
        RECT  1.310 2.670 1.690 3.070 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 3.310 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  2.450 -0.380 2.820 1.040 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.350 4.030 2.780 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.150 4.000 0.570 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.440 3.550 3.000 3.790 ;
        RECT  2.760 1.820 3.000 3.790 ;
        RECT  0.960 1.820 3.000 2.060 ;
        RECT  0.960 1.220 1.200 2.060 ;
        RECT  0.240 0.720 0.480 1.620 ;
        RECT  1.600 0.720 2.000 1.540 ;
        RECT  0.240 0.720 2.000 0.960 ;
    END
END OA12S

MACRO OA12T
    CLASS CORE ;
    FOREIGN OA12T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 1.400 4.800 1.640 ;
        RECT  3.090 2.940 4.800 3.180 ;
        RECT  3.890 1.400 4.170 3.180 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.030 0.550 2.430 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 2.260 1.760 2.740 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.260 2.310 3.300 ;
        RECT  2.020 2.260 2.310 2.660 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.760 -0.380 4.140 1.080 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  2.410 -0.380 2.810 1.100 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.410 4.040 2.810 5.420 ;
        RECT  3.770 4.130 4.200 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.150 4.110 0.570 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.440 3.550 2.850 3.790 ;
        RECT  2.610 1.780 2.850 3.790 ;
        RECT  2.610 2.150 3.030 2.550 ;
        RECT  0.880 1.780 2.850 2.020 ;
        RECT  0.880 1.540 1.280 2.020 ;
        RECT  1.600 1.060 2.000 1.540 ;
        RECT  0.160 1.060 0.560 1.500 ;
        RECT  0.160 1.060 2.000 1.300 ;
    END
END OA12T

MACRO OA13
    CLASS CORE ;
    FOREIGN OA13 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 2.790 4.790 3.190 ;
        RECT  4.510 0.620 4.790 3.300 ;
        RECT  4.480 1.490 4.790 1.890 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 2.140 0.550 2.740 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 1.740 1.690 2.370 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 2.160 2.340 2.740 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.890 3.060 2.290 ;
        RECT  2.650 1.740 2.930 2.290 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 -0.380 2.070 0.560 ;
        RECT  3.910 -0.380 4.260 1.060 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.800 4.010 4.200 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.160 3.840 0.600 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.160 3.540 3.660 3.780 ;
        RECT  3.420 1.180 3.660 3.780 ;
        RECT  3.420 2.130 4.030 2.530 ;
        RECT  3.250 1.180 3.660 1.580 ;
        RECT  0.880 1.260 2.850 1.500 ;
    END
END OA13

MACRO OA13P
    CLASS CORE ;
    FOREIGN OA13P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.490 4.790 3.190 ;
        RECT  4.380 2.790 4.790 3.190 ;
        RECT  4.480 1.490 4.790 1.890 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 2.140 0.550 2.740 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 1.740 1.690 2.370 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 2.160 2.340 2.740 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.740 2.930 2.390 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 -0.380 2.070 0.560 ;
        RECT  3.770 -0.380 4.170 0.990 ;
        RECT  5.020 -0.380 5.420 0.990 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.680 4.140 4.080 5.420 ;
        RECT  5.020 4.180 5.420 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.180 4.260 0.580 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.160 3.540 3.500 3.780 ;
        RECT  3.260 1.260 3.500 3.780 ;
        RECT  3.260 2.130 4.000 2.530 ;
        RECT  3.020 1.260 3.500 1.500 ;
        RECT  0.880 1.260 2.700 1.500 ;
    END
END OA13P

MACRO OA13S
    CLASS CORE ;
    FOREIGN OA13S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.850 2.810 4.170 3.210 ;
        RECT  3.890 0.620 4.170 3.300 ;
        RECT  3.860 0.660 4.170 1.060 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 2.110 0.780 2.350 ;
        RECT  0.160 1.180 0.460 2.350 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.740 ;
        RECT  1.190 2.160 1.690 2.560 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 2.160 2.340 2.740 ;
        RECT  1.930 2.160 2.340 2.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.630 2.160 2.950 3.300 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 -0.380 2.060 0.940 ;
        RECT  3.000 -0.380 3.370 1.010 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.160 -0.380 0.560 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.960 4.110 3.370 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.160 3.710 0.600 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.100 3.540 3.460 3.780 ;
        RECT  3.220 1.490 3.460 3.780 ;
        RECT  3.220 2.150 3.580 2.550 ;
        RECT  3.170 1.490 3.460 1.890 ;
        RECT  2.420 1.260 2.660 1.890 ;
        RECT  0.930 1.260 1.170 1.890 ;
        RECT  0.930 1.260 2.660 1.500 ;
    END
END OA13S

MACRO OA13T
    CLASS CORE ;
    FOREIGN OA13T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.400 1.570 6.040 1.810 ;
        RECT  4.300 2.870 6.040 3.110 ;
        RECT  5.130 1.570 5.410 3.110 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 2.140 0.550 2.740 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 1.740 1.690 2.370 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 2.160 2.340 2.740 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.740 2.930 2.390 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 -0.380 2.070 0.560 ;
        RECT  3.770 -0.380 4.170 0.990 ;
        RECT  5.020 -0.380 5.420 0.990 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.680 4.140 4.080 5.420 ;
        RECT  5.020 4.180 5.420 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.180 4.260 0.580 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.160 3.540 3.500 3.780 ;
        RECT  3.260 1.260 3.500 3.780 ;
        RECT  3.260 2.130 4.000 2.530 ;
        RECT  3.020 1.260 3.500 1.500 ;
        RECT  0.880 1.260 2.700 1.500 ;
    END
END OA13T

MACRO OA22
    CLASS CORE ;
    FOREIGN OA22 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.760 3.120 4.170 3.520 ;
        RECT  3.890 0.620 4.170 3.860 ;
        RECT  3.860 1.410 4.170 1.810 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.610 3.020 2.010 ;
        RECT  2.650 1.610 2.970 2.180 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.010 2.300 2.330 2.880 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.300 1.690 3.300 ;
        RECT  1.260 2.480 1.690 2.880 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.880 0.490 2.280 ;
        RECT  0.170 1.740 0.450 2.760 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.200 -0.380 3.600 1.010 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  1.590 -0.380 2.030 0.670 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.970 4.020 3.390 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.150 4.390 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.750 3.540 3.460 3.780 ;
        RECT  3.220 2.230 3.460 3.780 ;
        RECT  0.750 1.400 0.990 3.780 ;
        RECT  3.220 2.230 3.650 2.630 ;
        RECT  0.750 1.400 1.350 1.640 ;
        RECT  1.670 1.820 2.140 2.060 ;
        RECT  1.670 0.920 1.910 2.060 ;
        RECT  0.240 0.920 0.480 1.500 ;
        RECT  1.670 1.000 2.810 1.240 ;
        RECT  0.240 0.920 1.910 1.160 ;
    END
END OA22

MACRO OA222
    CLASS CORE ;
    FOREIGN OA222 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.100 3.000 5.410 3.400 ;
        RECT  5.130 0.620 5.410 3.860 ;
        RECT  5.100 1.290 5.410 1.690 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 3.300 ;
        RECT  1.980 2.410 2.310 2.810 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.300 2.930 3.300 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.080 0.490 2.480 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.300 1.690 3.300 ;
        RECT  1.210 2.460 1.690 2.860 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.400 3.590 2.800 ;
        RECT  3.270 2.300 3.550 3.300 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.460 4.270 2.860 ;
        RECT  3.890 2.300 4.170 3.300 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.300 -0.380 4.700 1.130 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  2.860 -0.380 3.260 1.130 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.340 4.090 4.740 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  1.500 4.110 1.900 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.540 4.770 3.780 ;
        RECT  4.530 1.830 4.770 3.780 ;
        RECT  0.730 1.220 0.970 3.780 ;
        RECT  4.530 1.830 4.880 2.230 ;
        RECT  0.470 1.220 0.970 1.460 ;
        RECT  2.040 1.440 2.440 1.860 ;
        RECT  2.040 1.440 3.900 1.680 ;
        RECT  3.660 0.810 3.900 1.680 ;
        RECT  1.340 0.680 1.580 1.940 ;
        RECT  1.340 0.680 1.590 1.080 ;
    END
END OA222

MACRO OA222P
    CLASS CORE ;
    FOREIGN OA222P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 0.620 6.030 3.860 ;
        RECT  5.740 1.270 6.030 1.670 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 3.300 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.400 3.030 2.800 ;
        RECT  2.650 2.300 2.930 3.300 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.270 0.560 2.670 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.300 1.690 3.300 ;
        RECT  1.300 2.460 1.690 2.860 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.300 4.170 3.300 ;
        RECT  3.790 2.390 4.170 2.790 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.740 4.790 2.740 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.930 -0.380 5.330 0.920 ;
        RECT  6.320 -0.380 6.650 0.970 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  3.340 -0.380 3.660 1.530 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.990 4.100 5.430 5.420 ;
        RECT  6.220 4.100 6.670 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  1.590 4.120 1.990 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.540 5.390 3.780 ;
        RECT  5.150 2.180 5.390 3.780 ;
        RECT  0.810 1.140 1.050 3.780 ;
        RECT  5.150 2.180 5.490 2.580 ;
        RECT  2.380 1.770 4.140 2.010 ;
        RECT  3.900 1.230 4.140 2.010 ;
        RECT  3.900 1.230 4.540 1.470 ;
        RECT  1.640 0.680 1.880 1.980 ;
    END
END OA222P

MACRO OA222S
    CLASS CORE ;
    FOREIGN OA222S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.100 3.000 5.410 3.400 ;
        RECT  5.130 0.620 5.410 3.860 ;
        RECT  5.100 1.210 5.410 1.610 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 3.300 ;
        RECT  1.980 2.410 2.310 2.810 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.300 2.930 3.300 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.490 2.650 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.300 1.690 3.300 ;
        RECT  1.210 2.460 1.690 2.860 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.400 3.580 2.800 ;
        RECT  3.270 2.300 3.550 3.300 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.460 4.260 2.860 ;
        RECT  3.890 2.300 4.170 3.300 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.300 -0.380 4.700 1.470 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  2.860 -0.380 3.180 1.550 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 4.060 4.650 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  1.430 4.030 1.850 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.540 4.770 3.780 ;
        RECT  4.530 1.830 4.770 3.780 ;
        RECT  0.730 1.120 0.970 3.780 ;
        RECT  4.530 1.830 4.880 2.230 ;
        RECT  0.550 1.120 0.970 1.520 ;
        RECT  2.040 1.790 3.660 2.030 ;
        RECT  3.420 1.150 3.660 2.030 ;
        RECT  2.040 1.620 2.440 2.030 ;
        RECT  3.420 1.230 3.980 1.470 ;
        RECT  1.340 0.680 1.580 1.940 ;
        RECT  1.340 0.680 1.590 1.080 ;
    END
END OA222S

MACRO OA222T
    CLASS CORE ;
    FOREIGN OA222T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.540 1.370 7.280 1.610 ;
        RECT  5.600 3.050 7.280 3.290 ;
        RECT  6.370 1.370 6.650 3.290 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 3.300 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.400 3.030 2.800 ;
        RECT  2.650 2.300 2.930 3.300 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.270 0.560 2.670 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.300 1.690 3.300 ;
        RECT  1.300 2.460 1.690 2.860 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.300 4.170 3.300 ;
        RECT  3.720 2.390 4.170 2.790 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.740 4.790 2.740 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.930 -0.380 5.330 0.820 ;
        RECT  6.320 -0.380 6.650 0.900 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  3.340 -0.380 3.660 1.530 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.960 4.100 5.400 5.420 ;
        RECT  6.220 4.100 6.670 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  1.590 4.140 1.990 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.540 5.360 3.780 ;
        RECT  5.120 2.180 5.360 3.780 ;
        RECT  0.810 1.140 1.050 3.780 ;
        RECT  5.120 2.180 5.490 2.580 ;
        RECT  2.380 1.770 4.140 2.010 ;
        RECT  3.900 1.230 4.140 2.010 ;
        RECT  3.900 1.230 4.540 1.470 ;
        RECT  1.620 0.680 1.860 1.980 ;
    END
END OA222T

MACRO OA22P
    CLASS CORE ;
    FOREIGN OA22P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 0.620 4.790 3.300 ;
        RECT  4.390 2.900 4.790 3.300 ;
        RECT  4.380 1.410 4.790 1.810 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.740 3.550 2.740 ;
        RECT  3.180 2.180 3.550 2.580 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.740 2.930 2.740 ;
        RECT  2.320 2.180 2.930 2.580 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.180 1.690 3.300 ;
        RECT  1.310 2.180 1.690 2.580 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.180 0.580 2.740 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.710 -0.380 4.110 0.950 ;
        RECT  5.030 -0.380 5.450 1.030 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  2.120 -0.380 2.520 0.960 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.440 4.030 3.920 5.420 ;
        RECT  4.990 4.080 5.440 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.160 4.160 0.570 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.820 3.540 4.040 3.780 ;
        RECT  3.800 2.180 4.040 3.780 ;
        RECT  1.960 3.070 2.200 3.780 ;
        RECT  0.820 1.390 1.060 3.780 ;
        RECT  3.800 2.180 4.200 2.580 ;
        RECT  0.820 1.390 1.210 1.790 ;
        RECT  1.610 1.260 2.010 1.810 ;
        RECT  1.610 1.260 3.310 1.500 ;
        RECT  0.250 0.720 0.490 1.430 ;
        RECT  1.610 0.720 1.850 1.810 ;
        RECT  0.250 0.720 1.850 0.960 ;
    END
END OA22P

MACRO OA22S
    CLASS CORE ;
    FOREIGN OA22S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.860 3.100 4.170 3.500 ;
        RECT  3.890 1.180 4.170 3.860 ;
        RECT  3.860 1.490 4.170 1.890 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.740 2.970 2.140 ;
        RECT  2.650 1.550 2.930 2.180 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.010 2.300 2.330 2.880 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.300 1.690 3.300 ;
        RECT  1.260 2.480 1.690 2.880 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.320 0.490 2.720 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.200 -0.380 3.600 1.010 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  1.610 -0.380 2.010 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.970 4.040 3.390 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.150 4.390 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.750 3.540 3.530 3.780 ;
        RECT  3.290 2.230 3.530 3.780 ;
        RECT  0.750 1.820 0.990 3.780 ;
        RECT  3.290 2.230 3.650 2.630 ;
        RECT  0.750 1.820 1.350 2.060 ;
        RECT  1.670 1.820 2.070 2.060 ;
        RECT  1.670 0.990 1.910 2.060 ;
        RECT  0.240 0.990 0.480 1.500 ;
        RECT  0.240 0.990 2.800 1.230 ;
    END
END OA22S

MACRO OA22T
    CLASS CORE ;
    FOREIGN OA22T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.330 1.490 6.040 1.730 ;
        RECT  4.310 2.980 6.040 3.220 ;
        RECT  5.130 1.490 5.410 3.220 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.740 3.550 2.740 ;
        RECT  3.180 2.180 3.550 2.580 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.740 2.930 2.740 ;
        RECT  2.320 2.180 2.930 2.580 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.180 1.690 3.300 ;
        RECT  1.310 2.180 1.690 2.580 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.180 0.580 2.740 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.710 -0.380 4.110 1.000 ;
        RECT  5.030 -0.380 5.450 1.080 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  2.120 -0.380 2.520 0.960 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.440 4.030 3.920 5.420 ;
        RECT  4.990 4.080 5.440 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.160 4.160 0.570 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.820 3.540 4.040 3.780 ;
        RECT  3.800 2.180 4.040 3.780 ;
        RECT  1.960 3.070 2.200 3.780 ;
        RECT  0.820 1.390 1.060 3.780 ;
        RECT  3.800 2.180 4.200 2.580 ;
        RECT  0.820 1.390 1.210 1.790 ;
        RECT  1.610 1.260 2.010 1.810 ;
        RECT  1.610 1.260 3.310 1.500 ;
        RECT  0.250 0.720 0.490 1.430 ;
        RECT  1.610 0.720 1.850 1.810 ;
        RECT  0.250 0.720 1.850 0.960 ;
    END
END OA22T

MACRO OAI112H
    CLASS CORE ;
    FOREIGN OAI112H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.570 6.560 1.810 ;
        RECT  2.320 3.040 6.560 3.280 ;
        RECT  5.750 1.570 6.030 3.280 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.810 2.550 ;
        RECT  4.510 2.150 4.790 2.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.650 2.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.150 1.070 2.800 ;
        RECT  0.730 2.150 1.070 2.550 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.410 2.550 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.000 3.900 4.400 5.420 ;
        RECT  5.440 4.260 5.840 5.420 ;
        RECT  6.880 4.260 7.280 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.000 1.090 7.280 1.330 ;
        RECT  0.880 1.570 5.120 1.810 ;
        RECT  0.160 3.700 3.440 3.940 ;
    END
END OAI112H

MACRO OAI112HP
    CLASS CORE ;
    FOREIGN OAI112HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 1.570 12.140 1.810 ;
        RECT  3.760 3.040 12.140 3.280 ;
        RECT  10.090 1.570 10.370 3.280 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.150 8.530 2.550 ;
        RECT  8.230 2.150 8.510 2.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.150 11.610 2.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.310 2.800 ;
        RECT  1.970 2.150 2.310 2.550 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.890 2.550 ;
        RECT  4.510 2.150 4.790 2.800 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  5.920 -0.380 6.320 1.330 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.260 2.720 5.420 ;
        RECT  6.700 3.930 7.100 5.420 ;
        RECT  8.140 4.260 8.540 5.420 ;
        RECT  9.580 4.260 9.980 5.420 ;
        RECT  11.020 4.260 11.420 5.420 ;
        RECT  12.460 4.260 12.860 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.700 1.090 12.860 1.330 ;
        RECT  0.880 1.570 9.260 1.810 ;
        RECT  0.160 3.700 6.320 3.940 ;
    END
END OAI112HP

MACRO OAI112HS
    CLASS CORE ;
    FOREIGN OAI112HS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.340 3.690 3.550 3.930 ;
        RECT  3.270 1.570 4.180 1.810 ;
        RECT  3.270 1.570 3.550 3.930 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.150 2.930 2.790 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.150 4.170 2.790 ;
        RECT  3.860 2.150 4.170 2.550 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.150 0.510 2.550 ;
        RECT  0.170 2.150 0.450 2.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.150 1.690 2.800 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.340 4.170 2.740 5.420 ;
        RECT  3.780 4.260 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.190 3.000 1.430 ;
    END
END OAI112HS

MACRO OAI112HT
    CLASS CORE ;
    FOREIGN OAI112HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.220 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.850 1.570 18.340 1.810 ;
        RECT  5.200 3.040 18.340 3.280 ;
        RECT  15.050 1.570 15.330 3.280 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 2.150 12.870 2.550 ;
        RECT  12.570 2.150 12.850 2.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.910 2.150 17.190 2.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.310 2.800 ;
        RECT  1.970 2.150 2.310 2.550 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.750 2.550 ;
        RECT  6.370 2.150 6.650 2.800 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  5.920 -0.380 6.320 0.950 ;
        RECT  7.360 -0.380 7.760 0.950 ;
        RECT  8.800 -0.380 9.700 1.330 ;
        RECT  0.000 -0.380 19.220 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.260 2.720 5.420 ;
        RECT  3.760 4.260 4.160 5.420 ;
        RECT  9.520 3.930 10.420 5.420 ;
        RECT  11.460 4.260 11.860 5.420 ;
        RECT  12.900 4.260 13.300 5.420 ;
        RECT  14.340 4.260 14.740 5.420 ;
        RECT  15.780 4.260 16.180 5.420 ;
        RECT  17.220 4.260 17.620 5.420 ;
        RECT  18.660 4.260 19.060 5.420 ;
        RECT  0.000 4.660 19.220 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.020 1.090 19.060 1.330 ;
        RECT  0.880 1.570 14.020 1.810 ;
        RECT  0.160 3.700 9.200 3.940 ;
    END
END OAI112HT

MACRO OAI12H
    CLASS CORE ;
    FOREIGN OAI12H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.720 1.090 6.030 1.490 ;
        RECT  5.750 1.090 6.030 3.450 ;
        RECT  2.320 3.210 6.040 3.450 ;
        RECT  4.200 1.090 6.030 1.330 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.150 1.070 2.800 ;
        RECT  0.730 2.150 1.070 2.550 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.410 2.550 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.810 2.550 ;
        RECT  4.510 2.150 4.790 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.370 -0.380 3.770 0.950 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.960 4.170 4.360 5.420 ;
        RECT  5.640 4.260 6.040 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.570 5.320 1.810 ;
        RECT  0.160 3.780 3.440 4.020 ;
    END
END OAI12H

MACRO OAI12HP
    CLASS CORE ;
    FOREIGN OAI12HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.540 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.060 1.090 10.370 1.490 ;
        RECT  10.090 1.090 10.370 3.450 ;
        RECT  3.760 3.210 10.370 3.450 ;
        RECT  7.100 1.090 10.370 1.330 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.150 1.690 2.800 ;
        RECT  1.350 2.150 1.690 2.550 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.790 2.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.150 8.530 2.550 ;
        RECT  8.230 2.150 8.510 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  6.250 -0.380 6.650 0.950 ;
        RECT  0.000 -0.380 10.540 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.260 2.720 5.420 ;
        RECT  6.860 4.170 7.260 5.420 ;
        RECT  8.540 4.260 8.940 5.420 ;
        RECT  9.980 4.260 10.380 5.420 ;
        RECT  0.000 4.660 10.540 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.570 9.660 1.810 ;
        RECT  0.160 3.780 6.320 4.020 ;
    END
END OAI12HP

MACRO OAI12HS
    CLASS CORE ;
    FOREIGN OAI12HS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.240 3.290 3.550 3.690 ;
        RECT  3.270 1.490 3.550 3.690 ;
        RECT  1.480 3.450 3.550 3.690 ;
        RECT  3.240 1.490 3.550 1.890 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.510 2.650 ;
        RECT  0.170 2.250 0.450 2.890 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 1.690 2.900 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.250 2.930 2.890 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 1.110 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.440 3.930 2.840 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.570 2.840 1.810 ;
    END
END OAI12HS

MACRO OAI12HT
    CLASS CORE ;
    FOREIGN OAI12HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.400 1.090 14.710 1.490 ;
        RECT  14.430 1.090 14.710 3.450 ;
        RECT  5.200 3.210 14.710 3.450 ;
        RECT  9.890 1.090 14.710 1.330 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 2.150 7.270 2.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.570 2.150 12.870 2.550 ;
        RECT  12.570 2.150 12.850 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  5.920 -0.380 6.320 0.950 ;
        RECT  7.360 -0.380 7.760 0.950 ;
        RECT  9.130 -0.380 9.530 0.950 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.260 2.720 5.420 ;
        RECT  3.760 4.260 4.160 5.420 ;
        RECT  9.650 4.170 10.050 5.420 ;
        RECT  11.440 4.260 11.840 5.420 ;
        RECT  12.880 4.260 13.280 5.420 ;
        RECT  14.320 4.260 14.720 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.570 14.000 1.810 ;
        RECT  0.160 3.780 9.200 4.020 ;
    END
END OAI12HT

MACRO OAI13H
    CLASS CORE ;
    FOREIGN OAI13H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.060 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.160 3.700 5.060 3.940 ;
        RECT  6.860 1.190 7.270 1.590 ;
        RECT  6.990 1.190 7.270 3.610 ;
        RECT  4.820 3.370 7.900 3.610 ;
        RECT  4.820 3.370 5.060 3.940 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.690 2.250 6.030 2.650 ;
        RECT  5.750 1.860 6.030 2.650 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.210 2.130 3.550 2.530 ;
        RECT  3.270 1.890 3.550 2.530 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.010 1.690 2.650 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.510 2.250 7.890 2.650 ;
        RECT  7.610 2.010 7.890 2.650 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.940 1.110 ;
        RECT  5.340 -0.380 5.740 0.950 ;
        RECT  0.000 -0.380 8.060 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.780 3.850 7.180 5.420 ;
        RECT  0.000 4.660 8.060 5.420 ;
        RECT  5.300 3.910 5.700 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.350 5.020 1.590 ;
        RECT  6.140 0.710 6.380 1.430 ;
        RECT  4.780 1.190 6.380 1.430 ;
        RECT  6.140 0.710 7.900 0.950 ;
        RECT  3.040 3.220 4.580 3.460 ;
        RECT  4.340 2.890 4.580 3.460 ;
        RECT  4.340 2.890 6.420 3.130 ;
        RECT  0.880 4.180 4.160 4.420 ;
    END
END OAI13H

MACRO OAI13HP
    CLASS CORE ;
    FOREIGN OAI13HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.400 1.190 15.240 1.430 ;
        RECT  0.880 3.370 15.240 3.610 ;
        RECT  14.430 1.190 14.710 3.610 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.710 1.670 10.990 2.650 ;
        RECT  10.650 2.030 10.990 2.430 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.690 2.130 6.030 2.530 ;
        RECT  5.750 1.890 6.030 2.530 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.250 2.370 2.650 ;
        RECT  2.030 2.010 2.310 2.650 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.570 2.250 15.950 2.650 ;
        RECT  15.670 2.010 15.950 2.650 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.110 -0.380 4.510 0.950 ;
        RECT  5.550 -0.380 5.950 0.950 ;
        RECT  6.990 -0.380 7.390 0.950 ;
        RECT  8.140 -0.380 8.540 0.950 ;
        RECT  9.580 -0.380 9.980 0.950 ;
        RECT  11.020 -0.380 11.920 0.950 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  11.240 4.260 11.640 5.420 ;
        RECT  12.680 4.260 13.080 5.420 ;
        RECT  14.120 4.200 14.520 5.420 ;
        RECT  15.560 4.260 15.960 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  9.800 3.910 10.200 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.190 13.000 1.430 ;
        RECT  12.760 0.710 13.000 1.430 ;
        RECT  12.760 0.710 15.960 0.950 ;
        RECT  5.200 2.890 13.800 3.130 ;
        RECT  0.160 3.850 9.200 4.090 ;
    END
END OAI13HP

MACRO OAI13HS
    CLASS CORE ;
    FOREIGN OAI13HS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 3.700 5.230 3.940 ;
        RECT  6.340 1.490 6.650 1.890 ;
        RECT  6.340 3.270 6.650 3.670 ;
        RECT  4.990 3.430 6.650 3.670 ;
        RECT  6.370 1.490 6.650 3.770 ;
        RECT  4.990 3.430 5.230 3.940 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.450 2.250 4.790 2.650 ;
        RECT  4.510 1.930 4.790 2.650 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.590 2.250 2.930 2.650 ;
        RECT  2.650 2.010 2.930 2.650 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.130 2.650 ;
        RECT  0.790 2.010 1.070 2.650 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 2.010 6.030 2.650 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.690 -0.380 3.090 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.470 3.910 5.870 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  3.760 4.260 4.160 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 1.190 5.940 1.430 ;
        RECT  2.320 3.220 4.720 3.460 ;
        RECT  4.480 2.950 4.720 3.460 ;
        RECT  4.480 2.950 4.880 3.190 ;
        RECT  0.160 4.180 3.440 4.420 ;
    END
END OAI13HS

MACRO OAI13HT
    CLASS CORE ;
    FOREIGN OAI13HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.320 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  18.160 1.190 21.440 1.430 ;
        RECT  0.160 3.370 22.160 3.610 ;
        RECT  20.010 1.190 20.290 3.610 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.050 1.670 15.330 2.650 ;
        RECT  14.990 2.030 15.330 2.430 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.790 2.130 9.130 2.530 ;
        RECT  8.850 1.890 9.130 2.530 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.250 2.990 2.650 ;
        RECT  2.650 2.010 2.930 2.650 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  21.250 1.790 21.530 2.570 ;
        RECT  21.150 2.030 21.530 2.430 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.480 -0.380 5.380 0.950 ;
        RECT  6.050 -0.380 6.450 0.950 ;
        RECT  7.490 -0.380 7.890 0.950 ;
        RECT  8.930 -0.380 9.330 0.950 ;
        RECT  10.370 -0.380 10.770 0.950 ;
        RECT  11.530 -0.380 11.930 0.950 ;
        RECT  12.970 -0.380 13.370 0.950 ;
        RECT  14.410 -0.380 14.810 0.950 ;
        RECT  15.850 -0.380 16.750 0.950 ;
        RECT  0.000 -0.380 22.320 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  15.280 4.260 15.680 5.420 ;
        RECT  16.720 4.260 17.120 5.420 ;
        RECT  18.160 4.260 18.560 5.420 ;
        RECT  19.600 4.200 20.000 5.420 ;
        RECT  21.040 4.260 21.440 5.420 ;
        RECT  0.000 4.660 22.320 5.420 ;
        RECT  13.840 3.910 14.240 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.190 17.760 1.430 ;
        RECT  17.520 0.710 17.760 1.430 ;
        RECT  17.520 0.710 22.160 0.950 ;
        RECT  7.360 2.890 19.280 3.130 ;
        RECT  0.880 3.850 12.800 4.090 ;
    END
END OAI13HT

MACRO OAI222H
    CLASS CORE ;
    FOREIGN OAI222H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.320 3.170 9.130 3.410 ;
        RECT  8.440 1.570 10.280 1.810 ;
        RECT  8.850 1.570 9.130 3.410 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.770 2.550 ;
        RECT  6.370 2.150 6.650 2.790 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.930 2.550 ;
        RECT  4.510 2.150 4.790 2.790 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.150 8.530 2.550 ;
        RECT  8.230 2.150 8.510 2.790 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.150 10.370 2.790 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.410 2.550 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.150 1.070 2.800 ;
        RECT  0.730 2.150 1.070 2.550 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 1.070 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.280 4.260 6.680 5.420 ;
        RECT  9.880 4.260 10.280 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.840 1.190 7.960 1.430 ;
        RECT  7.720 0.710 7.960 1.430 ;
        RECT  7.720 0.710 11.000 0.950 ;
        RECT  7.720 3.780 11.000 4.020 ;
        RECT  0.880 1.310 4.520 1.550 ;
        RECT  4.280 0.710 4.520 1.550 ;
        RECT  4.280 0.710 7.400 0.950 ;
        RECT  4.120 3.780 7.400 4.020 ;
        RECT  0.160 3.780 3.440 4.020 ;
    END
END OAI222H

MACRO OAI222HP
    CLASS CORE ;
    FOREIGN OAI222HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.840 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.760 3.170 16.080 3.410 ;
        RECT  14.240 1.570 18.960 1.810 ;
        RECT  15.670 1.570 15.950 3.410 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.150 11.610 2.790 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.150 8.510 2.790 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 2.150 14.730 2.550 ;
        RECT  14.430 2.150 14.710 2.790 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  18.150 2.150 18.430 2.790 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.890 2.550 ;
        RECT  4.510 2.150 4.790 2.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.150 1.690 2.800 ;
        RECT  1.350 2.150 1.690 2.550 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  5.920 -0.380 6.320 1.070 ;
        RECT  0.000 -0.380 19.840 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.260 2.720 5.420 ;
        RECT  10.600 4.260 11.000 5.420 ;
        RECT  12.040 4.260 12.440 5.420 ;
        RECT  17.120 4.260 17.520 5.420 ;
        RECT  18.560 4.260 18.960 5.420 ;
        RECT  0.000 4.660 19.840 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.720 1.570 13.760 1.810 ;
        RECT  13.520 1.090 13.760 1.810 ;
        RECT  13.520 1.090 19.680 1.330 ;
        RECT  13.520 3.780 19.680 4.020 ;
        RECT  0.880 1.310 7.400 1.550 ;
        RECT  7.160 1.090 13.160 1.330 ;
        RECT  7.000 3.780 13.160 4.020 ;
        RECT  0.160 3.780 6.320 4.020 ;
    END
END OAI222HP

MACRO OAI222HT
    CLASS CORE ;
    FOREIGN OAI222HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 28.520 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.200 3.170 23.390 3.410 ;
        RECT  20.040 1.570 27.640 1.810 ;
        RECT  23.110 1.570 23.390 3.410 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 2.150 16.570 2.790 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.150 12.230 2.790 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  21.250 2.150 21.530 2.790 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  26.210 2.150 26.490 2.790 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.650 2.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  5.920 -0.380 6.320 0.950 ;
        RECT  7.360 -0.380 7.760 0.950 ;
        RECT  8.800 -0.380 9.200 1.070 ;
        RECT  0.000 -0.380 28.520 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.260 2.720 5.420 ;
        RECT  3.760 4.260 4.160 5.420 ;
        RECT  14.920 4.260 15.320 5.420 ;
        RECT  16.360 4.260 16.760 5.420 ;
        RECT  17.800 4.260 18.200 5.420 ;
        RECT  24.360 4.260 24.760 5.420 ;
        RECT  25.800 4.260 26.200 5.420 ;
        RECT  27.240 4.260 27.640 5.420 ;
        RECT  0.000 4.660 28.520 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.600 1.570 19.560 1.810 ;
        RECT  19.320 1.090 19.560 1.810 ;
        RECT  19.320 1.090 28.360 1.330 ;
        RECT  19.320 3.780 28.360 4.020 ;
        RECT  0.880 1.310 10.280 1.550 ;
        RECT  10.040 1.090 18.920 1.330 ;
        RECT  9.880 3.780 18.920 4.020 ;
        RECT  0.160 3.780 9.200 4.020 ;
    END
END OAI222HT

MACRO OAI222S
    CLASS CORE ;
    FOREIGN OAI222S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.180 4.790 3.780 ;
        RECT  2.150 3.540 5.340 3.780 ;
        RECT  4.370 1.480 4.790 1.880 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.320 2.250 3.560 2.650 ;
        RECT  3.270 2.300 3.550 3.300 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.300 2.930 3.300 ;
        RECT  2.450 2.250 2.690 2.650 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 2.250 5.410 3.300 ;
        RECT  5.030 2.250 5.410 2.650 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.250 4.270 2.650 ;
        RECT  3.890 2.250 4.170 3.300 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 1.730 2.650 ;
        RECT  1.410 2.250 1.690 3.300 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.070 3.270 ;
        RECT  0.690 2.250 1.070 2.650 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.140 -0.380 0.580 0.940 ;
        RECT  1.470 -0.380 1.940 0.940 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.240 -0.380 0.480 1.020 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.480 4.060 3.900 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.170 3.920 0.570 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.090 0.700 5.390 1.700 ;
        RECT  2.210 1.110 2.790 1.350 ;
        RECT  2.550 0.700 2.790 1.350 ;
        RECT  3.760 0.700 4.160 0.950 ;
        RECT  2.550 0.700 5.390 0.940 ;
        RECT  0.720 1.600 3.420 1.840 ;
        RECT  3.020 1.550 3.420 1.840 ;
        RECT  0.720 1.560 1.120 1.840 ;
    END
END OAI222S

MACRO OAI22H
    CLASS CORE ;
    FOREIGN OAI22H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.320 3.300 5.410 3.540 ;
        RECT  4.720 1.370 6.560 1.610 ;
        RECT  5.130 1.370 5.410 3.540 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.150 1.070 2.800 ;
        RECT  0.730 2.150 1.070 2.550 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.410 2.550 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.810 2.550 ;
        RECT  4.510 2.150 4.790 2.790 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.650 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 1.330 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.160 4.260 6.560 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.570 4.320 1.810 ;
        RECT  4.080 0.890 4.320 1.810 ;
        RECT  4.080 0.890 7.280 1.130 ;
        RECT  4.000 3.780 7.280 4.020 ;
        RECT  0.160 3.780 3.440 4.020 ;
    END
END OAI22H

MACRO OAI22HP
    CLASS CORE ;
    FOREIGN OAI22HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.020 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.760 3.300 9.750 3.540 ;
        RECT  7.420 1.370 12.140 1.610 ;
        RECT  9.470 1.370 9.750 3.540 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.150 1.690 2.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.150 4.790 2.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.150 8.510 2.790 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.150 11.610 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.050 -0.380 3.450 0.950 ;
        RECT  3.040 0.710 3.450 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  5.920 -0.380 6.320 1.070 ;
        RECT  0.000 -0.380 13.020 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.260 2.720 5.420 ;
        RECT  10.300 4.260 10.700 5.420 ;
        RECT  11.740 4.260 12.140 5.420 ;
        RECT  0.000 4.660 13.020 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.570 7.020 1.810 ;
        RECT  6.780 0.890 7.020 1.810 ;
        RECT  6.780 0.890 12.860 1.130 ;
        RECT  6.700 3.780 12.860 4.020 ;
        RECT  0.160 3.780 6.320 4.020 ;
    END
END OAI22HP

MACRO OAI22HT
    CLASS CORE ;
    FOREIGN OAI22HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.220 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.200 3.300 14.090 3.540 ;
        RECT  10.740 1.370 18.340 1.610 ;
        RECT  13.810 1.370 14.090 3.540 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.150 2.310 2.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 2.150 6.650 2.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.150 12.230 2.790 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.290 2.150 16.570 2.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.480 -0.380 4.880 0.950 ;
        RECT  5.930 -0.380 6.330 0.950 ;
        RECT  5.920 0.710 6.330 0.950 ;
        RECT  7.360 -0.380 7.760 0.950 ;
        RECT  8.800 -0.380 9.700 1.070 ;
        RECT  0.000 -0.380 19.220 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.260 2.720 5.420 ;
        RECT  3.760 4.260 4.160 5.420 ;
        RECT  15.060 4.260 15.460 5.420 ;
        RECT  16.500 4.260 16.900 5.420 ;
        RECT  17.940 4.260 18.340 5.420 ;
        RECT  0.000 4.660 19.220 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 1.570 10.340 1.810 ;
        RECT  10.100 0.890 10.340 1.810 ;
        RECT  10.100 0.890 19.060 1.130 ;
        RECT  10.020 3.780 19.060 4.020 ;
        RECT  0.160 3.780 9.200 4.020 ;
    END
END OAI22HT

MACRO OAI22S
    CLASS CORE ;
    FOREIGN OAI22S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.980 4.100 2.930 4.340 ;
        RECT  2.650 1.180 2.930 4.420 ;
        RECT  2.520 1.320 2.930 1.720 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.700 2.230 1.070 2.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.230 1.730 2.630 ;
        RECT  1.410 2.230 1.690 3.300 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.230 2.410 2.630 ;
        RECT  2.030 2.230 2.310 3.300 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.740 3.550 2.740 ;
        RECT  3.190 2.230 3.550 2.630 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.790 1.270 1.340 1.510 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.790 -0.380 1.070 1.510 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.240 3.830 3.560 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.300 4.020 0.700 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.240 1.750 2.040 1.990 ;
        RECT  1.800 0.700 2.040 1.990 ;
        RECT  0.240 1.260 0.480 1.990 ;
        RECT  3.160 0.700 3.560 1.060 ;
        RECT  1.800 0.700 3.560 0.940 ;
    END
END OAI22S

MACRO OR2
    CLASS CORE ;
    FOREIGN OR2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 1.490 2.330 1.890 ;
        RECT  2.030 2.790 2.310 4.420 ;
        RECT  2.090 1.490 2.330 3.190 ;
        RECT  2.000 2.790 2.330 3.190 ;
        RECT  2.030 0.620 2.310 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.530 0.480 2.930 ;
        RECT  0.170 2.300 0.450 2.930 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.110 1.250 2.350 ;
        RECT  0.790 2.110 1.070 2.770 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  1.340 -0.380 1.740 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  1.410 4.180 1.730 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.170 1.760 3.410 ;
        RECT  1.520 1.570 1.760 3.410 ;
        RECT  1.520 2.130 1.850 2.530 ;
        RECT  0.440 1.570 1.760 1.810 ;
    END
END OR2

MACRO OR2B1
    CLASS CORE ;
    FOREIGN OR2B1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.240 2.790 3.530 3.190 ;
        RECT  3.290 1.180 3.530 3.300 ;
        RECT  3.240 1.450 3.530 1.850 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.640 1.690 2.280 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.230 0.480 2.630 ;
        RECT  0.170 2.230 0.450 2.940 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.270 -0.380 2.670 0.560 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.970 -0.380 1.370 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.160 4.400 2.670 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.340 3.500 2.900 3.740 ;
        RECT  2.660 1.160 2.900 3.740 ;
        RECT  2.660 2.230 3.030 2.630 ;
        RECT  1.740 1.160 2.900 1.400 ;
        RECT  0.610 3.400 1.050 3.640 ;
        RECT  0.810 1.160 1.050 3.640 ;
        RECT  0.810 2.980 2.350 3.220 ;
        RECT  2.110 1.830 2.350 3.220 ;
        RECT  0.180 1.160 1.050 1.400 ;
    END
END OR2B1

MACRO OR2B1P
    CLASS CORE ;
    FOREIGN OR2B1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.240 1.260 4.170 1.540 ;
        RECT  3.890 1.260 4.170 3.220 ;
        RECT  3.190 2.940 4.170 3.220 ;
        RECT  3.240 1.260 3.480 1.840 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.640 2.310 2.280 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.230 0.480 2.630 ;
        RECT  0.170 1.970 0.450 2.830 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.950 -0.380 1.350 0.560 ;
        RECT  1.680 -0.380 2.080 0.560 ;
        RECT  2.370 -0.380 2.770 0.560 ;
        RECT  3.780 -0.380 4.180 0.940 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.300 -0.380 0.700 0.390 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 4.130 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.420 4.130 0.820 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.430 2.980 2.900 3.220 ;
        RECT  2.660 1.080 2.900 3.220 ;
        RECT  2.660 2.310 3.450 2.550 ;
        RECT  1.740 1.080 2.900 1.320 ;
        RECT  0.750 3.190 1.050 3.590 ;
        RECT  0.810 1.240 1.050 3.590 ;
        RECT  0.810 1.820 1.690 2.060 ;
        RECT  0.180 1.240 1.050 1.480 ;
    END
END OR2B1P

MACRO OR2B1S
    CLASS CORE ;
    FOREIGN OR2B1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.100 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.180 2.930 3.220 ;
        RECT  1.740 2.940 2.930 3.220 ;
        RECT  2.620 1.180 2.930 1.580 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.020 0.480 2.420 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.540 1.690 2.180 ;
        RECT  1.400 1.720 1.690 2.120 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.100 0.380 ;
        RECT  1.020 -0.380 1.420 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 3.910 2.940 5.420 ;
        RECT  0.000 4.660 3.100 5.420 ;
        RECT  0.950 4.060 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.540 0.960 3.780 ;
        RECT  0.720 1.260 0.960 3.780 ;
        RECT  0.720 2.420 2.400 2.660 ;
        RECT  0.160 1.260 0.960 1.500 ;
    END
END OR2B1S

MACRO OR2B1T
    CLASS CORE ;
    FOREIGN OR2B1T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.260 6.030 3.220 ;
        RECT  4.900 1.260 6.660 1.540 ;
        RECT  5.020 2.940 6.660 3.220 ;
        RECT  4.900 1.190 5.140 1.590 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.040 3.550 2.740 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.950 0.480 2.840 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.590 -0.380 2.990 1.320 ;
        RECT  1.230 -0.380 3.720 0.490 ;
        RECT  4.100 -0.380 4.500 0.940 ;
        RECT  5.540 -0.380 5.940 0.940 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  1.230 -0.380 1.470 1.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.260 4.220 3.660 5.420 ;
        RECT  4.500 4.120 4.900 5.420 ;
        RECT  5.750 4.120 6.150 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  0.480 4.160 0.880 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.820 2.960 2.910 3.200 ;
        RECT  2.670 1.560 2.910 3.200 ;
        RECT  4.410 2.180 5.430 2.420 ;
        RECT  4.410 1.560 4.650 2.420 ;
        RECT  1.950 1.560 4.650 1.800 ;
        RECT  3.390 1.000 3.630 1.800 ;
        RECT  1.950 1.000 2.190 1.800 ;
        RECT  1.300 3.770 2.940 4.010 ;
        RECT  3.860 2.980 4.100 3.980 ;
        RECT  2.700 3.740 4.100 3.980 ;
        RECT  0.570 3.360 1.050 3.760 ;
        RECT  0.810 1.680 1.050 3.760 ;
        RECT  0.810 2.170 2.230 2.410 ;
        RECT  0.750 1.240 0.990 1.920 ;
        RECT  0.320 1.240 0.990 1.480 ;
    END
END OR2B1T

MACRO OR2P
    CLASS CORE ;
    FOREIGN OR2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.620 2.790 2.930 3.190 ;
        RECT  2.650 0.620 2.930 3.300 ;
        RECT  2.520 1.490 2.930 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.550 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 2.100 1.690 2.500 ;
        RECT  1.410 1.740 1.690 2.500 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.720 -0.380 2.120 1.020 ;
        RECT  3.190 -0.380 3.560 1.030 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.160 -0.380 0.560 1.500 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.160 4.140 3.560 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  1.530 4.050 1.930 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.320 3.520 2.270 3.760 ;
        RECT  2.030 1.260 2.270 3.760 ;
        RECT  0.320 2.980 0.560 3.760 ;
        RECT  0.160 2.980 0.560 3.220 ;
        RECT  0.880 1.260 2.270 1.500 ;
    END
END OR2P

MACRO OR2S
    CLASS CORE ;
    FOREIGN OR2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.370 2.310 3.580 ;
        RECT  2.000 3.180 2.310 3.580 ;
        RECT  2.000 1.370 2.310 1.770 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.490 0.480 2.890 ;
        RECT  0.170 2.120 0.450 3.100 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.910 1.150 2.310 ;
        RECT  0.790 1.660 1.070 2.830 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.450 -0.380 1.610 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.900 4.480 1.300 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 4.180 0.660 4.420 ;
        RECT  0.420 3.520 0.660 4.420 ;
        RECT  0.420 3.520 1.760 3.760 ;
        RECT  1.520 1.040 1.760 3.760 ;
        RECT  1.520 2.490 1.790 2.890 ;
        RECT  0.450 1.040 1.760 1.280 ;
    END
END OR2S

MACRO OR2T
    CLASS CORE ;
    FOREIGN OR2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.260 6.040 1.540 ;
        RECT  3.890 2.940 6.040 3.220 ;
        RECT  5.130 1.260 5.410 3.220 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.720 2.100 1.070 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.100 3.000 2.740 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.920 -0.380 2.320 1.500 ;
        RECT  3.480 -0.380 3.880 0.940 ;
        RECT  4.920 -0.380 5.320 0.940 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.410 -0.380 0.810 1.500 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.880 3.810 4.280 5.420 ;
        RECT  5.130 4.120 5.530 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  2.280 4.260 2.680 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.900 2.980 1.140 3.920 ;
        RECT  0.900 2.980 3.530 3.220 ;
        RECT  3.290 1.260 3.530 3.220 ;
        RECT  1.310 1.100 1.550 3.220 ;
        RECT  3.290 2.140 4.770 2.540 ;
        RECT  2.640 1.260 3.530 1.500 ;
        RECT  1.210 1.100 1.550 1.500 ;
        RECT  0.280 4.160 1.790 4.400 ;
        RECT  1.550 3.460 1.790 4.400 ;
        RECT  0.280 2.980 0.520 4.400 ;
        RECT  1.550 3.460 3.400 3.700 ;
        RECT  0.200 2.980 0.600 3.220 ;
    END
END OR2T

MACRO OR3
    CLASS CORE ;
    FOREIGN OR3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.240 2.790 3.550 3.190 ;
        RECT  3.270 1.180 3.550 3.300 ;
        RECT  3.240 1.350 3.550 1.750 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.740 ;
        RECT  1.350 1.910 1.690 2.310 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.740 2.310 2.740 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.740 1.070 2.740 ;
        RECT  0.670 1.910 1.070 2.310 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.650 -0.380 3.050 0.980 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  1.020 -0.380 1.420 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  2.320 4.090 2.720 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.190 2.790 0.480 3.190 ;
        RECT  0.190 1.260 0.430 3.190 ;
        RECT  2.760 2.250 3.030 2.650 ;
        RECT  2.760 1.260 3.000 2.650 ;
        RECT  0.190 1.260 3.000 1.500 ;
    END
END OR3

MACRO OR3B1
    CLASS CORE ;
    FOREIGN OR3B1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 2.790 4.790 3.190 ;
        RECT  4.510 1.180 4.790 3.300 ;
        RECT  4.480 1.490 4.790 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 1.690 3.300 ;
        RECT  1.220 2.250 1.690 2.650 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.480 2.540 ;
        RECT  0.170 1.740 0.450 2.740 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 -0.380 2.600 0.560 ;
        RECT  3.680 -0.380 4.080 0.970 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.020 -0.380 1.420 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.680 4.180 4.080 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  1.040 4.030 1.440 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.040 2.790 3.280 3.190 ;
        RECT  3.040 2.790 4.150 3.030 ;
        RECT  3.910 1.390 4.150 3.030 ;
        RECT  1.610 1.390 4.150 1.630 ;
        RECT  0.720 3.540 2.790 3.780 ;
        RECT  2.550 2.030 2.790 3.780 ;
        RECT  0.160 3.430 0.960 3.670 ;
        RECT  0.720 1.260 0.960 3.780 ;
        RECT  2.550 2.030 3.030 2.430 ;
        RECT  0.160 1.260 0.960 1.500 ;
    END
END OR3B1

MACRO OR3B1P
    CLASS CORE ;
    FOREIGN OR3B1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 2.790 4.790 3.190 ;
        RECT  4.510 0.620 4.790 3.300 ;
        RECT  4.480 1.490 4.790 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.740 2.310 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 1.690 3.300 ;
        RECT  1.220 2.250 1.690 2.650 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.480 2.540 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 -0.380 2.700 0.640 ;
        RECT  3.780 -0.380 4.180 0.990 ;
        RECT  5.060 -0.380 5.380 1.070 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.820 -0.380 1.220 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 4.140 4.180 5.420 ;
        RECT  5.020 4.140 5.420 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  1.040 4.150 1.440 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.070 2.960 4.150 3.200 ;
        RECT  3.910 1.260 4.150 3.200 ;
        RECT  3.070 2.790 3.310 3.200 ;
        RECT  1.610 1.260 4.150 1.500 ;
        RECT  0.160 3.540 2.790 3.780 ;
        RECT  2.550 2.030 2.790 3.780 ;
        RECT  0.720 1.260 0.960 3.780 ;
        RECT  2.550 2.030 2.980 2.430 ;
        RECT  0.160 1.260 0.960 1.500 ;
    END
END OR3B1P

MACRO OR3B1S
    CLASS CORE ;
    FOREIGN OR3B1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 3.150 4.790 3.550 ;
        RECT  4.510 0.620 4.790 3.860 ;
        RECT  4.480 0.770 4.790 1.170 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.250 2.320 2.650 ;
        RECT  2.030 1.740 2.310 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.740 ;
        RECT  1.400 2.250 1.690 2.650 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.700 0.480 3.100 ;
        RECT  0.170 2.660 0.450 3.300 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.380 2.940 1.020 ;
        RECT  3.680 -0.380 4.080 1.170 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.960 -0.380 1.360 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.680 3.510 4.080 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  1.020 4.020 1.420 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.040 2.790 3.280 3.190 ;
        RECT  3.040 2.790 4.150 3.030 ;
        RECT  3.910 1.570 4.150 3.030 ;
        RECT  3.200 1.570 4.150 1.810 ;
        RECT  3.200 1.260 3.440 1.810 ;
        RECT  1.750 1.260 3.440 1.500 ;
        RECT  0.160 3.540 2.800 3.780 ;
        RECT  2.560 2.050 2.800 3.780 ;
        RECT  0.720 1.260 0.960 3.780 ;
        RECT  2.560 2.050 3.010 2.450 ;
        RECT  0.160 1.260 0.960 1.500 ;
    END
END OR3B1S

MACRO OR3B1T
    CLASS CORE ;
    FOREIGN OR3B1T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 2.870 4.720 3.270 ;
        RECT  5.130 1.570 5.410 3.110 ;
        RECT  4.480 1.570 6.040 1.810 ;
        RECT  4.480 2.870 6.040 3.110 ;
        RECT  4.480 1.410 4.720 1.810 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.740 2.310 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 1.690 3.300 ;
        RECT  1.220 2.250 1.690 2.650 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.480 2.540 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 -0.380 2.700 0.640 ;
        RECT  3.780 -0.380 4.180 0.990 ;
        RECT  5.060 -0.380 5.380 1.070 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.820 -0.380 1.220 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 4.140 4.180 5.420 ;
        RECT  5.020 4.140 5.420 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  1.040 4.150 1.440 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.070 2.950 4.150 3.190 ;
        RECT  3.910 1.260 4.150 3.190 ;
        RECT  3.070 2.790 3.310 3.190 ;
        RECT  1.610 1.260 4.150 1.500 ;
        RECT  0.160 3.540 2.790 3.780 ;
        RECT  2.550 2.030 2.790 3.780 ;
        RECT  0.720 1.260 0.960 3.780 ;
        RECT  2.550 2.030 2.980 2.430 ;
        RECT  0.160 1.260 0.960 1.500 ;
    END
END OR3B1T

MACRO OR3B2
    CLASS CORE ;
    FOREIGN OR3B2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.640 3.050 2.930 3.330 ;
        RECT  2.650 0.620 2.930 3.830 ;
        RECT  2.650 3.550 3.560 3.830 ;
        RECT  1.520 0.700 2.930 0.940 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.160 0.550 2.750 ;
        RECT  0.170 1.740 0.450 2.750 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.300 3.550 3.300 ;
        RECT  3.170 2.320 3.550 2.720 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.010 2.300 2.410 2.770 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.200 -0.380 3.560 0.860 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.610 -0.380 1.010 1.090 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 4.130 2.820 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  1.040 4.130 1.440 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.540 1.050 3.780 ;
        RECT  0.810 1.490 1.050 3.780 ;
        RECT  0.810 2.420 1.730 2.660 ;
        RECT  0.690 1.490 1.050 1.890 ;
    END
END OR3B2

MACRO OR3B2P
    CLASS CORE ;
    FOREIGN OR3B2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.020 1.260 6.030 1.540 ;
        RECT  5.750 1.260 6.030 3.220 ;
        RECT  5.100 2.940 6.030 3.220 ;
        RECT  5.100 2.880 5.340 3.280 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.960 1.690 2.620 ;
        RECT  1.310 1.960 1.690 2.360 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.730 1.070 3.430 ;
        RECT  0.720 2.910 1.070 3.310 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.720 4.330 2.740 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.670 1.360 1.050 1.760 ;
        RECT  0.810 -0.380 2.560 0.560 ;
        RECT  4.400 -0.380 4.800 0.780 ;
        RECT  5.640 -0.380 6.040 0.780 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.810 -0.380 1.050 1.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.400 4.260 4.800 5.420 ;
        RECT  5.640 4.260 6.040 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  1.190 4.260 1.590 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.930 3.620 4.810 3.860 ;
        RECT  4.570 2.200 4.810 3.860 ;
        RECT  2.930 1.360 3.170 3.860 ;
        RECT  4.570 2.200 5.220 2.440 ;
        RECT  1.310 1.440 3.170 1.680 ;
        RECT  3.410 2.980 3.900 3.380 ;
        RECT  3.410 1.080 3.650 3.380 ;
        RECT  3.410 1.080 3.930 1.480 ;
        RECT  0.190 3.770 2.260 4.010 ;
        RECT  2.020 2.030 2.260 4.010 ;
        RECT  0.190 0.620 0.430 4.010 ;
        RECT  0.160 0.620 0.560 0.860 ;
    END
END OR3B2P

MACRO OR3B2S
    CLASS CORE ;
    FOREIGN OR3B2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.220 2.930 3.330 ;
        RECT  1.640 3.050 3.560 3.330 ;
        RECT  1.520 1.220 2.930 1.500 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.800 0.570 3.300 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.170 2.300 3.550 2.810 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.010 1.740 2.410 2.770 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.160 -0.380 3.560 0.560 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.380 -0.380 0.780 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.370 4.480 2.770 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  1.040 4.480 1.440 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.540 1.050 3.780 ;
        RECT  0.810 1.570 1.050 3.780 ;
        RECT  0.810 2.420 1.730 2.660 ;
        RECT  0.380 1.570 1.050 1.810 ;
    END
END OR3B2S

MACRO OR3B2T
    CLASS CORE ;
    FOREIGN OR3B2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.260 6.030 3.220 ;
        RECT  5.000 1.260 6.660 1.540 ;
        RECT  5.080 2.940 6.660 3.220 ;
        RECT  5.080 2.940 5.320 3.340 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.030 1.690 2.730 ;
        RECT  1.310 2.030 1.690 2.430 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.730 1.070 3.430 ;
        RECT  0.670 2.910 1.070 3.310 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.330 2.520 ;
        RECT  3.890 1.720 4.170 2.740 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.670 1.360 1.050 1.760 ;
        RECT  0.810 -0.380 2.560 0.560 ;
        RECT  4.380 -0.380 4.780 0.780 ;
        RECT  5.620 -0.380 6.020 0.780 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  0.810 -0.380 1.050 1.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.380 4.260 4.780 5.420 ;
        RECT  5.620 4.260 6.020 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  1.030 4.260 1.430 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.930 3.620 4.840 3.860 ;
        RECT  4.600 2.200 4.840 3.860 ;
        RECT  2.930 1.360 3.170 3.860 ;
        RECT  4.600 2.200 5.200 2.440 ;
        RECT  1.420 1.440 3.170 1.680 ;
        RECT  3.410 2.980 3.910 3.380 ;
        RECT  3.410 1.080 3.650 3.380 ;
        RECT  3.410 1.080 3.910 1.480 ;
        RECT  0.190 3.770 2.260 4.010 ;
        RECT  2.020 2.060 2.260 4.010 ;
        RECT  0.190 0.620 0.430 4.010 ;
        RECT  0.160 0.620 0.560 0.860 ;
    END
END OR3B2T

MACRO OR3P
    CLASS CORE ;
    FOREIGN OR3P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 0.620 3.550 3.300 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.740 ;
        RECT  1.350 1.910 1.690 2.310 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.740 2.310 2.740 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.740 1.070 2.740 ;
        RECT  0.670 1.910 1.070 2.310 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.380 2.940 0.980 ;
        RECT  3.810 -0.380 4.180 0.980 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  1.020 -0.380 1.420 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 4.090 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  2.200 4.090 2.600 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.190 2.790 0.480 3.190 ;
        RECT  0.190 1.260 0.430 3.190 ;
        RECT  2.670 2.250 2.980 2.650 ;
        RECT  2.670 1.260 2.910 2.650 ;
        RECT  0.190 1.260 2.910 1.500 ;
    END
END OR3P

MACRO OR3S
    CLASS CORE ;
    FOREIGN OR3S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.240 2.790 3.550 3.190 ;
        RECT  3.270 1.010 3.550 3.300 ;
        RECT  3.240 1.180 3.550 1.580 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.740 ;
        RECT  1.350 1.910 1.690 2.310 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.910 2.310 2.740 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.740 1.070 2.740 ;
        RECT  0.670 1.910 1.070 2.310 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.370 -0.380 2.770 0.560 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.950 -0.380 1.350 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  2.340 3.350 2.740 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.190 2.790 0.480 3.190 ;
        RECT  0.190 1.260 0.430 3.190 ;
        RECT  2.670 2.250 2.980 2.650 ;
        RECT  2.670 1.260 2.910 2.650 ;
        RECT  0.160 1.260 2.910 1.500 ;
    END
END OR3S

MACRO OR3T
    CLASS CORE ;
    FOREIGN OR3T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.140 1.430 4.800 1.670 ;
        RECT  3.140 2.870 4.800 3.110 ;
        RECT  3.890 1.430 4.170 3.110 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.740 1.690 2.740 ;
        RECT  1.320 1.910 1.690 2.310 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.740 2.310 2.740 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.740 1.070 2.740 ;
        RECT  0.640 1.910 1.070 2.310 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.470 -0.380 2.870 0.980 ;
        RECT  3.740 -0.380 4.110 0.980 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.020 -0.380 1.420 0.650 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.710 4.090 4.110 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  2.140 4.090 2.540 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 2.790 0.480 3.190 ;
        RECT  0.160 1.260 0.400 3.190 ;
        RECT  2.600 2.230 3.110 2.630 ;
        RECT  2.600 1.260 2.840 2.630 ;
        RECT  0.160 1.260 2.840 1.500 ;
    END
END OR3T

MACRO PDI
    CLASS CORE ;
    FOREIGN PDI 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 0.660 2.310 2.180 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.270 0.490 2.670 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END EB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.730 -0.380 1.130 1.050 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.790 3.590 1.070 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.810 1.490 1.050 3.190 ;
        RECT  0.810 2.080 1.170 2.480 ;
        RECT  0.710 1.490 1.050 1.890 ;
    END
END PDI

MACRO PDIX
    CLASS CORE ;
    FOREIGN PDIX 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 0.630 4.170 1.720 ;
        RECT  3.720 0.630 4.170 0.870 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.190 0.480 2.590 ;
        RECT  0.170 2.190 0.450 2.840 ;
        END
    END EB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.540 -0.380 1.940 0.950 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.520 -0.380 0.840 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 4.480 1.540 5.420 ;
        RECT  2.490 4.480 2.890 5.420 ;
        RECT  3.840 4.480 4.800 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.440 4.010 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.520 3.220 0.960 3.620 ;
        RECT  0.720 1.420 0.960 3.620 ;
        RECT  0.720 2.100 1.600 2.340 ;
        RECT  0.690 1.420 0.960 1.820 ;
    END
END PDIX

MACRO PUI
    CLASS CORE ;
    FOREIGN PUI 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 3.400 ;
        RECT  2.000 2.790 2.310 3.190 ;
        END
    END O
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.220 0.490 2.620 ;
        RECT  0.170 2.200 0.450 2.840 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.710 -0.380 1.150 1.030 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.690 4.110 1.660 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.730 2.790 1.050 3.190 ;
        RECT  0.810 1.490 1.050 3.190 ;
        RECT  0.810 2.080 1.170 2.480 ;
        RECT  0.710 1.490 1.050 1.890 ;
    END
END PUI

MACRO QDBHN
    CLASS CORE ;
    FOREIGN QDBHN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.410 0.450 2.500 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.840 2.930 2.870 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 1.130 7.270 3.190 ;
        RECT  6.960 2.790 7.270 3.190 ;
        RECT  6.960 1.490 7.270 1.890 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.270 -0.380 2.670 0.560 ;
        RECT  5.620 -0.380 6.020 0.560 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  1.480 -0.380 1.880 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.270 4.470 2.670 5.420 ;
        RECT  5.870 4.480 6.270 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.950 4.470 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.890 4.180 5.630 4.420 ;
        RECT  6.390 2.100 6.630 4.230 ;
        RECT  5.390 3.990 6.630 4.230 ;
        RECT  3.890 1.390 4.130 4.420 ;
        RECT  5.580 1.490 5.820 3.190 ;
        RECT  5.390 2.100 5.820 2.500 ;
        RECT  4.730 3.700 5.150 3.940 ;
        RECT  4.910 0.620 5.150 3.940 ;
        RECT  0.160 3.870 2.140 4.110 ;
        RECT  0.780 0.670 1.020 4.110 ;
        RECT  4.430 0.800 4.670 3.190 ;
        RECT  0.780 0.800 4.670 1.040 ;
        RECT  0.300 0.670 1.020 0.910 ;
        RECT  3.320 0.770 3.720 1.040 ;
        RECT  2.670 3.990 3.650 4.230 ;
        RECT  2.670 3.390 2.910 4.230 ;
        RECT  1.660 3.390 2.910 3.630 ;
        RECT  1.660 1.390 1.900 3.630 ;
        RECT  3.170 1.390 3.410 3.190 ;
    END
END QDBHN

MACRO QDBHS
    CLASS CORE ;
    FOREIGN QDBHS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.410 0.450 2.500 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.840 2.930 2.870 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 0.990 7.270 3.190 ;
        RECT  6.960 2.790 7.270 3.190 ;
        RECT  6.960 1.490 7.270 1.890 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 -0.380 2.700 0.560 ;
        RECT  5.740 -0.380 6.140 0.560 ;
        RECT  6.820 -0.380 7.220 0.560 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  1.480 -0.380 1.880 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 4.470 2.700 5.420 ;
        RECT  6.010 4.480 6.410 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.950 4.470 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.890 4.180 5.770 4.420 ;
        RECT  6.390 2.100 6.630 4.230 ;
        RECT  5.530 3.990 6.630 4.230 ;
        RECT  3.890 1.390 4.130 4.420 ;
        RECT  5.580 1.490 5.820 3.190 ;
        RECT  5.390 2.100 5.820 2.500 ;
        RECT  4.730 3.700 5.150 3.940 ;
        RECT  4.910 0.620 5.150 3.940 ;
        RECT  0.160 3.870 1.810 4.110 ;
        RECT  0.780 0.670 1.020 4.110 ;
        RECT  4.430 0.800 4.670 3.190 ;
        RECT  0.780 0.800 4.670 1.040 ;
        RECT  0.300 0.670 1.020 0.910 ;
        RECT  2.050 3.990 3.650 4.230 ;
        RECT  2.050 3.390 2.290 4.230 ;
        RECT  1.260 3.390 2.290 3.630 ;
        RECT  1.260 1.390 1.500 3.630 ;
        RECT  3.170 1.390 3.410 3.190 ;
    END
END QDBHS

MACRO QDFFN
    CLASS CORE ;
    FOREIGN QDFFN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.540 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.970 2.230 2.310 2.630 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.660 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.360 0.620 9.640 1.540 ;
        RECT  9.470 1.260 9.750 3.200 ;
        RECT  9.240 2.800 9.750 3.200 ;
        RECT  9.240 0.620 9.640 1.020 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.310 -0.380 2.710 0.560 ;
        RECT  7.890 -0.380 8.130 0.640 ;
        RECT  9.880 -0.380 10.280 0.940 ;
        RECT  0.000 -0.380 10.540 0.380 ;
        RECT  0.910 -0.380 1.310 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 4.040 2.780 5.420 ;
        RECT  5.970 4.480 6.370 5.420 ;
        RECT  7.680 4.480 8.080 5.420 ;
        RECT  9.880 4.260 10.280 5.420 ;
        RECT  0.000 4.660 10.540 5.420 ;
        RECT  0.190 4.260 0.590 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.650 3.850 9.050 4.090 ;
        RECT  8.730 1.370 8.970 4.090 ;
        RECT  7.890 2.480 8.970 2.720 ;
        RECT  7.360 0.890 8.820 1.130 ;
        RECT  8.420 0.730 8.820 1.130 ;
        RECT  4.800 0.620 5.040 1.020 ;
        RECT  7.360 0.620 7.600 1.130 ;
        RECT  4.800 0.620 7.600 0.860 ;
        RECT  4.720 4.000 8.380 4.240 ;
        RECT  8.140 3.080 8.380 4.240 ;
        RECT  4.000 3.520 4.240 4.160 ;
        RECT  4.000 3.520 7.780 3.760 ;
        RECT  7.410 1.660 7.650 3.760 ;
        RECT  4.320 0.620 4.560 3.760 ;
        RECT  7.350 1.660 7.650 2.060 ;
        RECT  3.810 0.620 4.560 0.860 ;
        RECT  5.790 3.040 7.110 3.280 ;
        RECT  6.870 1.100 7.110 3.280 ;
        RECT  5.790 2.120 6.030 3.280 ;
        RECT  5.630 2.120 6.030 2.360 ;
        RECT  6.560 1.100 7.110 1.340 ;
        RECT  4.800 1.500 5.040 3.200 ;
        RECT  6.290 2.260 6.630 2.660 ;
        RECT  6.290 1.580 6.530 2.660 ;
        RECT  4.800 1.580 6.530 1.820 ;
        RECT  0.940 3.240 1.230 3.640 ;
        RECT  0.940 1.100 1.180 3.640 ;
        RECT  3.840 1.100 4.080 3.200 ;
        RECT  0.190 1.100 4.080 1.340 ;
        RECT  3.180 1.580 3.420 4.360 ;
        RECT  3.040 1.580 3.440 1.820 ;
        RECT  1.660 4.040 2.130 4.280 ;
        RECT  1.890 3.560 2.130 4.280 ;
        RECT  1.890 3.560 2.930 3.800 ;
        RECT  2.550 3.400 2.930 3.800 ;
        RECT  2.550 1.580 2.790 3.800 ;
        RECT  1.660 1.580 2.790 1.820 ;
    END
END QDFFN

MACRO QDFFP
    CLASS CORE ;
    FOREIGN QDFFP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.230 1.930 2.630 ;
        RECT  1.410 2.120 1.690 2.840 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.550 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.650 1.280 11.280 1.520 ;
        RECT  10.650 2.960 11.280 3.200 ;
        RECT  10.650 1.280 11.050 3.200 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.040 -0.380 2.440 0.560 ;
        RECT  6.190 -0.380 6.590 0.860 ;
        RECT  9.100 -0.380 9.500 0.560 ;
        RECT  10.160 -0.380 10.560 0.800 ;
        RECT  11.600 -0.380 12.000 0.800 ;
        RECT  0.000 -0.380 12.400 0.380 ;
        RECT  0.880 -0.380 1.280 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.110 4.180 2.510 5.420 ;
        RECT  6.190 4.200 6.590 5.420 ;
        RECT  9.250 4.400 9.490 5.420 ;
        RECT  10.160 4.260 10.560 5.420 ;
        RECT  11.600 4.260 12.000 5.420 ;
        RECT  0.000 4.660 12.400 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.410 4.180 9.010 4.420 ;
        RECT  8.770 3.720 9.010 4.420 ;
        RECT  4.050 4.180 5.410 4.420 ;
        RECT  5.170 3.720 5.410 4.420 ;
        RECT  7.410 3.720 7.650 4.420 ;
        RECT  4.050 0.620 4.290 4.420 ;
        RECT  8.770 3.720 9.920 3.960 ;
        RECT  9.680 1.320 9.920 3.960 ;
        RECT  5.170 3.720 7.650 3.960 ;
        RECT  3.600 3.700 4.290 3.940 ;
        RECT  9.680 2.790 9.970 3.190 ;
        RECT  9.680 1.320 9.970 1.720 ;
        RECT  3.540 0.620 4.290 0.860 ;
        RECT  8.290 3.200 8.530 3.940 ;
        RECT  8.290 3.200 9.420 3.440 ;
        RECT  9.180 0.800 9.420 3.440 ;
        RECT  9.180 2.160 9.440 2.560 ;
        RECT  8.290 0.720 8.530 1.120 ;
        RECT  8.290 0.800 9.420 1.040 ;
        RECT  4.530 3.700 4.930 3.940 ;
        RECT  4.530 0.620 4.770 3.940 ;
        RECT  7.780 1.100 8.020 3.200 ;
        RECT  7.780 2.210 8.600 2.450 ;
        RECT  5.560 1.100 8.020 1.340 ;
        RECT  5.560 0.620 5.800 1.340 ;
        RECT  4.530 0.620 5.800 0.860 ;
        RECT  5.960 2.880 7.540 3.120 ;
        RECT  7.300 1.580 7.540 3.120 ;
        RECT  5.960 2.260 6.200 3.120 ;
        RECT  6.980 1.580 7.540 1.820 ;
        RECT  5.010 1.500 5.250 3.200 ;
        RECT  6.500 2.170 6.980 2.570 ;
        RECT  6.500 1.730 6.740 2.570 ;
        RECT  5.010 1.730 6.740 1.970 ;
        RECT  0.880 3.380 1.200 3.780 ;
        RECT  0.880 1.100 1.120 3.780 ;
        RECT  3.570 1.100 3.810 3.200 ;
        RECT  0.320 1.100 3.810 1.340 ;
        RECT  0.320 0.640 0.560 1.340 ;
        RECT  0.160 0.640 0.560 0.880 ;
        RECT  2.830 4.180 3.230 4.420 ;
        RECT  2.910 1.580 3.150 4.420 ;
        RECT  2.770 1.580 3.170 1.820 ;
        RECT  1.390 4.180 1.790 4.420 ;
        RECT  1.550 3.700 1.790 4.420 ;
        RECT  1.550 3.700 2.520 3.940 ;
        RECT  2.280 1.580 2.520 3.940 ;
        RECT  2.280 3.220 2.660 3.620 ;
        RECT  1.390 1.580 2.520 1.820 ;
    END
END QDFFP

MACRO QDFFRBN
    CLASS CORE ;
    FOREIGN QDFFRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.140 8.610 2.540 ;
        RECT  8.230 1.930 8.510 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.140 1.080 2.540 ;
        RECT  0.790 2.120 1.070 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 1.300 11.610 3.400 ;
        RECT  11.280 3.000 11.610 3.400 ;
        RECT  11.280 1.300 11.610 1.700 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  8.250 -0.380 8.650 0.560 ;
        RECT  10.480 -0.380 10.880 0.860 ;
        RECT  0.000 -0.380 11.780 0.380 ;
        RECT  1.100 -0.380 2.790 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.670 4.020 3.070 5.420 ;
        RECT  8.080 4.480 8.480 5.420 ;
        RECT  10.110 4.130 10.510 5.420 ;
        RECT  0.000 4.660 11.780 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.460 4.180 5.900 4.420 ;
        RECT  5.660 3.580 5.900 4.420 ;
        RECT  4.460 0.620 4.700 4.420 ;
        RECT  4.380 3.620 4.700 4.020 ;
        RECT  5.660 3.580 9.000 3.820 ;
        RECT  8.760 2.880 9.000 3.820 ;
        RECT  8.760 2.880 10.960 3.120 ;
        RECT  10.720 1.100 10.960 3.120 ;
        RECT  9.920 1.100 10.960 1.340 ;
        RECT  9.920 0.620 10.160 1.340 ;
        RECT  9.760 0.620 10.160 0.860 ;
        RECT  4.300 0.620 4.700 0.860 ;
        RECT  10.240 1.640 10.480 2.540 ;
        RECT  9.660 1.640 10.480 1.880 ;
        RECT  9.660 1.580 10.060 1.880 ;
        RECT  9.010 4.090 9.530 4.330 ;
        RECT  9.290 3.420 9.530 4.330 ;
        RECT  9.290 3.420 10.460 3.660 ;
        RECT  4.940 3.700 5.420 3.940 ;
        RECT  4.940 1.100 5.180 3.940 ;
        RECT  8.980 2.120 9.830 2.360 ;
        RECT  8.980 1.120 9.220 2.360 ;
        RECT  6.830 1.120 9.220 1.360 ;
        RECT  4.940 1.100 7.070 1.340 ;
        RECT  5.310 0.860 5.710 1.340 ;
        RECT  7.580 0.620 7.980 0.880 ;
        RECT  6.180 0.620 7.980 0.860 ;
        RECT  7.730 1.600 7.970 3.220 ;
        RECT  6.140 2.880 7.970 3.120 ;
        RECT  6.140 1.600 7.970 1.840 ;
        RECT  6.140 1.580 6.540 1.840 ;
        RECT  6.190 4.160 7.820 4.400 ;
        RECT  5.420 2.880 5.820 3.120 ;
        RECT  5.500 1.580 5.740 3.120 ;
        RECT  5.500 2.220 6.820 2.460 ;
        RECT  5.420 1.580 5.820 1.820 ;
        RECT  3.980 1.290 4.220 3.200 ;
        RECT  0.190 2.800 0.480 3.200 ;
        RECT  0.190 1.010 0.430 3.200 ;
        RECT  3.840 1.010 4.080 1.530 ;
        RECT  0.160 1.010 4.080 1.250 ;
        RECT  3.390 4.020 3.790 4.260 ;
        RECT  3.390 3.430 3.630 4.260 ;
        RECT  3.260 1.580 3.500 3.670 ;
        RECT  3.260 2.260 3.690 2.660 ;
        RECT  3.180 1.580 3.580 1.820 ;
        RECT  1.740 3.540 2.940 3.780 ;
        RECT  2.700 1.580 2.940 3.780 ;
        RECT  2.700 2.260 3.010 2.660 ;
        RECT  1.740 1.580 2.940 1.820 ;
    END
END QDFFRBN

MACRO QDFFRBP
    CLASS CORE ;
    FOREIGN QDFFRBP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.930 8.510 2.650 ;
        RECT  8.010 2.140 8.510 2.540 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.230 1.930 2.630 ;
        RECT  1.410 2.120 1.690 2.840 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.530 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 1.260 11.610 3.220 ;
        RECT  11.120 2.940 11.610 3.220 ;
        RECT  11.120 1.260 11.610 1.540 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  7.820 -0.380 8.220 0.560 ;
        RECT  10.400 -0.380 10.800 0.860 ;
        RECT  11.840 -0.380 12.240 0.860 ;
        RECT  0.000 -0.380 12.400 0.380 ;
        RECT  1.090 -0.380 2.440 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.310 4.020 2.710 5.420 ;
        RECT  7.720 4.480 8.120 5.420 ;
        RECT  9.380 4.480 9.780 5.420 ;
        RECT  10.190 4.480 10.590 5.420 ;
        RECT  11.840 4.260 12.240 5.420 ;
        RECT  0.000 4.660 12.400 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.100 4.180 5.540 4.420 ;
        RECT  5.300 3.580 5.540 4.420 ;
        RECT  4.100 0.620 4.340 4.420 ;
        RECT  4.020 3.620 4.340 4.020 ;
        RECT  5.300 3.580 10.880 3.820 ;
        RECT  10.640 1.100 10.880 3.820 ;
        RECT  9.840 1.100 10.880 1.340 ;
        RECT  9.840 0.620 10.080 1.340 ;
        RECT  9.680 0.620 10.080 0.860 ;
        RECT  3.940 0.620 4.340 0.860 ;
        RECT  8.590 3.100 10.400 3.340 ;
        RECT  10.160 1.650 10.400 3.340 ;
        RECT  9.250 1.650 10.400 1.890 ;
        RECT  9.250 1.490 9.490 1.890 ;
        RECT  4.580 3.700 5.060 3.940 ;
        RECT  4.580 1.100 4.820 3.940 ;
        RECT  8.770 2.220 9.410 2.460 ;
        RECT  8.770 1.120 9.010 2.460 ;
        RECT  6.470 1.120 9.010 1.360 ;
        RECT  4.580 1.100 6.710 1.340 ;
        RECT  4.950 0.860 5.350 1.340 ;
        RECT  7.370 1.600 7.610 3.220 ;
        RECT  5.780 2.880 7.610 3.120 ;
        RECT  5.780 1.600 7.610 1.840 ;
        RECT  5.780 1.580 6.180 1.840 ;
        RECT  7.150 0.620 7.550 0.880 ;
        RECT  5.820 0.620 7.550 0.860 ;
        RECT  5.830 4.160 7.460 4.400 ;
        RECT  5.060 2.880 5.460 3.120 ;
        RECT  5.140 1.580 5.380 3.120 ;
        RECT  5.140 2.220 6.460 2.460 ;
        RECT  5.060 1.580 5.460 1.820 ;
        RECT  0.820 3.130 1.200 3.530 ;
        RECT  3.620 1.290 3.860 3.200 ;
        RECT  0.820 1.010 1.060 3.530 ;
        RECT  3.480 1.010 3.720 1.530 ;
        RECT  0.160 1.010 3.720 1.250 ;
        RECT  3.110 3.370 3.350 4.340 ;
        RECT  2.910 1.570 3.150 3.610 ;
        RECT  2.910 2.260 3.340 2.660 ;
        RECT  2.820 1.570 3.220 1.810 ;
        RECT  1.520 3.930 1.920 4.170 ;
        RECT  1.680 3.540 1.920 4.170 ;
        RECT  1.680 3.540 2.580 3.780 ;
        RECT  2.340 1.570 2.580 3.780 ;
        RECT  2.340 2.260 2.660 2.660 ;
        RECT  1.390 1.570 2.580 1.810 ;
    END
END QDFFRBP

MACRO QDFFRBS
    CLASS CORE ;
    FOREIGN QDFFRBS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.140 8.590 2.540 ;
        RECT  8.230 1.930 8.510 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.140 1.080 2.540 ;
        RECT  0.790 2.120 1.070 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 0.650 11.610 3.400 ;
        RECT  11.280 3.000 11.610 3.400 ;
        RECT  11.280 0.650 11.610 1.050 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  8.230 -0.380 8.630 0.560 ;
        RECT  10.460 -0.380 10.860 0.860 ;
        RECT  0.000 -0.380 11.780 0.380 ;
        RECT  1.100 -0.380 2.790 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.670 4.020 3.070 5.420 ;
        RECT  8.060 4.480 8.460 5.420 ;
        RECT  10.090 4.130 10.490 5.420 ;
        RECT  0.000 4.660 11.780 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.440 4.180 5.880 4.420 ;
        RECT  5.640 3.580 5.880 4.420 ;
        RECT  4.440 0.620 4.680 4.420 ;
        RECT  4.360 3.620 4.680 4.020 ;
        RECT  5.640 3.580 8.980 3.820 ;
        RECT  8.740 2.880 8.980 3.820 ;
        RECT  8.740 2.880 10.940 3.120 ;
        RECT  10.700 1.100 10.940 3.120 ;
        RECT  9.900 1.100 10.940 1.340 ;
        RECT  9.900 0.620 10.140 1.340 ;
        RECT  9.740 0.620 10.140 0.860 ;
        RECT  4.280 0.620 4.680 0.860 ;
        RECT  10.220 1.640 10.460 2.540 ;
        RECT  9.640 1.640 10.460 1.880 ;
        RECT  9.640 1.580 10.040 1.880 ;
        RECT  8.990 4.090 9.510 4.330 ;
        RECT  9.270 3.420 9.510 4.330 ;
        RECT  9.270 3.420 10.440 3.660 ;
        RECT  4.920 3.700 5.400 3.940 ;
        RECT  4.920 1.100 5.160 3.940 ;
        RECT  8.960 2.120 9.810 2.360 ;
        RECT  8.960 1.120 9.200 2.360 ;
        RECT  6.810 1.120 9.200 1.360 ;
        RECT  4.920 1.100 7.050 1.340 ;
        RECT  5.290 0.860 5.690 1.340 ;
        RECT  7.560 0.620 7.960 0.880 ;
        RECT  6.160 0.620 7.960 0.860 ;
        RECT  7.710 1.600 7.950 3.220 ;
        RECT  6.120 2.880 7.950 3.120 ;
        RECT  6.120 1.600 7.950 1.840 ;
        RECT  6.120 1.580 6.520 1.840 ;
        RECT  6.170 4.160 7.800 4.400 ;
        RECT  5.400 2.880 5.800 3.120 ;
        RECT  5.480 1.580 5.720 3.120 ;
        RECT  5.480 2.220 6.800 2.460 ;
        RECT  5.400 1.580 5.800 1.820 ;
        RECT  3.960 1.290 4.200 3.200 ;
        RECT  0.190 2.800 0.480 3.200 ;
        RECT  0.190 1.010 0.430 3.200 ;
        RECT  3.820 1.010 4.060 1.530 ;
        RECT  0.160 1.010 4.060 1.250 ;
        RECT  3.370 4.020 3.790 4.260 ;
        RECT  3.370 3.430 3.610 4.260 ;
        RECT  3.240 1.580 3.480 3.670 ;
        RECT  3.240 2.260 3.690 2.660 ;
        RECT  3.160 1.580 3.560 1.820 ;
        RECT  1.740 3.540 2.920 3.780 ;
        RECT  2.680 1.580 2.920 3.780 ;
        RECT  2.680 2.260 2.990 2.660 ;
        RECT  1.740 1.580 2.920 1.820 ;
    END
END QDFFRBS

MACRO QDFFRBT
    CLASS CORE ;
    FOREIGN QDFFRBT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.640 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 1.930 8.510 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.910 2.230 2.310 2.630 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.470 2.820 11.710 3.220 ;
        RECT  11.470 1.260 13.230 1.540 ;
        RECT  12.510 1.260 12.910 3.220 ;
        RECT  12.510 1.260 13.230 1.580 ;
        RECT  11.470 2.940 13.230 3.220 ;
        RECT  11.470 1.260 11.710 1.660 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.250 -0.380 2.650 0.560 ;
        RECT  8.090 -0.380 8.490 0.560 ;
        RECT  10.670 -0.380 11.070 0.860 ;
        RECT  12.110 -0.380 12.510 0.860 ;
        RECT  0.000 -0.380 13.640 0.380 ;
        RECT  1.200 -0.380 1.600 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.020 2.720 5.420 ;
        RECT  8.070 4.480 8.470 5.420 ;
        RECT  9.650 4.480 10.050 5.420 ;
        RECT  10.470 4.480 10.870 5.420 ;
        RECT  12.110 4.260 12.510 5.420 ;
        RECT  0.000 4.660 13.640 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.320 4.180 5.760 4.420 ;
        RECT  5.520 3.580 5.760 4.420 ;
        RECT  4.320 0.620 4.560 4.420 ;
        RECT  4.240 3.620 4.560 4.020 ;
        RECT  5.520 3.580 11.230 3.820 ;
        RECT  10.990 1.100 11.230 3.820 ;
        RECT  10.110 1.100 11.230 1.340 ;
        RECT  10.110 0.620 10.350 1.340 ;
        RECT  9.950 0.620 10.350 0.860 ;
        RECT  4.160 0.620 4.560 0.860 ;
        RECT  8.860 3.100 10.750 3.340 ;
        RECT  10.510 1.640 10.750 3.340 ;
        RECT  9.440 1.640 10.750 1.880 ;
        RECT  9.440 1.570 9.840 1.880 ;
        RECT  4.800 3.700 5.280 3.940 ;
        RECT  4.800 1.100 5.040 3.940 ;
        RECT  8.840 2.220 9.690 2.460 ;
        RECT  8.840 1.120 9.080 2.460 ;
        RECT  6.690 1.120 9.080 1.360 ;
        RECT  4.800 1.100 6.930 1.340 ;
        RECT  5.170 0.860 5.570 1.340 ;
        RECT  7.590 2.820 7.830 3.220 ;
        RECT  6.000 2.880 7.830 3.120 ;
        RECT  7.510 1.600 7.750 3.120 ;
        RECT  6.000 1.600 7.750 1.840 ;
        RECT  6.000 1.580 6.400 1.840 ;
        RECT  7.350 0.620 7.750 0.880 ;
        RECT  6.040 0.620 7.750 0.860 ;
        RECT  6.050 4.160 7.680 4.400 ;
        RECT  5.280 2.880 5.680 3.120 ;
        RECT  5.360 1.580 5.600 3.120 ;
        RECT  5.360 2.220 6.680 2.460 ;
        RECT  5.280 1.580 5.680 1.820 ;
        RECT  3.840 1.290 4.080 3.200 ;
        RECT  0.960 1.020 1.200 3.190 ;
        RECT  3.700 1.020 3.940 1.530 ;
        RECT  0.160 1.020 3.940 1.260 ;
        RECT  3.120 1.580 3.360 4.340 ;
        RECT  3.120 2.260 3.550 2.660 ;
        RECT  3.040 1.580 3.440 1.820 ;
        RECT  1.530 3.930 1.930 4.170 ;
        RECT  1.690 3.540 1.930 4.170 ;
        RECT  1.690 3.540 2.800 3.780 ;
        RECT  2.560 1.580 2.800 3.780 ;
        RECT  2.560 2.260 2.870 2.660 ;
        RECT  1.600 1.580 2.800 1.820 ;
    END
END QDFFRBT

MACRO QDFFRSBN
    CLASS CORE ;
    FOREIGN QDFFRSBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.640 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.370 3.210 ;
        RECT  9.690 2.140 10.370 2.540 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.300 13.470 3.400 ;
        RECT  13.160 3.000 13.470 3.400 ;
        RECT  13.160 1.300 13.470 1.700 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.090 1.620 9.330 2.450 ;
        RECT  7.360 2.210 9.330 2.450 ;
        RECT  10.090 1.100 10.330 1.860 ;
        RECT  9.090 1.620 10.330 1.860 ;
        RECT  10.090 1.100 11.610 1.340 ;
        RECT  11.330 1.100 11.610 2.210 ;
        RECT  7.360 2.140 7.600 2.540 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 -0.380 2.780 0.560 ;
        RECT  8.970 -0.380 9.370 0.560 ;
        RECT  12.360 -0.380 12.760 0.860 ;
        RECT  0.000 -0.380 13.640 0.380 ;
        RECT  1.410 -0.380 1.810 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 4.030 2.920 5.420 ;
        RECT  9.400 4.480 9.800 5.420 ;
        RECT  12.120 4.130 12.520 5.420 ;
        RECT  0.000 4.660 13.640 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.450 4.180 5.890 4.420 ;
        RECT  5.650 3.580 5.890 4.420 ;
        RECT  4.450 0.620 4.690 4.420 ;
        RECT  4.370 3.620 4.690 4.020 ;
        RECT  8.420 3.580 10.910 3.820 ;
        RECT  10.670 2.940 10.910 3.820 ;
        RECT  5.650 3.580 7.290 3.820 ;
        RECT  7.050 3.360 8.660 3.600 ;
        RECT  10.670 2.940 12.920 3.180 ;
        RECT  12.680 1.100 12.920 3.180 ;
        RECT  11.880 1.100 12.920 1.340 ;
        RECT  11.880 0.620 12.120 1.340 ;
        RECT  11.080 0.620 12.120 0.860 ;
        RECT  4.290 0.620 4.690 0.860 ;
        RECT  10.720 2.450 12.440 2.690 ;
        RECT  12.200 2.140 12.440 2.690 ;
        RECT  10.720 1.580 10.960 2.690 ;
        RECT  10.570 1.580 10.970 1.820 ;
        RECT  10.330 4.090 11.390 4.330 ;
        RECT  11.150 3.480 11.390 4.330 ;
        RECT  11.150 3.480 12.340 3.720 ;
        RECT  4.930 3.700 5.410 3.940 ;
        RECT  4.930 1.100 5.170 3.940 ;
        RECT  6.820 1.120 9.850 1.360 ;
        RECT  9.610 0.620 9.850 1.360 ;
        RECT  4.930 1.100 7.060 1.340 ;
        RECT  5.300 0.860 5.700 1.340 ;
        RECT  9.610 0.620 10.700 0.860 ;
        RECT  9.050 2.820 9.290 3.220 ;
        RECT  6.130 2.880 9.290 3.120 ;
        RECT  6.880 1.600 7.120 3.120 ;
        RECT  6.130 1.600 8.650 1.840 ;
        RECT  6.130 1.580 6.530 1.840 ;
        RECT  6.180 4.160 9.140 4.400 ;
        RECT  7.660 3.840 8.060 4.400 ;
        RECT  8.330 0.620 8.730 0.880 ;
        RECT  6.170 0.620 8.730 0.860 ;
        RECT  5.410 2.880 5.810 3.120 ;
        RECT  5.490 1.580 5.730 3.120 ;
        RECT  6.400 2.140 6.640 2.540 ;
        RECT  5.490 2.220 6.640 2.460 ;
        RECT  5.410 1.580 5.810 1.820 ;
        RECT  3.970 1.290 4.210 3.200 ;
        RECT  0.960 1.010 1.200 3.190 ;
        RECT  3.830 1.010 4.070 1.530 ;
        RECT  0.160 1.010 4.070 1.250 ;
        RECT  3.250 3.950 3.560 4.350 ;
        RECT  3.250 1.580 3.490 4.350 ;
        RECT  3.250 2.260 3.680 2.660 ;
        RECT  3.170 1.580 3.570 1.820 ;
        RECT  1.730 3.930 2.130 4.170 ;
        RECT  1.890 3.540 2.130 4.170 ;
        RECT  1.890 3.540 2.930 3.780 ;
        RECT  2.690 1.580 2.930 3.780 ;
        RECT  2.690 2.260 3.000 2.660 ;
        RECT  1.730 1.580 2.930 1.820 ;
    END
END QDFFRSBN

MACRO QDFFS
    CLASS CORE ;
    FOREIGN QDFFS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.540 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.970 2.230 2.310 2.630 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.660 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.360 0.620 9.640 1.540 ;
        RECT  9.470 1.260 9.750 3.200 ;
        RECT  9.240 2.800 9.750 3.200 ;
        RECT  9.240 0.620 9.640 1.020 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.310 -0.380 2.710 0.560 ;
        RECT  7.890 -0.380 8.130 0.640 ;
        RECT  9.880 -0.380 10.280 0.940 ;
        RECT  0.000 -0.380 10.540 0.380 ;
        RECT  0.910 -0.380 1.310 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 4.040 2.780 5.420 ;
        RECT  5.970 4.480 6.370 5.420 ;
        RECT  7.680 4.480 8.080 5.420 ;
        RECT  9.880 4.130 10.280 5.420 ;
        RECT  0.000 4.660 10.540 5.420 ;
        RECT  0.190 4.260 0.590 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.650 4.100 9.050 4.340 ;
        RECT  8.730 1.370 8.970 4.340 ;
        RECT  7.890 2.480 8.970 2.720 ;
        RECT  7.360 0.890 8.820 1.130 ;
        RECT  8.420 0.730 8.820 1.130 ;
        RECT  4.800 0.620 5.040 1.020 ;
        RECT  7.360 0.620 7.600 1.130 ;
        RECT  4.800 0.620 7.600 0.860 ;
        RECT  4.720 4.000 8.380 4.240 ;
        RECT  8.140 3.080 8.380 4.240 ;
        RECT  4.000 3.520 4.240 4.160 ;
        RECT  4.000 3.520 7.780 3.760 ;
        RECT  7.410 1.660 7.650 3.760 ;
        RECT  4.320 0.620 4.560 3.760 ;
        RECT  7.350 1.660 7.650 2.060 ;
        RECT  3.810 0.620 4.560 0.860 ;
        RECT  5.790 3.040 7.110 3.280 ;
        RECT  6.870 1.100 7.110 3.280 ;
        RECT  5.790 2.120 6.030 3.280 ;
        RECT  5.630 2.120 6.030 2.360 ;
        RECT  6.560 1.100 7.110 1.340 ;
        RECT  4.800 1.500 5.040 3.200 ;
        RECT  6.290 2.260 6.630 2.660 ;
        RECT  6.290 1.580 6.530 2.660 ;
        RECT  4.800 1.580 6.530 1.820 ;
        RECT  0.940 3.240 1.230 3.640 ;
        RECT  0.940 1.100 1.180 3.640 ;
        RECT  3.840 1.100 4.080 3.200 ;
        RECT  0.190 1.100 4.080 1.340 ;
        RECT  3.180 1.580 3.420 4.360 ;
        RECT  3.040 1.580 3.440 1.820 ;
        RECT  1.660 4.040 2.130 4.280 ;
        RECT  1.890 3.560 2.130 4.280 ;
        RECT  1.890 3.560 2.930 3.800 ;
        RECT  2.550 3.400 2.930 3.800 ;
        RECT  2.550 1.580 2.790 3.800 ;
        RECT  1.660 1.580 2.790 1.820 ;
    END
END QDFFS

MACRO QDFZN
    CLASS CORE ;
    FOREIGN QDFZN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        RECT  3.830 2.230 4.170 2.630 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.220 2.310 2.620 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.220 0.620 11.500 1.540 ;
        RECT  11.330 1.260 11.610 3.200 ;
        RECT  11.100 2.800 11.610 3.200 ;
        RECT  11.100 0.620 11.500 1.020 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.170 -0.380 4.570 0.560 ;
        RECT  9.750 -0.380 9.990 0.640 ;
        RECT  11.740 -0.380 12.140 0.940 ;
        RECT  0.000 -0.380 12.400 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.240 4.020 4.640 5.420 ;
        RECT  7.830 4.480 8.230 5.420 ;
        RECT  9.540 4.480 9.940 5.420 ;
        RECT  11.740 4.260 12.140 5.420 ;
        RECT  0.000 4.660 12.400 5.420 ;
        RECT  2.010 4.480 2.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.590 1.370 10.830 4.170 ;
        RECT  9.750 2.480 10.830 2.720 ;
        RECT  9.220 0.890 10.680 1.130 ;
        RECT  10.280 0.730 10.680 1.130 ;
        RECT  6.660 0.620 6.900 1.020 ;
        RECT  9.220 0.620 9.460 1.130 ;
        RECT  6.660 0.620 9.460 0.860 ;
        RECT  6.580 4.000 10.240 4.240 ;
        RECT  10.000 3.080 10.240 4.240 ;
        RECT  5.860 3.520 6.100 4.160 ;
        RECT  5.860 3.520 9.640 3.760 ;
        RECT  9.270 1.660 9.510 3.760 ;
        RECT  6.180 0.620 6.420 3.760 ;
        RECT  9.210 1.660 9.510 2.060 ;
        RECT  5.670 0.620 6.420 0.860 ;
        RECT  7.650 3.040 8.970 3.280 ;
        RECT  8.730 1.100 8.970 3.280 ;
        RECT  7.650 2.130 7.890 3.280 ;
        RECT  7.490 2.130 7.890 2.370 ;
        RECT  8.420 1.100 8.970 1.340 ;
        RECT  6.660 1.500 6.900 3.200 ;
        RECT  8.150 2.260 8.490 2.660 ;
        RECT  8.150 1.590 8.390 2.660 ;
        RECT  6.660 1.590 8.390 1.830 ;
        RECT  5.700 1.100 5.940 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.040 1.580 5.280 4.340 ;
        RECT  4.900 1.580 5.300 1.820 ;
        RECT  3.520 4.020 3.920 4.260 ;
        RECT  3.680 3.540 3.920 4.260 ;
        RECT  3.680 3.540 4.650 3.780 ;
        RECT  4.410 1.580 4.650 3.780 ;
        RECT  4.410 3.220 4.790 3.620 ;
        RECT  3.520 1.580 4.650 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END QDFZN

MACRO QDFZP
    CLASS CORE ;
    FOREIGN QDFZP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        RECT  3.830 2.230 4.170 2.630 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.220 2.310 2.620 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.130 1.280 13.530 3.200 ;
        RECT  12.970 2.960 13.530 3.200 ;
        RECT  12.970 1.280 13.530 1.520 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.170 -0.380 4.570 0.560 ;
        RECT  8.280 -0.380 8.680 0.860 ;
        RECT  11.190 -0.380 11.590 0.560 ;
        RECT  12.250 -0.380 12.650 0.800 ;
        RECT  13.690 -0.380 14.090 0.800 ;
        RECT  0.000 -0.380 14.260 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.240 4.020 4.640 5.420 ;
        RECT  8.280 4.200 8.680 5.420 ;
        RECT  11.340 4.400 11.580 5.420 ;
        RECT  12.250 4.260 12.650 5.420 ;
        RECT  13.690 4.260 14.090 5.420 ;
        RECT  0.000 4.660 14.260 5.420 ;
        RECT  2.010 4.480 2.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.500 4.180 11.100 4.420 ;
        RECT  10.860 3.720 11.100 4.420 ;
        RECT  6.180 4.180 7.540 4.420 ;
        RECT  7.300 3.720 7.540 4.420 ;
        RECT  9.500 3.720 9.740 4.420 ;
        RECT  6.180 0.620 6.420 4.420 ;
        RECT  10.860 3.720 12.010 3.960 ;
        RECT  11.770 1.320 12.010 3.960 ;
        RECT  7.300 3.720 9.740 3.960 ;
        RECT  5.730 3.700 6.420 3.940 ;
        RECT  11.770 2.790 12.060 3.190 ;
        RECT  11.770 1.320 12.060 1.720 ;
        RECT  5.670 0.620 6.420 0.860 ;
        RECT  10.380 3.200 10.620 3.940 ;
        RECT  10.380 3.200 11.510 3.440 ;
        RECT  11.270 0.800 11.510 3.440 ;
        RECT  11.270 2.160 11.530 2.560 ;
        RECT  10.380 0.720 10.620 1.120 ;
        RECT  10.380 0.800 11.510 1.040 ;
        RECT  6.660 3.700 7.060 3.940 ;
        RECT  6.660 0.620 6.900 3.940 ;
        RECT  9.870 1.100 10.110 3.200 ;
        RECT  9.870 2.210 10.690 2.450 ;
        RECT  7.690 1.100 10.110 1.340 ;
        RECT  7.690 0.620 7.930 1.340 ;
        RECT  6.660 0.620 7.930 0.860 ;
        RECT  8.050 2.880 9.630 3.120 ;
        RECT  9.390 1.580 9.630 3.120 ;
        RECT  8.050 2.260 8.290 3.120 ;
        RECT  9.070 1.580 9.630 1.820 ;
        RECT  7.140 1.500 7.380 3.200 ;
        RECT  8.590 2.170 9.070 2.570 ;
        RECT  8.590 1.730 8.830 2.570 ;
        RECT  7.140 1.730 8.830 1.970 ;
        RECT  5.700 1.100 5.940 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.040 1.580 5.280 4.340 ;
        RECT  4.900 1.580 5.300 1.820 ;
        RECT  3.520 4.020 3.920 4.260 ;
        RECT  3.680 3.520 3.920 4.260 ;
        RECT  3.680 3.520 4.650 3.760 ;
        RECT  4.410 1.580 4.650 3.760 ;
        RECT  4.410 3.220 4.790 3.620 ;
        RECT  3.520 1.580 4.650 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END QDFZP

MACRO QDFZRBN
    CLASS CORE ;
    FOREIGN QDFZRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.640 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.470 2.540 ;
        RECT  10.090 1.930 10.370 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.270 2.310 2.670 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.200 13.470 3.840 ;
        RECT  13.140 3.440 13.470 3.840 ;
        RECT  13.140 1.200 13.470 1.600 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.380 4.650 0.560 ;
        RECT  10.110 -0.380 10.510 0.560 ;
        RECT  12.340 -0.380 12.740 0.860 ;
        RECT  0.000 -0.380 13.640 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 4.030 4.720 5.420 ;
        RECT  9.940 4.480 10.340 5.420 ;
        RECT  11.970 4.130 12.370 5.420 ;
        RECT  0.000 4.660 13.640 5.420 ;
        RECT  2.090 4.480 2.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 4.180 7.760 4.420 ;
        RECT  7.520 3.580 7.760 4.420 ;
        RECT  6.320 0.620 6.560 4.420 ;
        RECT  6.240 3.620 6.560 4.020 ;
        RECT  7.520 3.580 10.860 3.820 ;
        RECT  10.620 2.880 10.860 3.820 ;
        RECT  10.620 2.880 12.820 3.120 ;
        RECT  12.580 1.100 12.820 3.120 ;
        RECT  11.780 1.100 12.820 1.340 ;
        RECT  11.780 0.620 12.020 1.340 ;
        RECT  11.620 0.620 12.020 0.860 ;
        RECT  6.160 0.620 6.560 0.860 ;
        RECT  12.100 1.640 12.340 2.540 ;
        RECT  11.520 1.640 12.340 1.880 ;
        RECT  11.520 1.580 11.920 1.880 ;
        RECT  10.870 4.090 11.390 4.330 ;
        RECT  11.150 3.420 11.390 4.330 ;
        RECT  11.150 3.420 12.320 3.660 ;
        RECT  6.800 3.700 7.280 3.940 ;
        RECT  6.800 1.100 7.040 3.940 ;
        RECT  10.840 2.120 11.690 2.360 ;
        RECT  10.840 1.120 11.080 2.360 ;
        RECT  8.690 1.120 11.080 1.360 ;
        RECT  6.800 1.100 8.930 1.340 ;
        RECT  7.170 0.860 7.570 1.340 ;
        RECT  9.440 0.620 9.840 0.880 ;
        RECT  8.040 0.620 9.840 0.860 ;
        RECT  9.590 1.600 9.830 3.220 ;
        RECT  8.000 2.880 9.830 3.120 ;
        RECT  8.000 1.600 9.830 1.840 ;
        RECT  8.000 1.580 8.400 1.840 ;
        RECT  8.050 4.160 9.680 4.400 ;
        RECT  7.280 2.880 7.680 3.120 ;
        RECT  7.360 1.580 7.600 3.120 ;
        RECT  7.360 2.220 8.680 2.460 ;
        RECT  7.280 1.580 7.680 1.820 ;
        RECT  5.840 1.290 6.080 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.700 1.290 6.080 1.530 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.120 1.580 5.360 4.350 ;
        RECT  5.120 2.260 5.550 2.660 ;
        RECT  5.040 1.580 5.440 1.820 ;
        RECT  3.600 4.030 4.000 4.270 ;
        RECT  3.760 3.540 4.000 4.270 ;
        RECT  3.760 3.540 4.800 3.780 ;
        RECT  4.560 1.580 4.800 3.780 ;
        RECT  4.560 2.260 4.870 2.660 ;
        RECT  3.600 1.580 4.800 1.820 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.280 3.700 ;
        RECT  2.880 3.940 3.280 4.420 ;
        RECT  1.230 3.940 3.280 4.180 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
    END
END QDFZRBN

MACRO QDFZRBP
    CLASS CORE ;
    FOREIGN QDFZRBP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.470 2.540 ;
        RECT  10.090 1.930 10.370 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.270 2.310 2.670 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 1.260 14.090 3.780 ;
        RECT  13.470 3.500 14.090 3.780 ;
        RECT  13.470 1.260 14.090 1.540 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.380 4.650 0.560 ;
        RECT  10.110 -0.380 10.510 0.560 ;
        RECT  12.750 -0.380 13.150 0.860 ;
        RECT  14.190 -0.380 14.590 0.860 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 4.020 4.720 5.420 ;
        RECT  9.940 4.480 10.340 5.420 ;
        RECT  11.660 4.480 12.060 5.420 ;
        RECT  12.470 4.480 12.870 5.420 ;
        RECT  14.190 4.260 14.590 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  2.090 4.480 2.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 4.180 7.760 4.420 ;
        RECT  7.520 3.580 7.760 4.420 ;
        RECT  6.320 0.620 6.560 4.420 ;
        RECT  6.240 3.620 6.560 4.020 ;
        RECT  7.520 3.580 13.230 3.820 ;
        RECT  12.990 1.100 13.230 3.820 ;
        RECT  12.190 1.100 13.230 1.340 ;
        RECT  12.190 0.620 12.430 1.340 ;
        RECT  12.030 0.620 12.430 0.860 ;
        RECT  6.160 0.620 6.560 0.860 ;
        RECT  10.870 3.100 12.750 3.340 ;
        RECT  12.510 1.640 12.750 3.340 ;
        RECT  11.520 1.640 12.750 1.880 ;
        RECT  11.520 1.570 11.920 1.880 ;
        RECT  6.800 3.700 7.280 3.940 ;
        RECT  6.800 1.100 7.040 3.940 ;
        RECT  10.840 2.220 11.690 2.460 ;
        RECT  10.840 1.120 11.080 2.460 ;
        RECT  8.690 1.120 11.080 1.360 ;
        RECT  6.800 1.100 8.930 1.340 ;
        RECT  7.170 0.860 7.570 1.340 ;
        RECT  9.440 0.620 9.840 0.880 ;
        RECT  8.040 0.620 9.840 0.860 ;
        RECT  9.590 1.600 9.830 3.220 ;
        RECT  8.000 2.880 9.830 3.120 ;
        RECT  8.000 1.600 9.830 1.840 ;
        RECT  8.000 1.580 8.400 1.840 ;
        RECT  8.050 4.160 9.680 4.400 ;
        RECT  7.280 2.880 7.680 3.120 ;
        RECT  7.360 1.580 7.600 3.120 ;
        RECT  7.360 2.220 8.680 2.460 ;
        RECT  7.280 1.580 7.680 1.820 ;
        RECT  5.840 1.290 6.080 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.700 1.290 6.080 1.530 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.120 1.580 5.360 4.340 ;
        RECT  5.120 2.260 5.550 2.660 ;
        RECT  5.040 1.580 5.440 1.820 ;
        RECT  3.600 4.020 4.000 4.260 ;
        RECT  3.760 3.540 4.000 4.260 ;
        RECT  3.760 3.540 4.800 3.780 ;
        RECT  4.560 1.580 4.800 3.780 ;
        RECT  4.560 2.260 4.870 2.660 ;
        RECT  3.600 1.580 4.800 1.820 ;
        RECT  0.160 4.140 0.990 4.380 ;
        RECT  0.750 3.460 0.990 4.380 ;
        RECT  0.750 3.460 3.280 3.700 ;
        RECT  2.880 3.940 3.280 4.420 ;
        RECT  1.230 3.940 3.280 4.180 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
    END
END QDFZRBP

MACRO QDFZRBS
    CLASS CORE ;
    FOREIGN QDFZRBS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.640 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.470 2.540 ;
        RECT  10.090 1.930 10.370 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.270 2.310 2.670 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 0.750 13.470 3.670 ;
        RECT  13.160 3.270 13.470 3.670 ;
        RECT  13.160 0.750 13.470 1.150 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.380 4.650 0.560 ;
        RECT  10.110 -0.380 10.510 0.560 ;
        RECT  12.340 -0.380 12.740 0.860 ;
        RECT  0.000 -0.380 13.640 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 4.030 4.720 5.420 ;
        RECT  9.940 4.480 10.340 5.420 ;
        RECT  11.970 4.130 12.370 5.420 ;
        RECT  0.000 4.660 13.640 5.420 ;
        RECT  2.090 4.480 2.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 4.180 7.760 4.420 ;
        RECT  7.520 3.580 7.760 4.420 ;
        RECT  6.320 0.620 6.560 4.420 ;
        RECT  6.240 3.620 6.560 4.020 ;
        RECT  7.520 3.580 10.860 3.820 ;
        RECT  10.620 2.880 10.860 3.820 ;
        RECT  10.620 2.880 12.820 3.120 ;
        RECT  12.580 1.100 12.820 3.120 ;
        RECT  11.780 1.100 12.820 1.340 ;
        RECT  11.780 0.620 12.020 1.340 ;
        RECT  11.620 0.620 12.020 0.860 ;
        RECT  6.160 0.620 6.560 0.860 ;
        RECT  12.100 1.640 12.340 2.540 ;
        RECT  11.520 1.640 12.340 1.880 ;
        RECT  11.520 1.580 11.920 1.880 ;
        RECT  10.870 4.090 11.390 4.330 ;
        RECT  11.150 3.420 11.390 4.330 ;
        RECT  11.150 3.420 12.320 3.660 ;
        RECT  6.800 3.700 7.280 3.940 ;
        RECT  6.800 1.100 7.040 3.940 ;
        RECT  10.840 2.120 11.690 2.360 ;
        RECT  10.840 1.120 11.080 2.360 ;
        RECT  8.690 1.120 11.080 1.360 ;
        RECT  6.800 1.100 8.930 1.340 ;
        RECT  7.170 0.860 7.570 1.340 ;
        RECT  9.440 0.620 9.840 0.880 ;
        RECT  8.040 0.620 9.840 0.860 ;
        RECT  9.590 1.600 9.830 3.220 ;
        RECT  8.000 2.880 9.830 3.120 ;
        RECT  8.000 1.600 9.830 1.840 ;
        RECT  8.000 1.580 8.400 1.840 ;
        RECT  8.050 4.160 9.680 4.400 ;
        RECT  7.280 2.880 7.680 3.120 ;
        RECT  7.360 1.580 7.600 3.120 ;
        RECT  7.360 2.220 8.680 2.460 ;
        RECT  7.280 1.580 7.680 1.820 ;
        RECT  5.840 1.290 6.080 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.700 1.290 6.080 1.530 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.120 1.580 5.360 4.350 ;
        RECT  5.120 2.260 5.550 2.660 ;
        RECT  5.040 1.580 5.440 1.820 ;
        RECT  3.600 4.030 4.000 4.270 ;
        RECT  3.760 3.540 4.000 4.270 ;
        RECT  3.760 3.540 4.800 3.780 ;
        RECT  4.560 1.580 4.800 3.780 ;
        RECT  4.560 2.260 4.870 2.660 ;
        RECT  3.600 1.580 4.800 1.820 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.280 3.700 ;
        RECT  2.880 3.940 3.280 4.420 ;
        RECT  1.230 3.940 3.280 4.180 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
    END
END QDFZRBS

MACRO QDFZRBT
    CLASS CORE ;
    FOREIGN QDFZRBT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.140 10.470 2.540 ;
        RECT  10.090 1.930 10.370 2.650 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.270 2.310 2.670 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.050 1.260 15.330 3.780 ;
        RECT  13.470 3.500 15.330 3.780 ;
        RECT  13.470 1.260 15.330 1.540 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.380 4.650 0.560 ;
        RECT  10.110 -0.380 10.510 0.560 ;
        RECT  12.750 -0.380 13.150 0.860 ;
        RECT  14.190 -0.380 14.590 0.860 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 4.020 4.720 5.420 ;
        RECT  10.080 4.480 10.480 5.420 ;
        RECT  11.660 4.480 12.060 5.420 ;
        RECT  12.470 4.480 12.870 5.420 ;
        RECT  14.190 4.260 14.590 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  2.090 4.480 2.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 4.180 7.760 4.420 ;
        RECT  7.520 3.580 7.760 4.420 ;
        RECT  6.320 0.620 6.560 4.420 ;
        RECT  6.240 3.620 6.560 4.020 ;
        RECT  7.520 3.580 13.230 3.820 ;
        RECT  12.990 1.100 13.230 3.820 ;
        RECT  12.190 1.100 13.230 1.340 ;
        RECT  12.190 0.620 12.430 1.340 ;
        RECT  12.030 0.620 12.430 0.860 ;
        RECT  6.160 0.620 6.560 0.860 ;
        RECT  10.870 3.100 12.750 3.340 ;
        RECT  12.510 1.640 12.750 3.340 ;
        RECT  11.520 1.640 12.750 1.880 ;
        RECT  11.520 1.570 11.920 1.880 ;
        RECT  6.800 3.700 7.280 3.940 ;
        RECT  6.800 1.100 7.040 3.940 ;
        RECT  10.840 2.220 11.690 2.460 ;
        RECT  10.840 1.120 11.080 2.460 ;
        RECT  8.690 1.120 11.080 1.360 ;
        RECT  6.800 1.100 8.930 1.340 ;
        RECT  7.170 0.860 7.570 1.340 ;
        RECT  9.440 0.620 9.840 0.880 ;
        RECT  8.040 0.620 9.840 0.860 ;
        RECT  9.590 1.600 9.830 3.220 ;
        RECT  8.000 2.880 9.830 3.120 ;
        RECT  8.000 1.600 9.830 1.840 ;
        RECT  8.000 1.580 8.400 1.840 ;
        RECT  8.050 4.160 9.680 4.400 ;
        RECT  7.280 2.880 7.680 3.120 ;
        RECT  7.360 1.580 7.600 3.120 ;
        RECT  7.360 2.220 8.680 2.460 ;
        RECT  7.280 1.580 7.680 1.820 ;
        RECT  5.840 1.290 6.080 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.700 1.290 6.080 1.530 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.120 1.580 5.360 4.340 ;
        RECT  5.120 2.260 5.550 2.660 ;
        RECT  5.040 1.580 5.440 1.820 ;
        RECT  3.600 4.020 4.000 4.260 ;
        RECT  3.760 3.540 4.000 4.260 ;
        RECT  3.760 3.540 4.800 3.780 ;
        RECT  4.560 1.580 4.800 3.780 ;
        RECT  4.560 2.260 4.870 2.660 ;
        RECT  3.600 1.580 4.800 1.820 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.280 3.700 ;
        RECT  2.880 3.940 3.280 4.420 ;
        RECT  1.230 3.940 3.280 4.180 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
    END
END QDFZRBT

MACRO QDFZRSBN
    CLASS CORE ;
    FOREIGN QDFZRSBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.950 2.140 12.230 3.210 ;
        RECT  11.560 2.140 12.230 2.540 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.270 2.310 2.670 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.050 1.300 15.330 3.400 ;
        RECT  15.020 3.000 15.330 3.400 ;
        RECT  15.020 1.300 15.330 1.700 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.960 1.620 11.200 2.450 ;
        RECT  9.230 2.210 11.200 2.450 ;
        RECT  11.960 1.100 12.200 1.860 ;
        RECT  10.960 1.620 12.200 1.860 ;
        RECT  11.960 1.100 13.470 1.340 ;
        RECT  13.190 1.100 13.470 2.210 ;
        RECT  9.230 2.140 9.470 2.540 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.380 4.650 0.560 ;
        RECT  10.840 -0.380 11.240 0.560 ;
        RECT  14.220 -0.380 14.620 0.860 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 4.030 4.720 5.420 ;
        RECT  11.270 4.480 11.670 5.420 ;
        RECT  13.990 4.130 14.390 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  2.090 4.480 2.490 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 4.180 7.760 4.420 ;
        RECT  7.520 3.580 7.760 4.420 ;
        RECT  6.320 0.620 6.560 4.420 ;
        RECT  6.240 3.620 6.560 4.020 ;
        RECT  10.290 3.580 12.710 3.820 ;
        RECT  12.470 2.940 12.710 3.820 ;
        RECT  7.520 3.580 9.160 3.820 ;
        RECT  8.920 3.360 10.530 3.600 ;
        RECT  12.470 2.940 14.780 3.180 ;
        RECT  14.540 1.100 14.780 3.180 ;
        RECT  13.740 1.100 14.780 1.340 ;
        RECT  13.740 0.620 13.980 1.340 ;
        RECT  12.940 0.620 13.980 0.860 ;
        RECT  6.160 0.620 6.560 0.860 ;
        RECT  12.590 2.450 14.300 2.690 ;
        RECT  14.060 2.140 14.300 2.690 ;
        RECT  12.590 1.580 12.830 2.690 ;
        RECT  12.440 1.580 12.840 1.820 ;
        RECT  12.200 4.090 13.190 4.330 ;
        RECT  12.950 3.480 13.190 4.330 ;
        RECT  12.950 3.480 14.210 3.720 ;
        RECT  6.800 3.700 7.280 3.940 ;
        RECT  6.800 1.100 7.040 3.940 ;
        RECT  8.690 1.120 11.720 1.360 ;
        RECT  11.480 0.620 11.720 1.360 ;
        RECT  6.800 1.100 8.930 1.340 ;
        RECT  7.170 0.860 7.570 1.340 ;
        RECT  11.480 0.620 12.570 0.860 ;
        RECT  10.920 2.820 11.160 3.220 ;
        RECT  8.000 2.880 11.160 3.120 ;
        RECT  8.750 1.600 8.990 3.120 ;
        RECT  8.000 1.600 10.520 1.840 ;
        RECT  8.000 1.580 8.400 1.840 ;
        RECT  8.050 4.160 11.010 4.400 ;
        RECT  9.530 3.840 9.930 4.400 ;
        RECT  10.200 0.620 10.600 0.880 ;
        RECT  8.040 0.620 10.600 0.860 ;
        RECT  7.280 2.880 7.680 3.120 ;
        RECT  7.360 1.580 7.600 3.120 ;
        RECT  8.270 2.140 8.510 2.540 ;
        RECT  7.360 2.220 8.510 2.460 ;
        RECT  7.280 1.580 7.680 1.820 ;
        RECT  5.840 1.290 6.080 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  5.700 1.290 6.080 1.530 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.120 1.580 5.360 4.350 ;
        RECT  5.120 2.260 5.550 2.660 ;
        RECT  5.040 1.580 5.440 1.820 ;
        RECT  3.600 4.030 4.000 4.270 ;
        RECT  3.760 3.540 4.000 4.270 ;
        RECT  3.760 3.540 4.800 3.780 ;
        RECT  4.560 1.580 4.800 3.780 ;
        RECT  4.560 2.260 4.870 2.660 ;
        RECT  3.600 1.580 4.800 1.820 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.280 3.700 ;
        RECT  2.880 3.940 3.280 4.420 ;
        RECT  1.230 3.940 3.280 4.180 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
    END
END QDFZRSBN

MACRO QDFZS
    CLASS CORE ;
    FOREIGN QDFZS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.120 4.170 2.840 ;
        RECT  3.830 2.230 4.170 2.630 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.120 2.310 2.840 ;
        RECT  1.940 2.220 2.310 2.620 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.140 0.630 2.540 ;
        RECT  0.170 2.120 0.450 2.840 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.220 0.620 11.500 1.540 ;
        RECT  11.330 1.260 11.610 3.200 ;
        RECT  11.100 2.800 11.610 3.200 ;
        RECT  11.100 0.620 11.500 1.020 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.140 2.970 2.540 ;
        RECT  2.650 2.120 2.930 2.840 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.170 -0.380 4.570 0.560 ;
        RECT  9.750 -0.380 9.990 0.640 ;
        RECT  11.740 -0.380 12.140 0.940 ;
        RECT  0.000 -0.380 12.400 0.380 ;
        RECT  1.850 -0.380 2.250 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.240 4.020 4.640 5.420 ;
        RECT  7.830 4.480 8.230 5.420 ;
        RECT  9.540 4.480 9.940 5.420 ;
        RECT  11.740 4.280 12.140 5.420 ;
        RECT  0.000 4.660 12.400 5.420 ;
        RECT  2.010 4.480 2.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.590 1.370 10.830 4.420 ;
        RECT  9.750 2.480 10.830 2.720 ;
        RECT  9.220 0.890 10.680 1.130 ;
        RECT  10.280 0.730 10.680 1.130 ;
        RECT  6.660 0.620 6.900 1.020 ;
        RECT  9.220 0.620 9.460 1.130 ;
        RECT  6.660 0.620 9.460 0.860 ;
        RECT  6.580 4.000 10.240 4.240 ;
        RECT  10.000 3.080 10.240 4.240 ;
        RECT  5.860 3.520 6.100 4.160 ;
        RECT  5.860 3.520 9.640 3.760 ;
        RECT  9.270 1.660 9.510 3.760 ;
        RECT  6.180 0.620 6.420 3.760 ;
        RECT  9.210 1.660 9.510 2.060 ;
        RECT  5.670 0.620 6.420 0.860 ;
        RECT  7.650 3.040 8.970 3.280 ;
        RECT  8.730 1.100 8.970 3.280 ;
        RECT  7.650 2.130 7.890 3.280 ;
        RECT  7.490 2.130 7.890 2.370 ;
        RECT  8.420 1.100 8.970 1.340 ;
        RECT  6.660 1.500 6.900 3.200 ;
        RECT  8.150 2.260 8.490 2.660 ;
        RECT  8.150 1.590 8.390 2.660 ;
        RECT  6.660 1.590 8.390 1.830 ;
        RECT  5.700 1.100 5.940 3.200 ;
        RECT  0.960 1.340 1.200 3.190 ;
        RECT  2.800 1.340 3.200 1.810 ;
        RECT  0.730 1.340 3.210 1.580 ;
        RECT  2.970 1.100 5.940 1.340 ;
        RECT  0.730 1.010 0.970 1.580 ;
        RECT  0.160 1.010 0.970 1.250 ;
        RECT  5.040 1.580 5.280 4.340 ;
        RECT  4.900 1.580 5.300 1.820 ;
        RECT  3.520 4.020 3.920 4.260 ;
        RECT  3.680 3.540 3.920 4.260 ;
        RECT  3.680 3.540 4.650 3.780 ;
        RECT  4.410 1.580 4.650 3.780 ;
        RECT  4.410 3.220 4.790 3.620 ;
        RECT  3.520 1.580 4.650 1.820 ;
        RECT  1.210 0.800 2.730 1.040 ;
        RECT  2.490 0.620 3.200 0.860 ;
        RECT  1.210 0.620 1.610 1.040 ;
        RECT  0.160 4.120 0.990 4.360 ;
        RECT  0.750 3.460 0.990 4.360 ;
        RECT  0.750 3.460 3.200 3.700 ;
        RECT  2.800 3.940 3.200 4.420 ;
        RECT  1.230 3.940 3.200 4.180 ;
    END
END QDFZS

MACRO QDLHN
    CLASS CORE ;
    FOREIGN QDLHN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.410 0.450 2.500 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.840 2.930 2.870 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 1.130 7.270 3.190 ;
        RECT  6.960 2.790 7.270 3.190 ;
        RECT  6.960 1.490 7.270 1.890 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.270 -0.380 2.670 0.560 ;
        RECT  5.620 -0.380 6.020 0.560 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  1.480 -0.380 1.880 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.270 4.470 2.670 5.420 ;
        RECT  5.870 4.480 6.270 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.950 4.470 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.890 4.180 5.630 4.420 ;
        RECT  6.390 2.100 6.630 4.230 ;
        RECT  5.390 3.990 6.630 4.230 ;
        RECT  3.890 1.390 4.130 4.420 ;
        RECT  5.580 1.490 5.820 3.190 ;
        RECT  5.390 2.100 5.820 2.500 ;
        RECT  4.730 3.700 5.150 3.940 ;
        RECT  4.910 0.620 5.150 3.940 ;
        RECT  4.430 0.800 4.670 3.190 ;
        RECT  1.660 0.800 1.900 3.190 ;
        RECT  1.660 0.800 4.670 1.040 ;
        RECT  3.320 0.770 3.720 1.040 ;
        RECT  0.160 3.990 3.650 4.230 ;
        RECT  0.780 0.670 1.020 4.230 ;
        RECT  0.780 3.430 2.140 3.670 ;
        RECT  0.300 0.670 1.020 0.910 ;
        RECT  3.170 1.390 3.410 3.190 ;
    END
END QDLHN

MACRO QDLHP
    CLASS CORE ;
    FOREIGN QDLHP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.060 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.410 0.450 2.500 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.200 2.790 2.600 ;
        RECT  2.030 1.840 2.310 2.870 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 1.490 7.270 3.190 ;
        RECT  6.860 2.790 7.270 3.190 ;
        RECT  6.860 1.490 7.270 1.890 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.170 -0.380 2.570 0.560 ;
        RECT  5.520 -0.380 5.920 0.560 ;
        RECT  7.500 -0.380 7.900 1.030 ;
        RECT  0.000 -0.380 8.060 0.380 ;
        RECT  1.380 -0.380 1.780 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.170 4.470 2.570 5.420 ;
        RECT  5.770 4.480 6.170 5.420 ;
        RECT  7.500 4.250 7.900 5.420 ;
        RECT  0.000 4.660 8.060 5.420 ;
        RECT  0.950 4.470 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.790 4.180 5.530 4.420 ;
        RECT  6.290 2.100 6.530 4.230 ;
        RECT  5.290 3.990 6.530 4.230 ;
        RECT  3.790 1.390 4.030 4.420 ;
        RECT  5.480 1.490 5.720 3.190 ;
        RECT  5.290 2.100 5.720 2.500 ;
        RECT  4.630 3.700 5.050 3.940 ;
        RECT  4.810 0.620 5.050 3.940 ;
        RECT  4.330 0.800 4.570 3.190 ;
        RECT  1.320 0.800 1.560 3.190 ;
        RECT  1.320 0.800 4.570 1.040 ;
        RECT  3.220 0.710 3.620 1.040 ;
        RECT  0.160 3.990 3.550 4.230 ;
        RECT  0.780 0.670 1.020 4.230 ;
        RECT  0.780 3.430 1.800 3.670 ;
        RECT  0.300 0.670 1.020 0.910 ;
        RECT  3.070 1.390 3.310 3.190 ;
    END
END QDLHP

MACRO QDLHRBN
    CLASS CORE ;
    FOREIGN QDLHRBN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.760 2.930 2.700 ;
        RECT  2.500 2.050 2.930 2.450 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.410 0.480 2.430 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.180 0.450 2.750 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.860 3.550 2.870 ;
        RECT  3.210 2.180 3.550 2.580 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.430 2.790 7.890 3.190 ;
        RECT  7.610 1.280 7.890 3.300 ;
        RECT  7.430 1.280 7.890 1.680 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.310 -0.380 6.710 0.560 ;
        RECT  8.120 -0.380 8.520 0.990 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  1.260 -0.380 2.330 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 4.480 2.940 5.420 ;
        RECT  6.630 4.480 7.030 5.420 ;
        RECT  8.120 4.260 8.520 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.760 4.180 6.250 4.420 ;
        RECT  6.950 2.020 7.190 4.230 ;
        RECT  6.010 3.990 7.190 4.230 ;
        RECT  4.760 0.620 5.000 4.420 ;
        RECT  2.020 0.800 2.260 3.190 ;
        RECT  2.020 0.800 2.810 1.040 ;
        RECT  4.630 0.620 5.000 1.020 ;
        RECT  2.570 0.620 5.000 0.860 ;
        RECT  5.830 2.870 6.440 3.110 ;
        RECT  5.830 1.460 6.070 3.110 ;
        RECT  5.830 1.460 6.440 1.700 ;
        RECT  5.350 3.700 5.750 3.940 ;
        RECT  5.350 0.620 5.590 3.940 ;
        RECT  4.280 1.750 4.520 4.420 ;
        RECT  1.200 3.430 4.520 3.670 ;
        RECT  1.200 2.790 1.440 3.670 ;
        RECT  1.260 1.310 1.500 3.030 ;
        RECT  3.790 1.210 4.030 3.190 ;
        RECT  0.160 3.910 0.560 4.380 ;
        RECT  0.160 3.910 3.920 4.150 ;
        RECT  0.720 2.050 0.960 4.150 ;
        RECT  0.780 0.670 1.020 2.290 ;
        RECT  0.190 0.670 1.020 0.910 ;
    END
END QDLHRBN

MACRO QDLHRBP
    CLASS CORE ;
    FOREIGN QDLHRBP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.300 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.760 2.930 2.700 ;
        RECT  2.500 2.050 2.930 2.450 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.410 0.480 2.430 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.180 0.450 2.750 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.860 3.550 2.870 ;
        RECT  3.210 2.180 3.550 2.580 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.200 1.460 8.540 3.110 ;
        RECT  8.020 2.870 8.540 3.110 ;
        RECT  8.020 1.460 8.540 1.700 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.310 -0.380 6.710 0.560 ;
        RECT  7.300 -0.380 7.700 0.920 ;
        RECT  8.740 -0.380 9.140 0.920 ;
        RECT  0.000 -0.380 9.300 0.380 ;
        RECT  1.260 -0.380 2.330 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 4.480 2.940 5.420 ;
        RECT  6.630 4.480 7.030 5.420 ;
        RECT  8.740 4.260 9.140 5.420 ;
        RECT  0.000 4.660 9.300 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.760 4.180 6.250 4.420 ;
        RECT  6.950 2.020 7.190 4.230 ;
        RECT  6.010 3.990 7.190 4.230 ;
        RECT  4.760 0.620 5.000 4.420 ;
        RECT  2.020 0.800 2.260 3.190 ;
        RECT  2.020 0.800 2.810 1.040 ;
        RECT  4.630 0.620 5.000 1.020 ;
        RECT  2.570 0.620 5.000 0.860 ;
        RECT  5.830 2.870 6.440 3.110 ;
        RECT  5.830 1.460 6.070 3.110 ;
        RECT  5.830 1.460 6.440 1.700 ;
        RECT  5.350 3.700 5.750 3.940 ;
        RECT  5.350 0.620 5.590 3.940 ;
        RECT  4.280 1.750 4.520 4.420 ;
        RECT  1.200 3.430 4.520 3.670 ;
        RECT  1.200 2.790 1.440 3.670 ;
        RECT  1.260 1.310 1.500 3.030 ;
        RECT  3.790 1.210 4.030 3.190 ;
        RECT  3.520 3.910 3.920 4.420 ;
        RECT  0.160 3.910 0.560 4.380 ;
        RECT  0.160 3.910 3.920 4.150 ;
        RECT  0.720 2.050 0.960 4.150 ;
        RECT  0.780 0.670 1.020 2.290 ;
        RECT  0.190 0.670 1.020 0.910 ;
    END
END QDLHRBP

MACRO QDLHRBS
    CLASS CORE ;
    FOREIGN QDLHRBS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.760 2.930 2.700 ;
        RECT  2.500 2.050 2.930 2.450 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.410 0.480 2.430 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.180 0.450 2.750 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.860 3.550 2.870 ;
        RECT  3.210 2.180 3.550 2.580 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.430 2.790 7.890 3.190 ;
        RECT  7.610 1.280 7.890 3.300 ;
        RECT  7.430 1.280 7.890 1.680 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  6.310 -0.380 6.710 0.560 ;
        RECT  8.120 -0.380 8.520 0.560 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  1.260 -0.380 2.330 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 4.480 2.940 5.420 ;
        RECT  6.630 4.480 7.030 5.420 ;
        RECT  8.120 4.480 8.520 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.760 4.180 6.250 4.420 ;
        RECT  6.950 2.020 7.190 4.230 ;
        RECT  6.010 3.990 7.190 4.230 ;
        RECT  4.760 0.620 5.000 4.420 ;
        RECT  2.020 0.800 2.260 3.190 ;
        RECT  2.020 0.800 2.810 1.040 ;
        RECT  4.630 0.620 5.000 1.020 ;
        RECT  2.570 0.620 5.000 0.860 ;
        RECT  5.830 2.870 6.440 3.110 ;
        RECT  5.830 1.460 6.070 3.110 ;
        RECT  5.830 1.460 6.440 1.700 ;
        RECT  5.350 3.700 5.750 3.940 ;
        RECT  5.350 0.620 5.590 3.940 ;
        RECT  4.280 1.750 4.520 4.420 ;
        RECT  1.200 3.430 4.520 3.670 ;
        RECT  1.200 2.790 1.440 3.670 ;
        RECT  1.260 1.310 1.500 3.030 ;
        RECT  3.790 1.210 4.030 3.190 ;
        RECT  0.160 3.910 0.560 4.380 ;
        RECT  0.160 3.910 3.920 4.150 ;
        RECT  0.720 2.050 0.960 4.150 ;
        RECT  0.780 0.670 1.020 2.290 ;
        RECT  0.190 0.670 1.020 0.910 ;
    END
END QDLHRBS

MACRO QDLHS
    CLASS CORE ;
    FOREIGN QDLHS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.440 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.410 0.450 2.500 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.840 2.930 2.870 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 0.990 7.270 3.190 ;
        RECT  6.960 2.790 7.270 3.190 ;
        RECT  6.960 1.490 7.270 1.890 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 -0.380 2.700 0.560 ;
        RECT  5.740 -0.380 6.140 0.560 ;
        RECT  6.820 -0.380 7.220 0.560 ;
        RECT  0.000 -0.380 7.440 0.380 ;
        RECT  1.480 -0.380 1.880 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 4.470 2.700 5.420 ;
        RECT  6.010 4.480 6.410 5.420 ;
        RECT  0.000 4.660 7.440 5.420 ;
        RECT  0.950 4.470 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.890 4.180 5.770 4.420 ;
        RECT  6.390 2.100 6.630 4.230 ;
        RECT  5.530 3.990 6.630 4.230 ;
        RECT  3.890 1.390 4.130 4.420 ;
        RECT  5.580 1.490 5.820 3.190 ;
        RECT  5.390 2.100 5.820 2.500 ;
        RECT  4.730 3.700 5.150 3.940 ;
        RECT  4.910 0.620 5.150 3.940 ;
        RECT  4.430 0.800 4.670 3.190 ;
        RECT  1.260 0.800 1.500 3.190 ;
        RECT  1.260 0.800 4.670 1.040 ;
        RECT  0.160 3.990 3.650 4.230 ;
        RECT  0.780 0.670 1.020 4.230 ;
        RECT  0.780 3.430 1.740 3.670 ;
        RECT  0.300 0.670 1.020 0.910 ;
        RECT  3.170 1.390 3.410 3.190 ;
    END
END QDLHS

MACRO QDLHSN
    CLASS CORE ;
    FOREIGN QDLHSN 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.480 2.500 ;
        RECT  0.170 1.410 0.540 1.810 ;
        RECT  0.170 1.180 0.450 2.750 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.860 4.170 2.870 ;
        END
    END D
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.640 3.550 2.700 ;
        RECT  3.250 2.050 3.550 2.450 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.200 2.870 8.510 3.270 ;
        RECT  8.230 1.180 8.510 3.300 ;
        RECT  8.200 1.490 8.510 1.890 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.290 -0.380 3.690 0.840 ;
        RECT  7.090 -0.380 7.490 0.560 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  1.240 -0.380 1.640 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.690 4.480 3.090 5.420 ;
        RECT  7.170 4.480 7.570 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.690 4.480 1.090 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.370 4.180 6.930 4.420 ;
        RECT  7.630 2.150 7.870 4.230 ;
        RECT  6.690 3.990 7.870 4.230 ;
        RECT  5.370 0.730 5.610 4.420 ;
        RECT  2.620 3.520 5.610 3.760 ;
        RECT  2.620 1.560 2.860 3.760 ;
        RECT  2.540 1.560 2.940 1.800 ;
        RECT  6.900 1.490 7.140 3.190 ;
        RECT  6.710 2.190 7.140 2.590 ;
        RECT  6.050 3.700 6.450 3.940 ;
        RECT  6.130 0.730 6.370 3.940 ;
        RECT  0.160 3.520 1.020 3.760 ;
        RECT  0.780 0.670 1.020 3.760 ;
        RECT  0.780 2.380 1.600 2.780 ;
        RECT  4.890 0.780 5.130 2.700 ;
        RECT  1.310 0.800 1.550 2.780 ;
        RECT  2.600 1.080 4.170 1.320 ;
        RECT  3.930 0.780 4.170 1.320 ;
        RECT  2.600 0.800 2.840 1.320 ;
        RECT  1.310 0.800 2.840 1.040 ;
        RECT  3.930 0.780 5.130 1.020 ;
        RECT  0.190 0.670 1.020 0.910 ;
        RECT  1.900 4.000 5.130 4.240 ;
        RECT  1.900 1.280 2.140 4.240 ;
        RECT  1.880 3.120 2.140 3.520 ;
        RECT  1.900 1.280 2.260 1.680 ;
        RECT  4.410 1.390 4.650 3.240 ;
    END
END QDLHSN

MACRO RAM2
    CLASS CORE ;
    FOREIGN RAM2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 2.220 7.490 2.620 ;
        RECT  6.990 2.220 7.270 2.740 ;
        END
    END RD
    PIN QBZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.110 3.650 8.510 3.890 ;
        RECT  8.230 2.820 9.750 3.060 ;
        RECT  9.470 0.620 9.750 4.380 ;
        RECT  9.350 4.140 9.750 4.380 ;
        RECT  8.060 0.620 9.760 0.860 ;
        RECT  8.230 2.820 8.510 3.890 ;
        END
    END QBZ
    PIN W
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 0.860 1.070 2.740 ;
        RECT  0.790 0.860 1.380 1.100 ;
        RECT  1.140 0.620 2.170 0.860 ;
        RECT  0.710 2.150 1.070 2.550 ;
        END
    END W
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 0.620 5.410 3.310 ;
        RECT  5.020 3.070 5.420 3.310 ;
        RECT  5.020 0.620 5.410 1.020 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 1.690 2.950 ;
        RECT  1.390 2.250 1.690 2.650 ;
        END
    END D
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.840 -0.380 4.240 0.560 ;
        RECT  5.740 -0.380 5.980 0.860 ;
        RECT  7.320 -0.380 7.720 0.860 ;
        RECT  0.000 -0.380 9.920 0.380 ;
        RECT  0.500 -0.380 0.900 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.200 4.480 4.600 5.420 ;
        RECT  5.630 4.260 6.030 5.420 ;
        RECT  6.980 4.080 7.380 5.420 ;
        RECT  0.000 4.660 9.920 5.420 ;
        RECT  0.840 4.470 1.240 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.930 1.100 9.170 1.700 ;
        RECT  6.260 1.100 6.660 1.470 ;
        RECT  6.260 1.100 9.170 1.340 ;
        RECT  7.630 4.130 9.060 4.370 ;
        RECT  8.820 3.300 9.060 4.370 ;
        RECT  7.630 3.550 7.870 4.370 ;
        RECT  6.340 3.550 7.870 3.790 ;
        RECT  8.820 3.300 9.170 3.700 ;
        RECT  6.340 2.980 6.580 3.790 ;
        RECT  7.640 2.850 7.970 3.250 ;
        RECT  7.730 1.580 7.970 3.250 ;
        RECT  7.730 2.340 9.110 2.580 ;
        RECT  7.610 1.580 8.010 1.820 ;
        RECT  3.770 3.720 6.010 3.960 ;
        RECT  5.770 2.120 6.010 3.960 ;
        RECT  3.770 3.310 4.600 3.960 ;
        RECT  3.770 1.750 4.010 3.960 ;
        RECT  3.610 2.690 4.010 3.090 ;
        RECT  3.770 1.750 4.410 1.990 ;
        RECT  2.090 4.020 2.650 4.420 ;
        RECT  2.410 0.800 2.650 4.420 ;
        RECT  2.410 2.790 2.890 3.190 ;
        RECT  4.540 2.310 4.890 2.710 ;
        RECT  4.650 1.260 4.890 2.710 ;
        RECT  2.260 1.280 2.660 1.520 ;
        RECT  4.540 0.800 4.780 1.500 ;
        RECT  2.410 0.800 4.780 1.040 ;
        RECT  2.890 3.540 3.370 3.940 ;
        RECT  3.130 2.360 3.370 3.940 ;
        RECT  3.050 1.280 3.290 2.600 ;
        RECT  2.980 1.280 3.380 1.520 ;
        RECT  1.930 1.760 2.170 3.190 ;
        RECT  1.700 1.280 1.940 2.000 ;
        RECT  1.540 1.280 1.940 1.520 ;
        RECT  1.410 3.430 2.160 3.670 ;
        RECT  0.120 3.300 1.650 3.540 ;
        RECT  0.120 2.900 0.480 3.540 ;
        RECT  0.120 1.320 0.360 3.540 ;
        RECT  0.120 1.320 0.480 1.720 ;
        RECT  1.450 3.990 1.850 4.350 ;
        RECT  0.290 3.990 1.850 4.230 ;
        RECT  0.290 3.870 0.690 4.230 ;
    END
END RAM2

MACRO RAM2S
    CLASS CORE ;
    FOREIGN RAM2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN RD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.100 8.510 3.300 ;
        RECT  8.200 2.220 8.510 2.620 ;
        END
    END RD
    PIN QBZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 1.260 7.480 1.540 ;
        RECT  6.370 2.940 7.480 3.220 ;
        RECT  6.370 1.260 6.650 3.220 ;
        END
    END QBZ
    PIN W
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 0.910 1.070 2.740 ;
        RECT  0.790 0.910 2.170 1.150 ;
        RECT  0.710 2.150 1.070 2.550 ;
        END
    END W
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 2.950 5.580 3.190 ;
        RECT  5.130 1.320 5.410 3.190 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.130 1.690 2.920 ;
        END
    END D
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.230 -0.380 4.630 0.560 ;
        RECT  5.660 -0.380 6.060 0.560 ;
        RECT  7.900 -0.380 8.300 0.560 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  0.970 -0.380 1.370 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.290 4.480 4.690 5.420 ;
        RECT  5.810 4.260 6.210 5.420 ;
        RECT  7.900 4.480 8.300 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.600 4.470 1.000 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.720 3.760 8.300 4.000 ;
        RECT  7.720 1.040 7.960 4.000 ;
        RECT  6.890 2.390 7.960 2.630 ;
        RECT  7.720 1.040 8.300 1.280 ;
        RECT  3.930 3.240 4.410 3.640 ;
        RECT  3.930 1.350 4.170 3.640 ;
        RECT  5.890 0.800 6.130 2.520 ;
        RECT  3.800 1.910 4.170 2.310 ;
        RECT  3.930 1.350 4.640 1.590 ;
        RECT  4.400 0.800 4.640 1.590 ;
        RECT  4.400 0.800 6.130 1.040 ;
        RECT  2.150 4.180 4.040 4.420 ;
        RECT  4.650 1.910 4.890 4.240 ;
        RECT  3.800 4.000 4.890 4.240 ;
        RECT  2.460 1.540 2.700 4.420 ;
        RECT  2.460 2.840 2.890 3.240 ;
        RECT  2.410 1.540 2.700 1.940 ;
        RECT  2.940 3.700 3.370 3.940 ;
        RECT  3.130 0.620 3.370 3.940 ;
        RECT  3.030 0.620 3.430 0.860 ;
        RECT  1.930 1.620 2.170 3.240 ;
        RECT  1.540 1.620 2.170 1.860 ;
        RECT  1.010 3.480 2.160 3.720 ;
        RECT  0.120 3.390 1.250 3.630 ;
        RECT  0.120 3.080 0.480 3.630 ;
        RECT  0.120 1.490 0.360 3.630 ;
        RECT  0.120 1.490 0.480 1.890 ;
        RECT  1.510 3.980 1.910 4.420 ;
        RECT  0.260 3.980 1.910 4.220 ;
        RECT  0.260 3.870 0.660 4.220 ;
    END
END RAM2S

MACRO RAM3
    CLASS CORE ;
    FOREIGN RAM3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.540 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN QZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 2.820 9.130 3.300 ;
        RECT  8.810 2.820 10.370 3.060 ;
        RECT  10.090 0.620 10.370 4.380 ;
        RECT  9.970 4.140 10.370 4.380 ;
        RECT  8.680 0.620 10.380 0.860 ;
        RECT  8.810 2.820 9.130 3.250 ;
        END
    END QZ
    PIN RD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.610 2.280 8.060 2.680 ;
        RECT  7.610 2.220 7.890 2.740 ;
        END
    END RD
    PIN W
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 0.910 1.070 2.740 ;
        RECT  0.790 0.910 2.220 1.150 ;
        RECT  0.710 2.150 1.070 2.550 ;
        END
    END W
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.060 1.690 2.740 ;
        RECT  1.390 2.300 1.690 2.700 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.500 6.030 3.270 ;
        RECT  5.450 2.870 6.030 3.270 ;
        RECT  5.600 1.500 6.030 1.740 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.220 -0.380 4.620 0.560 ;
        RECT  6.240 -0.380 6.640 0.780 ;
        RECT  7.500 -0.380 7.900 0.860 ;
        RECT  0.000 -0.380 10.540 0.380 ;
        RECT  0.970 -0.380 1.370 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.060 4.480 4.460 5.420 ;
        RECT  5.980 4.080 6.380 5.420 ;
        RECT  7.390 4.080 7.790 5.420 ;
        RECT  0.000 4.660 10.540 5.420 ;
        RECT  0.980 4.470 1.380 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.550 1.100 9.790 1.700 ;
        RECT  6.860 1.100 7.260 1.440 ;
        RECT  6.860 1.100 9.790 1.340 ;
        RECT  6.690 3.590 9.790 3.830 ;
        RECT  9.550 3.300 9.790 3.830 ;
        RECT  6.690 2.980 6.930 3.830 ;
        RECT  8.050 2.940 8.550 3.340 ;
        RECT  8.310 1.580 8.550 3.340 ;
        RECT  8.310 2.340 9.730 2.580 ;
        RECT  8.230 1.580 8.630 1.820 ;
        RECT  3.240 0.850 3.480 3.660 ;
        RECT  6.380 1.020 6.620 2.620 ;
        RECT  3.240 1.570 3.830 1.810 ;
        RECT  5.590 1.020 6.620 1.260 ;
        RECT  3.240 0.950 5.830 1.190 ;
        RECT  3.240 0.850 3.660 1.190 ;
        RECT  4.730 1.490 4.970 3.650 ;
        RECT  3.730 2.110 4.970 2.350 ;
        RECT  4.730 1.490 5.200 1.890 ;
        RECT  2.480 4.110 2.960 4.350 ;
        RECT  2.720 1.490 2.960 4.350 ;
        RECT  4.220 2.710 4.460 4.140 ;
        RECT  2.720 3.900 4.460 4.140 ;
        RECT  2.480 2.840 2.960 3.240 ;
        RECT  2.550 1.490 2.960 1.890 ;
        RECT  1.020 3.500 2.480 3.740 ;
        RECT  0.190 3.290 1.260 3.530 ;
        RECT  0.190 2.900 0.480 3.530 ;
        RECT  0.190 1.490 0.430 3.530 ;
        RECT  0.190 1.490 0.480 1.890 ;
        RECT  1.540 2.980 2.170 3.220 ;
        RECT  1.930 1.570 2.170 3.220 ;
        RECT  1.610 1.570 2.170 1.810 ;
        RECT  1.620 3.990 2.020 4.420 ;
        RECT  0.470 3.990 2.020 4.230 ;
        RECT  0.470 3.780 0.710 4.230 ;
    END
END RAM3

MACRO RAM3S
    CLASS CORE ;
    FOREIGN RAM3S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.300 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN QZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.990 1.260 8.010 1.540 ;
        RECT  6.990 2.940 8.040 3.220 ;
        RECT  6.990 1.260 7.270 3.220 ;
        END
    END QZ
    PIN RD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.850 2.100 9.130 3.300 ;
        RECT  8.820 2.220 9.130 2.620 ;
        END
    END RD
    PIN W
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 0.910 1.070 2.740 ;
        RECT  0.790 0.910 2.220 1.150 ;
        RECT  0.710 2.150 1.070 2.550 ;
        END
    END W
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.080 1.690 2.740 ;
        RECT  1.390 2.300 1.690 2.700 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.630 2.870 6.030 3.270 ;
        RECT  5.750 1.280 6.030 3.300 ;
        RECT  5.640 1.320 6.030 1.720 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.240 -0.380 5.210 0.560 ;
        RECT  6.100 -0.380 6.500 0.560 ;
        RECT  8.520 -0.380 8.920 0.560 ;
        RECT  0.000 -0.380 9.300 0.380 ;
        RECT  0.970 -0.380 1.370 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.040 4.480 4.440 5.420 ;
        RECT  6.330 4.080 6.770 5.420 ;
        RECT  8.520 4.480 8.920 5.420 ;
        RECT  0.000 4.660 9.300 5.420 ;
        RECT  0.980 4.470 1.380 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.310 3.760 8.920 4.000 ;
        RECT  8.310 1.040 8.550 4.000 ;
        RECT  7.510 2.390 8.550 2.630 ;
        RECT  8.310 1.040 8.920 1.280 ;
        RECT  3.330 0.800 3.570 3.660 ;
        RECT  6.350 0.800 6.590 2.520 ;
        RECT  3.330 1.570 3.850 1.810 ;
        RECT  3.260 0.850 3.660 1.090 ;
        RECT  3.330 0.800 6.590 1.040 ;
        RECT  4.910 1.490 5.150 3.650 ;
        RECT  3.920 2.110 5.150 2.350 ;
        RECT  2.480 4.110 2.960 4.350 ;
        RECT  2.720 1.490 2.960 4.350 ;
        RECT  4.420 2.710 4.660 4.140 ;
        RECT  2.720 3.900 4.660 4.140 ;
        RECT  2.480 2.840 2.960 3.240 ;
        RECT  2.550 1.490 2.960 1.890 ;
        RECT  1.040 3.500 2.480 3.740 ;
        RECT  0.220 3.300 1.280 3.540 ;
        RECT  0.220 2.900 0.480 3.540 ;
        RECT  0.220 1.490 0.460 3.540 ;
        RECT  0.220 1.490 0.480 1.890 ;
        RECT  1.540 2.980 2.170 3.220 ;
        RECT  1.930 1.570 2.170 3.220 ;
        RECT  1.610 1.570 2.170 1.810 ;
        RECT  1.620 3.990 2.020 4.420 ;
        RECT  0.390 3.990 2.020 4.230 ;
        RECT  0.390 3.870 0.790 4.230 ;
    END
END RAM3S

MACRO RAM5
    CLASS CORE ;
    FOREIGN RAM5 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN QZ1
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.550 2.870 14.090 3.110 ;
        RECT  13.810 0.620 14.090 4.420 ;
        RECT  13.690 4.180 14.090 4.420 ;
        RECT  12.420 0.620 14.100 0.860 ;
        RECT  12.550 2.870 12.790 3.270 ;
        END
    END QZ1
    PIN QZ0
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.490 2.940 6.030 3.180 ;
        RECT  5.750 2.820 7.270 3.060 ;
        RECT  7.030 2.820 7.270 3.250 ;
        RECT  5.570 0.620 7.430 0.860 ;
        RECT  5.750 0.620 6.030 3.180 ;
        END
    END QZ0
    PIN W
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.150 0.480 2.550 ;
        RECT  0.170 2.150 0.450 2.740 ;
        END
    END W
    PIN RD1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 2.280 11.790 2.680 ;
        RECT  11.330 2.220 11.610 2.740 ;
        END
    END RD1
    PIN RD0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.220 8.510 2.740 ;
        RECT  8.020 2.280 8.510 2.680 ;
        END
    END RD0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.050 1.690 2.740 ;
        RECT  1.250 2.300 1.690 2.700 ;
        END
    END D
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.220 -0.380 4.620 0.560 ;
        RECT  8.180 -0.380 8.580 0.860 ;
        RECT  9.680 -0.380 10.080 0.860 ;
        RECT  11.030 -0.380 11.430 0.860 ;
        RECT  0.000 -0.380 14.260 0.380 ;
        RECT  0.970 -0.380 1.370 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.060 4.480 4.460 5.420 ;
        RECT  8.090 4.480 8.490 5.420 ;
        RECT  9.690 4.080 10.090 5.420 ;
        RECT  11.110 4.080 11.510 5.420 ;
        RECT  0.000 4.660 14.260 5.420 ;
        RECT  0.980 4.470 1.380 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.440 3.590 13.510 3.830 ;
        RECT  13.270 3.350 13.510 3.830 ;
        RECT  10.440 2.980 10.680 3.830 ;
        RECT  11.790 2.940 12.270 3.340 ;
        RECT  12.030 1.580 12.270 3.340 ;
        RECT  12.030 2.390 13.450 2.630 ;
        RECT  11.690 1.580 12.270 1.820 ;
        RECT  13.140 1.100 13.380 1.700 ;
        RECT  10.390 1.100 10.790 1.440 ;
        RECT  10.390 1.100 13.380 1.340 ;
        RECT  4.820 3.980 9.070 4.220 ;
        RECT  8.830 3.540 9.070 4.220 ;
        RECT  3.240 3.940 5.060 4.180 ;
        RECT  3.240 1.600 3.480 4.180 ;
        RECT  8.830 3.540 9.950 3.780 ;
        RECT  9.710 2.220 9.950 3.780 ;
        RECT  9.700 2.220 9.950 2.620 ;
        RECT  3.240 1.600 3.830 1.840 ;
        RECT  6.310 3.500 8.590 3.740 ;
        RECT  8.350 3.060 8.590 3.740 ;
        RECT  6.310 3.300 6.550 3.740 ;
        RECT  8.350 3.060 9.420 3.300 ;
        RECT  6.290 1.100 6.530 1.700 ;
        RECT  8.820 1.100 9.220 1.440 ;
        RECT  6.290 1.100 9.220 1.340 ;
        RECT  7.530 3.020 8.070 3.260 ;
        RECT  7.530 1.580 7.770 3.260 ;
        RECT  6.350 2.340 7.770 2.580 ;
        RECT  7.450 1.580 7.850 1.820 ;
        RECT  4.720 2.790 5.140 3.650 ;
        RECT  4.900 1.520 5.140 3.650 ;
        RECT  3.730 2.790 5.140 3.030 ;
        RECT  4.900 1.520 5.200 1.920 ;
        RECT  2.480 4.110 2.960 4.350 ;
        RECT  2.720 0.800 2.960 4.350 ;
        RECT  2.480 2.840 2.960 3.240 ;
        RECT  4.220 2.060 4.660 2.460 ;
        RECT  4.220 0.800 4.460 2.460 ;
        RECT  2.550 1.490 2.960 1.890 ;
        RECT  2.720 0.800 4.460 1.040 ;
        RECT  1.030 3.500 2.480 3.740 ;
        RECT  1.030 2.980 1.270 3.740 ;
        RECT  0.160 2.980 1.270 3.220 ;
        RECT  0.770 1.570 1.010 3.220 ;
        RECT  0.160 1.570 1.010 1.810 ;
        RECT  0.390 0.910 0.790 1.270 ;
        RECT  0.390 0.910 2.220 1.150 ;
        RECT  1.540 2.980 2.170 3.220 ;
        RECT  1.930 1.570 2.170 3.220 ;
        RECT  1.610 1.570 2.170 1.810 ;
        RECT  1.620 3.990 2.020 4.420 ;
        RECT  0.470 3.990 2.020 4.230 ;
        RECT  0.470 3.460 0.710 4.230 ;
    END
END RAM5

MACRO RAM5S
    CLASS CORE ;
    FOREIGN RAM5S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN QZ1
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.830 4.140 12.230 4.380 ;
        RECT  11.840 1.430 12.240 1.670 ;
        RECT  11.950 1.430 12.230 4.380 ;
        END
    END QZ1
    PIN QZ0
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.430 6.030 3.250 ;
        RECT  5.620 2.850 6.030 3.250 ;
        RECT  5.600 1.430 6.030 1.670 ;
        END
    END QZ0
    PIN W
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.150 0.480 2.550 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END W
    PIN RD1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.090 2.280 10.550 2.680 ;
        RECT  10.090 2.220 10.370 2.740 ;
        END
    END RD1
    PIN RD0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.610 2.220 7.890 2.740 ;
        RECT  7.370 2.280 7.890 2.680 ;
        END
    END RD0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.050 1.690 2.740 ;
        RECT  1.250 2.300 1.690 2.700 ;
        END
    END D
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.220 -0.380 4.620 0.560 ;
        RECT  7.680 -0.380 8.080 0.860 ;
        RECT  9.740 -0.380 10.140 0.860 ;
        RECT  0.000 -0.380 12.400 0.380 ;
        RECT  0.970 -0.380 1.370 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.060 4.480 4.460 5.420 ;
        RECT  7.470 4.460 7.870 5.420 ;
        RECT  10.030 4.080 10.430 5.420 ;
        RECT  0.000 4.660 12.400 5.420 ;
        RECT  0.980 4.470 1.380 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.330 3.590 11.650 3.830 ;
        RECT  11.410 3.300 11.650 3.830 ;
        RECT  9.330 2.980 9.570 3.830 ;
        RECT  10.690 2.940 11.040 3.340 ;
        RECT  10.800 1.580 11.040 3.340 ;
        RECT  10.800 2.390 11.590 2.630 ;
        RECT  10.470 1.580 11.040 1.820 ;
        RECT  9.100 1.100 9.500 1.440 ;
        RECT  9.100 1.100 11.360 1.340 ;
        RECT  11.120 0.670 11.360 1.340 ;
        RECT  11.120 0.670 11.520 0.910 ;
        RECT  5.030 4.060 6.990 4.300 ;
        RECT  3.240 3.920 5.270 4.160 ;
        RECT  6.750 3.980 9.090 4.220 ;
        RECT  8.850 2.360 9.090 4.220 ;
        RECT  3.240 1.570 3.480 4.160 ;
        RECT  8.870 2.220 9.110 2.620 ;
        RECT  3.240 1.570 3.830 1.810 ;
        RECT  8.340 1.100 8.740 1.440 ;
        RECT  6.270 1.100 8.740 1.340 ;
        RECT  6.270 0.620 6.510 1.340 ;
        RECT  6.270 0.620 6.720 0.860 ;
        RECT  6.110 3.500 6.510 3.820 ;
        RECT  6.110 3.500 8.610 3.740 ;
        RECT  8.370 2.980 8.610 3.740 ;
        RECT  6.800 3.020 7.230 3.260 ;
        RECT  6.800 1.580 7.040 3.260 ;
        RECT  6.270 2.390 7.040 2.630 ;
        RECT  6.800 1.580 7.370 1.820 ;
        RECT  4.900 1.490 5.140 3.650 ;
        RECT  3.730 2.790 5.140 3.030 ;
        RECT  4.900 1.490 5.200 1.890 ;
        RECT  2.480 4.110 2.960 4.350 ;
        RECT  2.720 0.860 2.960 4.350 ;
        RECT  2.480 2.840 2.960 3.240 ;
        RECT  4.420 0.860 4.660 2.430 ;
        RECT  2.550 1.490 2.960 1.890 ;
        RECT  2.720 0.860 4.660 1.100 ;
        RECT  0.950 3.500 2.480 3.740 ;
        RECT  0.950 2.980 1.190 3.740 ;
        RECT  0.160 2.980 1.190 3.220 ;
        RECT  0.770 1.570 1.010 3.220 ;
        RECT  0.160 1.570 1.010 1.810 ;
        RECT  0.390 0.910 0.790 1.200 ;
        RECT  0.390 0.910 2.220 1.150 ;
        RECT  1.540 2.980 2.170 3.220 ;
        RECT  1.930 1.570 2.170 3.220 ;
        RECT  1.610 1.570 2.170 1.810 ;
        RECT  1.620 3.990 2.020 4.420 ;
        RECT  0.470 3.990 2.020 4.230 ;
        RECT  0.470 3.460 0.710 4.230 ;
    END
END RAM5S

MACRO TIE0
    CLASS CORE ;
    FOREIGN TIE0 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.860 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.490 0.480 1.890 ;
        RECT  0.170 1.180 0.450 2.260 ;
        END
    END O
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.860 0.380 ;
        RECT  0.930 -0.380 1.170 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 1.860 5.420 ;
        RECT  0.680 3.910 1.080 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 2.870 0.930 3.110 ;
        RECT  0.690 2.220 0.930 3.110 ;
    END
END TIE0

MACRO TIE1
    CLASS CORE ;
    FOREIGN TIE1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.860 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.840 0.480 3.240 ;
        RECT  0.170 2.220 0.450 3.300 ;
        END
    END O
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.860 0.380 ;
        RECT  0.930 -0.380 1.170 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 1.860 5.420 ;
        RECT  0.680 3.910 1.080 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.690 1.570 0.930 2.620 ;
        RECT  0.160 1.570 0.930 1.810 ;
    END
END TIE1

MACRO XNR2H
    CLASS CORE ;
    FOREIGN XNR2H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.390 1.570 6.630 3.110 ;
        RECT  3.290 2.870 6.630 3.110 ;
        RECT  3.190 1.570 6.630 1.810 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 2.110 2.650 ;
        RECT  1.410 2.250 1.690 2.890 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.230 2.250 8.510 2.890 ;
        RECT  7.990 2.250 8.510 2.650 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 -0.380 2.070 0.560 ;
        RECT  6.600 -0.380 7.000 0.780 ;
        RECT  8.120 -0.380 8.520 0.780 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 4.480 2.170 5.420 ;
        RECT  6.680 4.260 7.080 5.420 ;
        RECT  8.120 4.260 8.520 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.990 4.000 6.430 4.240 ;
        RECT  6.190 3.640 6.430 4.240 ;
        RECT  0.450 3.780 1.230 4.020 ;
        RECT  6.190 3.640 7.720 3.880 ;
        RECT  7.480 1.090 7.720 3.880 ;
        RECT  0.450 2.250 0.690 4.020 ;
        RECT  5.350 1.090 7.720 1.330 ;
        RECT  2.070 3.350 5.850 3.590 ;
        RECT  0.930 3.300 2.310 3.540 ;
        RECT  0.930 3.140 1.200 3.540 ;
        RECT  0.930 1.090 1.170 3.540 ;
        RECT  0.930 1.090 1.200 1.490 ;
        RECT  0.930 1.090 4.310 1.330 ;
        RECT  2.460 2.870 2.960 3.110 ;
        RECT  2.460 1.570 2.700 3.110 ;
        RECT  2.460 2.330 5.680 2.570 ;
        RECT  2.460 1.570 2.860 1.810 ;
    END
END XNR2H

MACRO XNR2HP
    CLASS CORE ;
    FOREIGN XNR2HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.490 2.870 11.670 3.110 ;
        RECT  5.620 1.570 11.800 1.810 ;
        RECT  11.330 1.570 11.610 3.110 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.230 3.550 2.870 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 2.250 14.090 2.890 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.110 -0.380 3.510 0.560 ;
        RECT  4.830 -0.380 5.230 0.560 ;
        RECT  12.050 -0.380 12.450 0.780 ;
        RECT  13.500 -0.380 13.900 0.780 ;
        RECT  14.940 -0.380 15.340 0.780 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.210 4.370 3.610 5.420 ;
        RECT  4.930 4.370 5.330 5.420 ;
        RECT  12.060 4.260 12.460 5.420 ;
        RECT  13.500 4.260 13.900 5.420 ;
        RECT  14.940 4.260 15.340 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.030 3.830 11.440 4.070 ;
        RECT  11.200 3.780 14.620 4.020 ;
        RECT  0.400 3.780 3.270 4.020 ;
        RECT  12.860 1.090 13.100 4.020 ;
        RECT  0.400 2.250 0.640 4.020 ;
        RECT  9.220 1.090 14.620 1.330 ;
        RECT  3.580 3.350 10.950 3.590 ;
        RECT  0.880 3.300 3.820 3.540 ;
        RECT  2.400 1.190 2.640 3.540 ;
        RECT  0.880 1.190 3.620 1.430 ;
        RECT  3.380 1.090 8.180 1.330 ;
        RECT  4.070 2.870 5.250 3.110 ;
        RECT  5.010 1.570 5.250 3.110 ;
        RECT  5.010 2.330 9.760 2.570 ;
        RECT  3.900 1.570 5.250 1.810 ;
    END
END XNR2HP

MACRO XNR2HS
    CLASS CORE ;
    FOREIGN XNR2HS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.950 1.850 4.150 2.090 ;
        RECT  3.910 1.850 4.150 3.110 ;
        RECT  2.780 2.870 4.150 3.110 ;
        RECT  2.950 1.570 3.350 2.090 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.850 1.690 2.820 ;
        RECT  1.330 2.190 1.690 2.590 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.070 2.890 ;
        RECT  0.650 2.250 1.070 2.650 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.230 -0.380 4.630 0.560 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  1.020 -0.380 1.420 0.810 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.130 4.480 4.530 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.500 3.830 5.340 4.070 ;
        RECT  5.100 0.800 5.340 4.070 ;
        RECT  3.750 0.800 5.340 1.040 ;
        RECT  2.230 0.680 3.990 0.920 ;
        RECT  2.060 3.780 2.460 4.080 ;
        RECT  0.170 3.780 2.770 4.020 ;
        RECT  2.530 3.350 2.770 4.020 ;
        RECT  0.170 3.620 0.480 4.020 ;
        RECT  0.170 1.050 0.410 4.020 ;
        RECT  2.530 3.350 4.780 3.590 ;
        RECT  4.540 1.340 4.780 3.590 ;
        RECT  3.670 1.340 4.780 1.580 ;
        RECT  0.170 1.050 0.480 1.450 ;
        RECT  1.560 3.060 2.170 3.460 ;
        RECT  1.930 1.370 2.170 3.460 ;
        RECT  1.930 2.330 3.540 2.570 ;
        RECT  1.530 1.370 2.170 1.610 ;
    END
END XNR2HS

MACRO XNR2HT
    CLASS CORE ;
    FOREIGN XNR2HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.320 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.790 1.570 16.830 1.810 ;
        RECT  7.880 2.870 16.920 3.110 ;
        RECT  16.290 1.570 16.570 3.110 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.230 5.410 2.630 ;
        RECT  4.510 2.230 4.790 3.060 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  20.010 1.860 20.290 2.690 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.550 -0.380 4.950 0.560 ;
        RECT  6.270 -0.380 6.670 0.560 ;
        RECT  17.420 -0.380 17.820 0.870 ;
        RECT  18.880 -0.380 19.280 0.780 ;
        RECT  20.320 -0.380 20.720 0.780 ;
        RECT  21.760 -0.380 22.160 0.780 ;
        RECT  0.000 -0.380 22.320 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.650 4.310 5.050 5.420 ;
        RECT  6.370 4.310 6.770 5.420 ;
        RECT  17.360 4.120 17.760 5.420 ;
        RECT  18.880 4.260 19.280 5.420 ;
        RECT  20.320 4.260 20.720 5.420 ;
        RECT  21.760 4.260 22.160 5.420 ;
        RECT  0.000 4.660 22.320 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.640 3.830 16.680 4.070 ;
        RECT  16.440 3.540 16.680 4.070 ;
        RECT  0.400 3.780 4.880 4.020 ;
        RECT  16.440 3.540 21.440 3.780 ;
        RECT  0.400 2.250 0.640 4.020 ;
        RECT  18.240 1.110 18.480 3.780 ;
        RECT  17.070 1.110 21.440 1.350 ;
        RECT  12.830 1.090 17.310 1.330 ;
        RECT  5.030 3.350 16.200 3.590 ;
        RECT  0.880 3.300 5.270 3.540 ;
        RECT  3.840 1.190 4.080 3.540 ;
        RECT  0.880 1.190 5.060 1.430 ;
        RECT  4.820 1.090 11.790 1.330 ;
        RECT  5.510 2.870 7.560 3.110 ;
        RECT  7.150 1.570 7.390 3.110 ;
        RECT  7.150 2.330 14.820 2.570 ;
        RECT  5.340 1.570 7.460 1.810 ;
    END
END XNR2HT

MACRO XNR3
    CLASS CORE ;
    FOREIGN XNR3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.710 1.180 10.990 3.300 ;
        RECT  10.680 2.900 10.990 3.300 ;
        RECT  10.680 1.180 10.990 1.580 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.280 0.580 2.680 ;
        RECT  0.170 2.170 0.450 2.870 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.690 2.990 ;
        RECT  1.300 2.120 1.690 2.520 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 2.300 9.750 3.020 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 1.060 ;
        RECT  9.300 -0.380 10.200 0.560 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.450 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.850 4.480 2.250 5.420 ;
        RECT  9.700 4.480 10.100 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.560 0.830 7.800 3.300 ;
        RECT  10.200 2.030 10.460 2.430 ;
        RECT  10.200 0.830 10.440 2.430 ;
        RECT  7.560 0.830 10.440 1.070 ;
        RECT  8.990 3.320 9.510 3.720 ;
        RECT  8.990 1.330 9.230 3.720 ;
        RECT  8.990 1.330 9.550 1.570 ;
        RECT  4.750 4.180 8.520 4.420 ;
        RECT  8.280 1.330 8.520 4.420 ;
        RECT  4.750 1.100 4.990 4.420 ;
        RECT  3.340 2.910 3.770 3.150 ;
        RECT  3.530 1.100 3.770 3.150 ;
        RECT  3.350 1.580 3.770 1.820 ;
        RECT  8.200 1.330 8.600 1.570 ;
        RECT  3.530 1.100 4.990 1.340 ;
        RECT  5.230 3.470 7.080 3.710 ;
        RECT  6.840 1.250 7.080 3.710 ;
        RECT  5.230 1.500 5.470 3.710 ;
        RECT  6.020 0.620 6.260 3.230 ;
        RECT  2.560 2.820 3.050 3.220 ;
        RECT  2.810 0.620 3.050 3.220 ;
        RECT  5.940 1.580 6.340 1.820 ;
        RECT  2.560 1.480 3.050 1.720 ;
        RECT  2.810 0.620 6.260 0.860 ;
        RECT  1.930 3.460 4.510 3.700 ;
        RECT  4.270 1.580 4.510 3.700 ;
        RECT  1.320 3.250 1.560 3.650 ;
        RECT  1.320 3.250 2.170 3.490 ;
        RECT  1.930 1.480 2.170 3.700 ;
        RECT  4.110 2.910 4.510 3.150 ;
        RECT  1.930 2.150 2.570 2.550 ;
        RECT  4.110 1.580 4.510 1.820 ;
        RECT  1.320 1.480 2.170 1.720 ;
        RECT  0.820 4.000 3.440 4.240 ;
        RECT  0.450 3.760 1.060 4.000 ;
        RECT  0.820 1.280 1.060 4.240 ;
        RECT  0.600 1.280 1.060 1.520 ;
    END
END XNR3

MACRO XNR3P
    CLASS CORE ;
    FOREIGN XNR3P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.710 1.180 10.990 3.300 ;
        RECT  10.580 2.900 10.990 3.300 ;
        RECT  10.580 1.180 10.990 1.580 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.280 0.580 2.680 ;
        RECT  0.170 2.170 0.450 2.870 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.690 2.990 ;
        RECT  1.300 2.120 1.690 2.520 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.400 2.620 9.750 3.020 ;
        RECT  9.470 2.300 9.750 3.020 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 1.060 ;
        RECT  9.200 -0.380 10.100 0.560 ;
        RECT  11.220 -0.380 11.620 0.950 ;
        RECT  0.000 -0.380 11.780 0.380 ;
        RECT  0.450 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.850 4.480 2.250 5.420 ;
        RECT  9.600 4.480 10.000 5.420 ;
        RECT  11.220 4.260 11.620 5.420 ;
        RECT  0.000 4.660 11.780 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.560 0.830 7.800 3.300 ;
        RECT  10.100 2.030 10.360 2.430 ;
        RECT  10.100 0.830 10.340 2.430 ;
        RECT  7.560 0.830 10.340 1.070 ;
        RECT  8.890 3.320 9.410 3.720 ;
        RECT  8.890 1.330 9.130 3.720 ;
        RECT  8.890 1.330 9.450 1.570 ;
        RECT  4.750 4.180 8.520 4.420 ;
        RECT  8.280 1.330 8.520 4.420 ;
        RECT  4.750 1.100 4.990 4.420 ;
        RECT  3.340 2.910 3.770 3.150 ;
        RECT  3.530 1.100 3.770 3.150 ;
        RECT  3.350 1.580 3.770 1.820 ;
        RECT  8.200 1.330 8.600 1.570 ;
        RECT  3.530 1.100 4.990 1.340 ;
        RECT  5.230 3.470 7.080 3.710 ;
        RECT  6.840 1.250 7.080 3.710 ;
        RECT  5.230 1.500 5.470 3.710 ;
        RECT  6.020 0.620 6.260 3.230 ;
        RECT  2.560 2.820 3.050 3.220 ;
        RECT  2.810 0.620 3.050 3.220 ;
        RECT  5.940 1.580 6.340 1.820 ;
        RECT  2.560 1.480 3.050 1.720 ;
        RECT  2.810 0.620 6.260 0.860 ;
        RECT  1.930 3.460 4.510 3.700 ;
        RECT  4.270 1.580 4.510 3.700 ;
        RECT  1.320 3.250 1.560 3.650 ;
        RECT  1.320 3.250 2.170 3.490 ;
        RECT  1.930 1.480 2.170 3.700 ;
        RECT  4.110 2.910 4.510 3.150 ;
        RECT  1.930 2.150 2.570 2.550 ;
        RECT  4.110 1.580 4.510 1.820 ;
        RECT  1.320 1.480 2.170 1.720 ;
        RECT  0.820 4.000 3.440 4.240 ;
        RECT  0.450 3.760 1.060 4.000 ;
        RECT  0.820 1.280 1.060 4.240 ;
        RECT  0.600 1.280 1.060 1.520 ;
    END
END XNR3P

MACRO XNR3S
    CLASS CORE ;
    FOREIGN XNR3S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.710 0.640 10.990 3.820 ;
        RECT  10.680 3.420 10.990 3.820 ;
        RECT  10.680 0.640 10.990 1.040 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.840 0.580 3.240 ;
        RECT  0.170 2.730 0.450 3.430 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.690 2.990 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 2.300 9.750 3.020 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.120 -0.380 2.520 0.840 ;
        RECT  9.300 -0.380 10.200 0.560 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.450 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.000 4.480 2.400 5.420 ;
        RECT  9.810 4.480 10.210 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.710 0.830 7.950 3.300 ;
        RECT  10.200 2.030 10.460 2.430 ;
        RECT  10.200 0.830 10.440 2.430 ;
        RECT  7.710 0.830 10.440 1.070 ;
        RECT  8.990 3.320 9.510 3.720 ;
        RECT  8.990 1.330 9.230 3.720 ;
        RECT  8.990 1.330 9.490 1.570 ;
        RECT  4.900 4.180 8.670 4.420 ;
        RECT  8.430 1.330 8.670 4.420 ;
        RECT  4.900 1.100 5.140 4.420 ;
        RECT  3.490 2.910 3.920 3.150 ;
        RECT  3.680 1.100 3.920 3.150 ;
        RECT  3.500 1.580 3.920 1.820 ;
        RECT  8.350 1.330 8.750 1.570 ;
        RECT  3.680 1.100 5.140 1.340 ;
        RECT  5.380 3.470 7.230 3.710 ;
        RECT  6.990 1.250 7.230 3.710 ;
        RECT  5.380 1.500 5.620 3.710 ;
        RECT  6.170 0.620 6.410 3.230 ;
        RECT  2.700 2.910 3.200 3.150 ;
        RECT  2.960 0.620 3.200 3.150 ;
        RECT  6.090 1.580 6.490 1.820 ;
        RECT  2.710 1.360 3.200 1.600 ;
        RECT  2.960 0.620 6.410 0.860 ;
        RECT  1.300 3.520 4.660 3.760 ;
        RECT  4.420 1.580 4.660 3.760 ;
        RECT  2.080 1.270 2.320 3.760 ;
        RECT  4.260 2.910 4.660 3.150 ;
        RECT  2.080 2.150 2.720 2.550 ;
        RECT  4.260 1.580 4.660 1.820 ;
        RECT  1.330 1.270 2.320 1.510 ;
        RECT  2.750 4.070 3.590 4.310 ;
        RECT  0.820 4.000 2.990 4.240 ;
        RECT  0.450 3.760 1.060 4.000 ;
        RECT  0.820 1.040 1.060 4.240 ;
        RECT  0.450 1.040 1.060 1.280 ;
    END
END XNR3S

MACRO XNR3T
    CLASS CORE ;
    FOREIGN XNR3T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 1.260 11.610 3.220 ;
        RECT  10.480 1.260 12.240 1.540 ;
        RECT  10.400 2.940 12.240 3.220 ;
        RECT  10.480 1.260 10.720 1.660 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.280 0.580 2.680 ;
        RECT  0.170 2.170 0.450 2.870 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.690 2.990 ;
        RECT  1.300 2.120 1.690 2.520 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.320 2.620 9.750 3.020 ;
        RECT  9.470 2.300 9.750 3.020 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 1.060 ;
        RECT  9.100 -0.380 10.000 0.560 ;
        RECT  11.120 -0.380 11.520 0.950 ;
        RECT  0.000 -0.380 12.400 0.380 ;
        RECT  0.450 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.850 4.480 2.250 5.420 ;
        RECT  9.500 4.480 9.900 5.420 ;
        RECT  11.120 4.260 11.520 5.420 ;
        RECT  0.000 4.660 12.400 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.560 0.830 7.800 3.300 ;
        RECT  9.990 2.030 10.260 2.430 ;
        RECT  9.990 0.830 10.230 2.430 ;
        RECT  7.560 0.830 10.230 1.070 ;
        RECT  8.840 3.320 9.270 3.720 ;
        RECT  8.840 1.330 9.080 3.720 ;
        RECT  8.790 1.940 9.080 2.340 ;
        RECT  8.840 1.330 9.350 1.570 ;
        RECT  4.750 4.180 8.520 4.420 ;
        RECT  8.280 1.330 8.520 4.420 ;
        RECT  4.750 1.100 4.990 4.420 ;
        RECT  3.340 2.910 3.770 3.150 ;
        RECT  3.530 1.100 3.770 3.150 ;
        RECT  3.350 1.580 3.770 1.820 ;
        RECT  8.200 1.330 8.600 1.570 ;
        RECT  3.530 1.100 4.990 1.340 ;
        RECT  5.230 3.470 7.080 3.710 ;
        RECT  6.840 1.250 7.080 3.710 ;
        RECT  5.230 1.500 5.470 3.710 ;
        RECT  6.020 0.620 6.260 3.230 ;
        RECT  2.560 2.820 3.050 3.220 ;
        RECT  2.810 0.620 3.050 3.220 ;
        RECT  5.940 1.580 6.340 1.820 ;
        RECT  2.560 1.480 3.050 1.720 ;
        RECT  2.810 0.620 6.260 0.860 ;
        RECT  1.930 3.460 4.510 3.700 ;
        RECT  4.270 1.580 4.510 3.700 ;
        RECT  1.320 3.250 1.560 3.650 ;
        RECT  1.320 3.250 2.170 3.490 ;
        RECT  1.930 1.480 2.170 3.700 ;
        RECT  4.110 2.910 4.510 3.150 ;
        RECT  1.930 2.150 2.570 2.550 ;
        RECT  4.110 1.580 4.510 1.820 ;
        RECT  1.320 1.480 2.170 1.720 ;
        RECT  0.820 4.000 3.440 4.240 ;
        RECT  0.450 3.760 1.060 4.000 ;
        RECT  0.820 1.280 1.060 4.240 ;
        RECT  0.600 1.280 1.060 1.520 ;
    END
END XNR3T

MACRO XNR4
    CLASS CORE ;
    FOREIGN XNR4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 0.620 9.750 3.300 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.450 2.740 ;
        RECT  0.120 2.280 0.580 2.740 ;
        RECT  0.120 3.910 2.910 4.150 ;
        RECT  4.110 3.910 4.510 4.320 ;
        RECT  2.670 4.080 4.510 4.320 ;
        RECT  0.120 2.280 0.360 4.150 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.940 1.690 2.740 ;
        RECT  1.300 1.940 1.690 2.340 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.300 2.280 14.760 2.740 ;
        RECT  14.520 2.280 14.760 4.240 ;
        RECT  11.770 4.000 14.760 4.240 ;
        RECT  11.770 4.000 12.170 4.340 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.940 13.580 2.340 ;
        RECT  13.190 1.940 13.470 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 0.560 ;
        RECT  7.870 -0.380 8.830 0.560 ;
        RECT  12.460 -0.380 12.860 0.560 ;
        RECT  14.030 -0.380 14.430 0.560 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  0.440 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 4.480 2.060 5.420 ;
        RECT  7.310 4.200 7.710 5.420 ;
        RECT  8.850 4.150 9.250 5.420 ;
        RECT  12.480 4.480 12.880 5.420 ;
        RECT  14.040 4.480 14.440 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  14.040 2.980 14.280 3.380 ;
        RECT  13.820 1.760 14.060 3.220 ;
        RECT  13.820 1.760 14.360 2.000 ;
        RECT  14.120 0.800 14.360 2.000 ;
        RECT  11.620 0.800 14.360 1.040 ;
        RECT  11.620 0.740 12.020 1.040 ;
        RECT  10.490 3.430 13.640 3.670 ;
        RECT  12.710 1.280 12.950 3.670 ;
        RECT  10.490 1.200 10.730 3.670 ;
        RECT  10.480 2.670 10.730 3.070 ;
        RECT  12.310 1.760 12.950 2.160 ;
        RECT  12.710 1.280 13.720 1.520 ;
        RECT  11.920 2.380 12.160 3.070 ;
        RECT  11.830 1.280 12.070 2.620 ;
        RECT  11.830 1.280 12.250 1.520 ;
        RECT  8.750 3.660 10.230 3.900 ;
        RECT  9.990 0.620 10.230 3.900 ;
        RECT  8.750 2.610 8.990 3.900 ;
        RECT  8.330 2.610 8.990 3.010 ;
        RECT  11.010 2.750 11.520 2.990 ;
        RECT  11.010 0.620 11.250 2.990 ;
        RECT  11.010 1.280 11.530 1.520 ;
        RECT  9.990 0.620 11.250 0.860 ;
        RECT  5.990 2.760 6.390 3.000 ;
        RECT  6.070 0.740 6.310 3.000 ;
        RECT  8.820 0.800 9.060 2.330 ;
        RECT  7.350 0.800 9.060 1.040 ;
        RECT  6.070 0.740 7.590 0.980 ;
        RECT  4.870 3.720 8.070 3.960 ;
        RECT  7.830 1.280 8.070 3.960 ;
        RECT  4.870 1.100 5.110 3.960 ;
        RECT  7.830 3.300 8.510 3.540 ;
        RECT  7.830 1.280 8.560 1.520 ;
        RECT  4.810 1.100 5.110 1.500 ;
        RECT  5.350 3.240 7.590 3.480 ;
        RECT  7.350 1.870 7.590 3.480 ;
        RECT  5.350 2.340 5.590 3.480 ;
        RECT  3.340 2.630 3.930 2.870 ;
        RECT  3.690 0.620 3.930 2.870 ;
        RECT  5.590 1.140 5.830 2.580 ;
        RECT  7.260 1.870 7.590 2.270 ;
        RECT  5.350 0.620 5.590 1.540 ;
        RECT  3.350 1.180 3.930 1.420 ;
        RECT  3.690 0.620 5.590 0.860 ;
        RECT  6.710 2.760 7.110 3.000 ;
        RECT  6.780 1.220 7.020 3.000 ;
        RECT  6.710 1.220 7.110 1.460 ;
        RECT  1.930 3.430 4.430 3.670 ;
        RECT  4.190 1.100 4.430 3.670 ;
        RECT  1.930 1.280 2.170 3.670 ;
        RECT  1.320 2.980 1.560 3.380 ;
        RECT  1.320 2.980 2.170 3.220 ;
        RECT  4.190 2.550 4.520 2.950 ;
        RECT  1.930 1.850 2.570 2.250 ;
        RECT  1.320 1.280 2.170 1.520 ;
        RECT  4.190 1.100 4.510 1.500 ;
        RECT  0.600 2.980 1.060 3.380 ;
        RECT  0.820 0.800 1.060 3.380 ;
        RECT  0.680 1.200 1.060 1.600 ;
        RECT  0.820 0.800 2.980 1.040 ;
        RECT  2.740 0.620 3.440 0.860 ;
        RECT  2.560 2.790 3.050 3.190 ;
        RECT  2.810 1.280 3.050 3.190 ;
        RECT  2.560 1.280 3.050 1.520 ;
    END
END XNR4

MACRO XNR4P
    CLASS CORE ;
    FOREIGN XNR4P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 1.250 9.900 1.650 ;
        RECT  9.470 2.810 9.920 3.210 ;
        RECT  9.470 0.620 9.750 3.300 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.450 2.740 ;
        RECT  0.120 2.280 0.580 2.740 ;
        RECT  0.120 3.910 2.910 4.150 ;
        RECT  4.250 3.910 4.650 4.320 ;
        RECT  2.670 4.080 4.790 4.320 ;
        RECT  0.120 2.280 0.360 4.150 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.940 1.690 2.740 ;
        RECT  1.300 1.940 1.690 2.340 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.920 2.280 15.380 2.740 ;
        RECT  15.140 2.280 15.380 4.150 ;
        RECT  12.470 3.910 15.380 4.150 ;
        RECT  12.470 3.910 12.850 4.420 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 1.940 14.200 2.340 ;
        RECT  13.810 1.940 14.090 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 0.560 ;
        RECT  8.040 -0.380 9.000 0.560 ;
        RECT  10.470 -0.380 10.870 0.560 ;
        RECT  13.080 -0.380 13.480 0.560 ;
        RECT  14.650 -0.380 15.050 0.560 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.440 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 4.480 2.060 5.420 ;
        RECT  7.480 4.200 7.880 5.420 ;
        RECT  8.980 4.150 9.380 5.420 ;
        RECT  10.290 4.480 10.690 5.420 ;
        RECT  13.100 4.480 13.500 5.420 ;
        RECT  14.660 4.480 15.060 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  14.440 2.980 14.900 3.380 ;
        RECT  14.440 1.760 14.680 3.380 ;
        RECT  14.440 1.760 14.980 2.000 ;
        RECT  14.740 0.800 14.980 2.000 ;
        RECT  12.240 0.800 14.980 1.040 ;
        RECT  12.240 0.740 12.640 1.040 ;
        RECT  11.110 3.430 13.570 3.670 ;
        RECT  13.330 1.280 13.570 3.670 ;
        RECT  11.110 1.280 11.350 3.670 ;
        RECT  13.940 2.980 14.180 3.380 ;
        RECT  13.330 3.060 14.180 3.300 ;
        RECT  11.020 2.750 11.420 2.990 ;
        RECT  12.930 1.760 13.570 2.160 ;
        RECT  13.330 1.280 14.340 1.520 ;
        RECT  11.030 1.280 11.430 1.520 ;
        RECT  12.540 2.380 12.780 3.070 ;
        RECT  12.450 1.280 12.690 2.620 ;
        RECT  12.450 1.280 12.870 1.520 ;
        RECT  8.920 3.660 10.780 3.900 ;
        RECT  10.540 0.800 10.780 3.900 ;
        RECT  8.920 2.610 9.160 3.900 ;
        RECT  8.500 2.610 9.160 3.010 ;
        RECT  11.670 2.750 12.140 2.990 ;
        RECT  11.670 0.800 11.910 2.990 ;
        RECT  11.670 1.280 12.150 1.520 ;
        RECT  10.540 0.800 11.910 1.040 ;
        RECT  6.160 2.760 6.560 3.000 ;
        RECT  6.240 0.740 6.480 3.000 ;
        RECT  8.990 0.800 9.230 2.330 ;
        RECT  7.520 0.800 9.230 1.040 ;
        RECT  6.240 0.740 7.760 0.980 ;
        RECT  5.040 3.720 8.240 3.960 ;
        RECT  8.000 1.280 8.240 3.960 ;
        RECT  5.040 1.700 5.280 3.960 ;
        RECT  8.000 3.300 8.680 3.540 ;
        RECT  5.040 1.700 5.520 2.100 ;
        RECT  8.000 1.280 8.730 1.520 ;
        RECT  5.520 3.240 7.760 3.480 ;
        RECT  7.520 1.870 7.760 3.480 ;
        RECT  5.520 2.340 5.760 3.480 ;
        RECT  3.340 2.630 3.930 2.870 ;
        RECT  3.690 0.620 3.930 2.870 ;
        RECT  5.760 1.220 6.000 2.580 ;
        RECT  7.430 1.870 7.760 2.270 ;
        RECT  5.440 1.220 6.000 1.460 ;
        RECT  3.350 1.180 3.930 1.420 ;
        RECT  5.440 0.620 5.680 1.460 ;
        RECT  3.690 0.620 5.680 0.860 ;
        RECT  6.880 2.760 7.280 3.000 ;
        RECT  6.950 1.220 7.190 3.000 ;
        RECT  6.880 1.220 7.280 1.460 ;
        RECT  1.930 3.430 4.650 3.670 ;
        RECT  4.410 1.180 4.650 3.670 ;
        RECT  1.930 1.280 2.170 3.670 ;
        RECT  1.320 2.980 1.560 3.380 ;
        RECT  1.320 2.980 2.170 3.220 ;
        RECT  4.200 2.630 4.650 2.870 ;
        RECT  1.930 1.850 2.570 2.250 ;
        RECT  1.320 1.280 2.170 1.520 ;
        RECT  4.190 1.180 4.650 1.420 ;
        RECT  0.600 2.980 1.060 3.380 ;
        RECT  0.820 0.800 1.060 3.380 ;
        RECT  0.680 1.200 1.060 1.600 ;
        RECT  0.820 0.800 2.980 1.040 ;
        RECT  2.740 0.620 3.440 0.860 ;
        RECT  2.560 2.790 3.050 3.190 ;
        RECT  2.810 1.280 3.050 3.190 ;
        RECT  2.560 1.280 3.050 1.520 ;
    END
END XNR4P

MACRO XNR4S
    CLASS CORE ;
    FOREIGN XNR4S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 0.620 9.750 3.300 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.450 2.740 ;
        RECT  0.120 2.280 0.580 2.740 ;
        RECT  0.120 3.910 2.910 4.150 ;
        RECT  4.030 3.910 4.430 4.320 ;
        RECT  2.670 4.080 4.430 4.320 ;
        RECT  0.120 2.280 0.360 4.150 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.940 1.690 2.740 ;
        RECT  1.300 1.940 1.690 2.340 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.300 2.280 14.760 2.740 ;
        RECT  14.520 2.280 14.760 4.150 ;
        RECT  11.850 3.910 14.760 4.150 ;
        RECT  11.850 3.910 12.230 4.420 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.940 13.580 2.340 ;
        RECT  13.190 1.940 13.470 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 0.560 ;
        RECT  7.870 -0.380 8.830 0.560 ;
        RECT  12.460 -0.380 12.860 0.560 ;
        RECT  14.030 -0.380 14.430 0.560 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  0.440 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 4.480 2.060 5.420 ;
        RECT  7.310 4.200 7.710 5.420 ;
        RECT  8.850 4.150 9.250 5.420 ;
        RECT  12.480 4.480 12.880 5.420 ;
        RECT  14.040 4.480 14.440 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.820 2.980 14.280 3.380 ;
        RECT  13.820 1.760 14.060 3.380 ;
        RECT  13.820 1.760 14.360 2.000 ;
        RECT  14.120 0.800 14.360 2.000 ;
        RECT  11.460 0.800 14.360 1.040 ;
        RECT  11.460 0.740 11.860 1.040 ;
        RECT  10.490 3.430 12.950 3.670 ;
        RECT  12.710 1.280 12.950 3.670 ;
        RECT  10.490 1.200 10.730 3.670 ;
        RECT  13.320 2.980 13.560 3.380 ;
        RECT  12.710 3.060 13.560 3.300 ;
        RECT  10.480 2.670 10.730 3.070 ;
        RECT  12.310 1.760 12.950 2.160 ;
        RECT  12.710 1.280 13.720 1.520 ;
        RECT  11.920 2.380 12.160 3.070 ;
        RECT  11.830 1.280 12.070 2.620 ;
        RECT  11.830 1.280 12.250 1.520 ;
        RECT  8.750 3.660 10.230 3.900 ;
        RECT  9.990 0.720 10.230 3.900 ;
        RECT  8.750 2.610 8.990 3.900 ;
        RECT  8.320 2.610 8.990 3.010 ;
        RECT  10.970 2.750 11.520 2.990 ;
        RECT  10.970 0.720 11.210 2.990 ;
        RECT  10.970 1.280 11.530 1.520 ;
        RECT  9.990 0.720 11.210 0.960 ;
        RECT  5.990 2.760 6.390 3.000 ;
        RECT  6.070 0.740 6.310 3.000 ;
        RECT  8.820 0.800 9.060 1.810 ;
        RECT  7.350 0.800 9.060 1.040 ;
        RECT  6.070 0.740 7.590 0.980 ;
        RECT  4.870 3.720 8.070 3.960 ;
        RECT  7.830 1.280 8.070 3.960 ;
        RECT  4.870 1.100 5.110 3.960 ;
        RECT  7.830 3.300 8.500 3.540 ;
        RECT  7.830 1.280 8.560 1.520 ;
        RECT  4.810 1.100 5.110 1.500 ;
        RECT  5.350 3.240 7.590 3.480 ;
        RECT  7.350 1.870 7.590 3.480 ;
        RECT  5.350 0.620 5.590 3.480 ;
        RECT  3.340 2.630 3.930 2.870 ;
        RECT  3.690 0.620 3.930 2.870 ;
        RECT  7.260 1.870 7.590 2.270 ;
        RECT  3.350 1.180 3.930 1.420 ;
        RECT  3.690 0.620 5.590 0.860 ;
        RECT  6.710 2.760 7.110 3.000 ;
        RECT  6.780 1.220 7.020 3.000 ;
        RECT  6.710 1.220 7.110 1.460 ;
        RECT  1.930 3.430 4.440 3.670 ;
        RECT  4.200 1.100 4.440 3.670 ;
        RECT  1.930 1.280 2.170 3.670 ;
        RECT  1.320 2.980 1.560 3.380 ;
        RECT  1.320 2.980 2.170 3.220 ;
        RECT  4.200 2.630 4.600 2.870 ;
        RECT  1.930 1.850 2.570 2.250 ;
        RECT  1.320 1.280 2.170 1.520 ;
        RECT  4.200 1.100 4.510 1.500 ;
        RECT  0.600 2.980 1.060 3.380 ;
        RECT  0.820 0.800 1.060 3.380 ;
        RECT  0.680 1.200 1.060 1.600 ;
        RECT  0.820 0.800 2.980 1.040 ;
        RECT  2.740 0.620 3.440 0.860 ;
        RECT  2.560 2.790 3.050 3.190 ;
        RECT  2.810 1.280 3.050 3.190 ;
        RECT  2.560 1.280 3.050 1.520 ;
    END
END XNR4S

MACRO XNR4T
    CLASS CORE ;
    FOREIGN XNR4T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.350 1.330 10.970 1.570 ;
        RECT  9.360 2.890 10.970 3.130 ;
        RECT  10.730 1.250 10.970 1.650 ;
        RECT  10.730 2.810 10.970 3.210 ;
        RECT  10.090 1.330 10.370 3.130 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.450 2.740 ;
        RECT  0.120 2.280 0.580 2.740 ;
        RECT  0.120 3.910 2.910 4.150 ;
        RECT  3.870 3.910 4.270 4.320 ;
        RECT  2.670 4.080 4.410 4.320 ;
        RECT  0.120 2.280 0.360 4.150 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.940 1.690 2.740 ;
        RECT  1.300 1.940 1.690 2.340 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.540 2.280 16.000 2.740 ;
        RECT  15.760 2.280 16.000 4.150 ;
        RECT  13.090 3.910 16.000 4.150 ;
        RECT  13.090 3.910 13.470 4.420 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 1.940 14.820 2.340 ;
        RECT  14.430 1.940 14.710 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 0.560 ;
        RECT  7.870 -0.380 8.830 0.560 ;
        RECT  9.990 -0.380 10.390 0.780 ;
        RECT  13.700 -0.380 14.100 0.560 ;
        RECT  15.270 -0.380 15.670 0.560 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  0.440 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 4.480 2.060 5.420 ;
        RECT  7.310 4.200 7.710 5.420 ;
        RECT  8.740 4.150 9.140 5.420 ;
        RECT  10.010 4.150 10.410 5.420 ;
        RECT  13.720 4.480 14.120 5.420 ;
        RECT  15.280 4.480 15.680 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  15.060 2.980 15.520 3.380 ;
        RECT  15.060 1.760 15.300 3.380 ;
        RECT  15.060 1.760 15.600 2.000 ;
        RECT  15.360 0.800 15.600 2.000 ;
        RECT  12.710 0.800 15.600 1.040 ;
        RECT  12.710 0.740 13.110 1.040 ;
        RECT  11.730 3.430 14.190 3.670 ;
        RECT  13.950 1.280 14.190 3.670 ;
        RECT  11.730 1.200 11.970 3.670 ;
        RECT  14.560 2.980 14.800 3.380 ;
        RECT  13.950 3.060 14.800 3.300 ;
        RECT  11.720 2.670 11.970 3.070 ;
        RECT  13.550 1.760 14.190 2.160 ;
        RECT  13.950 1.280 14.960 1.520 ;
        RECT  13.160 2.380 13.400 3.070 ;
        RECT  13.070 1.280 13.310 2.620 ;
        RECT  13.070 1.280 13.490 1.520 ;
        RECT  8.750 3.660 11.450 3.900 ;
        RECT  11.210 0.720 11.450 3.900 ;
        RECT  8.750 2.610 8.990 3.900 ;
        RECT  8.320 2.610 8.990 3.010 ;
        RECT  12.220 2.750 12.760 2.990 ;
        RECT  12.220 0.720 12.460 2.990 ;
        RECT  12.220 1.280 12.770 1.520 ;
        RECT  11.210 0.720 12.460 0.960 ;
        RECT  5.990 2.760 6.390 3.000 ;
        RECT  6.070 0.740 6.310 3.000 ;
        RECT  8.820 0.800 9.060 2.330 ;
        RECT  7.350 0.800 9.060 1.040 ;
        RECT  6.070 0.740 7.590 0.980 ;
        RECT  4.870 3.720 8.070 3.960 ;
        RECT  7.830 1.280 8.070 3.960 ;
        RECT  4.870 1.100 5.110 3.960 ;
        RECT  7.830 3.300 8.500 3.540 ;
        RECT  7.830 1.280 8.490 1.520 ;
        RECT  4.810 1.100 5.110 1.500 ;
        RECT  5.350 3.240 7.590 3.480 ;
        RECT  7.350 1.870 7.590 3.480 ;
        RECT  5.350 0.620 5.590 3.480 ;
        RECT  3.340 2.630 3.930 2.870 ;
        RECT  3.690 0.620 3.930 2.870 ;
        RECT  7.260 1.870 7.590 2.270 ;
        RECT  3.350 1.180 3.930 1.420 ;
        RECT  3.690 0.620 5.590 0.860 ;
        RECT  6.710 2.760 7.110 3.000 ;
        RECT  6.780 1.220 7.020 3.000 ;
        RECT  6.710 1.220 7.110 1.460 ;
        RECT  1.930 3.430 4.440 3.670 ;
        RECT  4.200 1.100 4.440 3.670 ;
        RECT  1.930 1.280 2.170 3.670 ;
        RECT  1.320 2.980 1.560 3.380 ;
        RECT  1.320 2.980 2.170 3.220 ;
        RECT  4.200 2.550 4.520 2.950 ;
        RECT  1.930 1.850 2.570 2.250 ;
        RECT  1.320 1.280 2.170 1.520 ;
        RECT  4.200 1.100 4.510 1.500 ;
        RECT  0.600 2.980 1.060 3.380 ;
        RECT  0.820 0.800 1.060 3.380 ;
        RECT  0.680 1.200 1.060 1.600 ;
        RECT  0.820 0.800 2.980 1.040 ;
        RECT  2.740 0.620 3.440 0.860 ;
        RECT  2.560 2.790 3.050 3.190 ;
        RECT  2.810 1.280 3.050 3.190 ;
        RECT  2.560 1.280 3.050 1.520 ;
    END
END XNR4T

MACRO XOR2H
    CLASS CORE ;
    FOREIGN XOR2H 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.390 1.570 6.630 3.110 ;
        RECT  3.120 2.870 6.630 3.110 ;
        RECT  3.190 1.570 6.630 1.810 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 2.110 2.650 ;
        RECT  1.410 2.250 1.690 2.890 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.250 0.690 2.650 ;
        RECT  0.170 2.250 0.450 2.890 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 -0.380 2.070 0.560 ;
        RECT  6.670 -0.380 7.070 0.780 ;
        RECT  8.120 -0.380 8.520 0.780 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  6.510 4.310 6.910 5.420 ;
        RECT  8.120 4.260 8.520 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.840 4.110 6.270 4.350 ;
        RECT  6.030 3.830 6.270 4.350 ;
        RECT  6.030 3.830 7.720 4.070 ;
        RECT  7.480 1.020 7.720 4.070 ;
        RECT  5.350 1.020 7.720 1.260 ;
        RECT  0.930 3.780 3.600 4.020 ;
        RECT  3.360 3.350 3.600 4.020 ;
        RECT  0.930 3.620 1.200 4.020 ;
        RECT  0.930 0.800 1.170 4.020 ;
        RECT  3.360 3.350 7.240 3.590 ;
        RECT  7.000 2.250 7.240 3.590 ;
        RECT  0.930 0.800 1.200 1.200 ;
        RECT  0.930 0.800 4.310 1.040 ;
        RECT  2.470 1.570 2.710 3.390 ;
        RECT  2.470 2.330 5.680 2.570 ;
        RECT  2.460 1.570 2.860 1.810 ;
    END
END XOR2H

MACRO XOR2HP
    CLASS CORE ;
    FOREIGN XOR2HP 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.490 2.870 11.670 3.110 ;
        RECT  5.620 1.570 11.800 1.810 ;
        RECT  11.330 1.570 11.610 3.110 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.250 3.550 2.890 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.250 1.690 2.890 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.110 -0.380 3.510 0.560 ;
        RECT  4.830 -0.380 5.230 0.560 ;
        RECT  12.050 -0.380 12.450 0.780 ;
        RECT  13.500 -0.380 13.900 0.780 ;
        RECT  14.940 -0.380 15.340 0.780 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.760 4.260 5.160 5.420 ;
        RECT  11.890 4.310 12.290 5.420 ;
        RECT  13.500 4.260 13.900 5.420 ;
        RECT  14.940 4.260 15.340 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.210 4.110 11.540 4.350 ;
        RECT  11.300 3.830 11.540 4.350 ;
        RECT  11.300 3.830 13.180 4.070 ;
        RECT  14.380 1.090 14.620 4.020 ;
        RECT  12.860 3.780 14.620 4.020 ;
        RECT  9.220 1.090 14.620 1.330 ;
        RECT  0.880 3.780 5.940 4.020 ;
        RECT  5.700 3.350 5.940 4.020 ;
        RECT  2.400 1.190 2.640 4.020 ;
        RECT  5.700 3.350 12.420 3.590 ;
        RECT  12.180 2.410 12.420 3.590 ;
        RECT  12.180 2.410 13.960 2.650 ;
        RECT  13.220 2.250 13.960 2.650 ;
        RECT  0.880 1.190 3.620 1.430 ;
        RECT  3.380 1.090 8.180 1.330 ;
        RECT  3.900 2.890 5.250 3.130 ;
        RECT  5.010 1.570 5.250 3.130 ;
        RECT  5.010 2.330 9.760 2.570 ;
        RECT  3.900 1.570 5.250 1.810 ;
    END
END XOR2HP

MACRO XOR2HS
    CLASS CORE ;
    FOREIGN XOR2HS 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.950 1.840 4.150 2.080 ;
        RECT  3.910 1.840 4.150 3.110 ;
        RECT  2.880 2.870 4.150 3.110 ;
        RECT  2.950 1.540 3.350 2.080 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.010 1.690 2.750 ;
        RECT  1.330 2.250 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.070 2.890 ;
        RECT  0.650 2.250 1.070 2.650 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.230 -0.380 4.630 0.620 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  1.020 -0.380 1.420 0.810 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.130 4.480 4.530 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.880 4.260 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.160 4.110 3.890 4.350 ;
        RECT  3.650 3.830 3.890 4.350 ;
        RECT  3.650 3.830 5.340 4.070 ;
        RECT  5.100 1.340 5.340 4.070 ;
        RECT  3.670 1.340 5.340 1.580 ;
        RECT  0.170 3.630 2.870 3.870 ;
        RECT  2.630 3.350 2.870 3.870 ;
        RECT  0.170 3.470 0.480 3.870 ;
        RECT  2.630 3.350 4.780 3.590 ;
        RECT  4.540 2.250 4.780 3.590 ;
        RECT  0.170 1.050 0.410 3.870 ;
        RECT  0.170 1.050 0.480 1.450 ;
        RECT  0.170 1.050 2.630 1.290 ;
        RECT  2.100 0.680 2.630 1.290 ;
        RECT  1.560 2.990 2.170 3.390 ;
        RECT  1.930 1.530 2.170 3.390 ;
        RECT  1.930 2.330 3.540 2.570 ;
        RECT  1.530 1.530 2.170 1.770 ;
    END
END XOR2HS

MACRO XOR2HT
    CLASS CORE ;
    FOREIGN XOR2HT 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.320 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.710 2.870 16.750 3.110 ;
        RECT  7.790 1.570 16.830 1.810 ;
        RECT  16.290 1.570 16.570 3.110 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.250 5.410 2.650 ;
        RECT  4.510 2.250 4.790 3.130 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.250 2.310 3.130 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  3.040 -0.380 3.440 0.950 ;
        RECT  4.550 -0.380 4.950 0.560 ;
        RECT  6.270 -0.380 6.670 0.560 ;
        RECT  17.420 -0.380 17.820 0.850 ;
        RECT  18.880 -0.380 19.280 0.780 ;
        RECT  20.320 -0.380 20.730 0.780 ;
        RECT  21.760 -0.380 22.160 0.780 ;
        RECT  0.000 -0.380 22.320 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.260 2.000 5.420 ;
        RECT  3.040 4.260 3.440 5.420 ;
        RECT  4.480 4.260 4.880 5.420 ;
        RECT  6.200 4.260 6.600 5.420 ;
        RECT  17.360 4.310 17.760 5.420 ;
        RECT  18.880 4.260 19.280 5.420 ;
        RECT  20.320 4.260 20.720 5.420 ;
        RECT  21.760 4.260 22.160 5.420 ;
        RECT  0.000 4.660 22.320 5.420 ;
        RECT  0.160 4.260 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.430 4.110 16.560 4.350 ;
        RECT  16.320 3.830 16.560 4.350 ;
        RECT  16.320 3.830 18.560 4.070 ;
        RECT  21.200 1.090 21.440 4.020 ;
        RECT  18.240 3.780 21.440 4.020 ;
        RECT  12.830 1.090 21.440 1.330 ;
        RECT  0.880 3.780 8.160 4.020 ;
        RECT  7.920 3.350 8.160 4.020 ;
        RECT  3.840 1.190 4.080 4.020 ;
        RECT  7.920 3.350 17.270 3.590 ;
        RECT  17.030 2.130 17.270 3.590 ;
        RECT  17.030 2.130 20.150 2.370 ;
        RECT  19.410 1.970 20.150 2.370 ;
        RECT  0.880 1.190 5.060 1.430 ;
        RECT  4.820 1.090 11.790 1.330 ;
        RECT  5.340 2.890 7.390 3.130 ;
        RECT  7.150 1.570 7.390 3.130 ;
        RECT  7.150 2.330 14.820 2.570 ;
        RECT  5.340 1.570 7.460 1.810 ;
    END
END XOR2HT

MACRO XOR3
    CLASS CORE ;
    FOREIGN XOR3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.710 1.180 10.990 3.300 ;
        RECT  10.680 2.900 10.990 3.300 ;
        RECT  10.680 1.180 10.990 1.580 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.280 0.580 2.680 ;
        RECT  0.170 2.170 0.450 2.870 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.720 2.520 ;
        RECT  1.410 2.120 1.690 2.990 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 2.300 9.750 3.020 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.050 -0.380 2.450 1.060 ;
        RECT  9.300 -0.380 10.200 0.560 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.450 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.030 4.480 2.430 5.420 ;
        RECT  9.700 4.480 10.100 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.740 0.830 7.980 3.300 ;
        RECT  10.200 2.030 10.460 2.430 ;
        RECT  10.200 0.830 10.440 2.430 ;
        RECT  7.740 0.830 10.440 1.070 ;
        RECT  8.990 3.320 9.520 3.720 ;
        RECT  8.990 1.870 9.230 3.720 ;
        RECT  9.020 1.330 9.260 2.110 ;
        RECT  9.020 1.330 9.550 1.570 ;
        RECT  4.930 4.180 8.700 4.420 ;
        RECT  8.460 1.330 8.700 4.420 ;
        RECT  4.930 1.100 5.170 4.420 ;
        RECT  3.520 2.910 3.950 3.150 ;
        RECT  3.710 1.100 3.950 3.150 ;
        RECT  3.530 1.580 3.950 1.820 ;
        RECT  8.380 1.330 8.780 1.570 ;
        RECT  3.710 1.100 5.170 1.340 ;
        RECT  5.410 3.470 7.260 3.710 ;
        RECT  7.020 1.250 7.260 3.710 ;
        RECT  5.410 1.500 5.650 3.710 ;
        RECT  6.200 0.620 6.440 3.230 ;
        RECT  2.810 2.830 3.230 3.230 ;
        RECT  2.990 0.620 3.230 3.230 ;
        RECT  6.120 1.580 6.520 1.820 ;
        RECT  2.740 1.480 3.230 1.720 ;
        RECT  2.990 0.620 6.440 0.860 ;
        RECT  2.110 3.470 4.690 3.710 ;
        RECT  4.450 1.580 4.690 3.710 ;
        RECT  1.410 3.250 1.650 3.650 ;
        RECT  1.410 3.250 2.350 3.490 ;
        RECT  2.110 1.480 2.350 3.710 ;
        RECT  4.290 2.910 4.690 3.150 ;
        RECT  2.110 2.150 2.750 2.550 ;
        RECT  4.290 1.580 4.690 1.820 ;
        RECT  1.360 1.480 2.350 1.720 ;
        RECT  0.820 4.000 3.620 4.240 ;
        RECT  0.450 3.760 1.060 4.000 ;
        RECT  0.820 1.280 1.060 4.240 ;
        RECT  0.600 1.280 1.060 1.520 ;
    END
END XOR3

MACRO XOR3P
    CLASS CORE ;
    FOREIGN XOR3P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.710 1.180 10.990 3.300 ;
        RECT  10.580 2.900 10.990 3.300 ;
        RECT  10.580 1.180 10.990 1.580 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.280 0.580 2.680 ;
        RECT  0.170 2.170 0.450 2.870 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.720 2.520 ;
        RECT  1.410 2.120 1.690 2.990 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 2.300 9.750 3.020 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.050 -0.380 2.450 1.060 ;
        RECT  9.200 -0.380 10.100 0.560 ;
        RECT  11.220 -0.380 11.620 0.950 ;
        RECT  0.000 -0.380 11.780 0.380 ;
        RECT  0.450 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.030 4.480 2.430 5.420 ;
        RECT  9.600 4.480 10.000 5.420 ;
        RECT  11.220 4.260 11.620 5.420 ;
        RECT  0.000 4.660 11.780 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.740 0.830 7.980 3.300 ;
        RECT  10.100 2.030 10.460 2.430 ;
        RECT  10.100 0.830 10.340 2.430 ;
        RECT  7.740 0.830 10.340 1.070 ;
        RECT  8.990 3.320 9.520 3.720 ;
        RECT  8.990 1.870 9.230 3.720 ;
        RECT  9.020 1.330 9.260 2.110 ;
        RECT  9.020 1.330 9.500 1.570 ;
        RECT  4.930 4.180 8.700 4.420 ;
        RECT  8.460 1.330 8.700 4.420 ;
        RECT  4.930 1.100 5.170 4.420 ;
        RECT  3.520 2.910 3.950 3.150 ;
        RECT  3.710 1.100 3.950 3.150 ;
        RECT  3.530 1.580 3.950 1.820 ;
        RECT  8.380 1.330 8.780 1.570 ;
        RECT  3.710 1.100 5.170 1.340 ;
        RECT  5.410 3.470 7.260 3.710 ;
        RECT  7.020 1.250 7.260 3.710 ;
        RECT  5.410 1.500 5.650 3.710 ;
        RECT  6.200 0.620 6.440 3.230 ;
        RECT  2.810 2.830 3.230 3.230 ;
        RECT  2.990 0.620 3.230 3.230 ;
        RECT  6.120 1.580 6.520 1.820 ;
        RECT  2.740 1.480 3.230 1.720 ;
        RECT  2.990 0.620 6.440 0.860 ;
        RECT  2.110 3.470 4.690 3.710 ;
        RECT  4.450 1.580 4.690 3.710 ;
        RECT  1.410 3.250 1.650 3.650 ;
        RECT  1.410 3.250 2.350 3.490 ;
        RECT  2.110 1.480 2.350 3.710 ;
        RECT  4.290 2.910 4.690 3.150 ;
        RECT  2.110 2.150 2.750 2.550 ;
        RECT  4.290 1.580 4.690 1.820 ;
        RECT  1.360 1.480 2.350 1.720 ;
        RECT  0.820 4.000 3.620 4.240 ;
        RECT  0.450 3.760 1.060 4.000 ;
        RECT  0.820 1.280 1.060 4.240 ;
        RECT  0.600 1.280 1.060 1.520 ;
    END
END XOR3P

MACRO XOR3S
    CLASS CORE ;
    FOREIGN XOR3S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.710 1.230 10.990 3.820 ;
        RECT  10.680 3.420 10.990 3.820 ;
        RECT  10.680 1.230 10.990 1.630 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.280 0.580 2.680 ;
        RECT  0.170 2.170 0.450 2.870 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.720 2.520 ;
        RECT  1.410 2.120 1.690 2.990 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 2.300 9.750 3.020 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.050 -0.380 2.450 0.960 ;
        RECT  9.300 -0.380 10.200 0.560 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  0.450 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.030 4.480 2.430 5.420 ;
        RECT  9.770 4.340 10.170 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.740 0.830 7.980 3.300 ;
        RECT  10.200 2.030 10.460 2.430 ;
        RECT  10.200 0.830 10.440 2.430 ;
        RECT  7.740 0.830 10.440 1.070 ;
        RECT  8.990 3.320 9.520 3.720 ;
        RECT  8.990 1.870 9.230 3.720 ;
        RECT  9.020 1.330 9.260 2.110 ;
        RECT  9.020 1.330 9.540 1.570 ;
        RECT  4.930 4.180 8.700 4.420 ;
        RECT  8.460 1.330 8.700 4.420 ;
        RECT  4.930 1.100 5.170 4.420 ;
        RECT  3.520 2.910 3.950 3.150 ;
        RECT  3.710 1.100 3.950 3.150 ;
        RECT  3.530 1.580 3.950 1.820 ;
        RECT  8.380 1.330 8.780 1.570 ;
        RECT  3.710 1.100 5.170 1.340 ;
        RECT  5.410 3.470 7.260 3.710 ;
        RECT  7.020 1.250 7.260 3.710 ;
        RECT  5.410 1.500 5.650 3.710 ;
        RECT  6.200 0.620 6.440 3.230 ;
        RECT  2.810 2.830 3.230 3.230 ;
        RECT  2.990 0.620 3.230 3.230 ;
        RECT  6.120 1.580 6.520 1.820 ;
        RECT  2.740 1.480 3.230 1.720 ;
        RECT  2.990 0.620 6.440 0.860 ;
        RECT  1.330 3.520 4.690 3.760 ;
        RECT  4.450 1.580 4.690 3.760 ;
        RECT  2.110 1.480 2.350 3.760 ;
        RECT  4.290 2.910 4.690 3.150 ;
        RECT  2.110 2.150 2.750 2.550 ;
        RECT  4.290 1.580 4.690 1.820 ;
        RECT  1.360 1.480 2.350 1.720 ;
        RECT  0.820 4.000 3.620 4.240 ;
        RECT  0.450 3.760 1.060 4.000 ;
        RECT  0.820 1.280 1.060 4.240 ;
        RECT  0.600 1.280 1.060 1.520 ;
    END
END XOR3S

MACRO XOR3T
    CLASS CORE ;
    FOREIGN XOR3T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.330 1.260 11.610 3.220 ;
        RECT  10.480 1.260 12.240 1.540 ;
        RECT  10.400 2.940 12.240 3.220 ;
        RECT  10.480 1.260 10.720 1.660 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.280 0.580 2.680 ;
        RECT  0.170 2.170 0.450 2.870 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.120 1.700 2.520 ;
        RECT  1.410 2.120 1.690 2.990 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.400 2.620 9.750 3.020 ;
        RECT  9.470 2.300 9.750 3.020 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.030 -0.380 2.430 1.060 ;
        RECT  9.100 -0.380 10.000 0.560 ;
        RECT  11.120 -0.380 11.520 0.950 ;
        RECT  0.000 -0.380 12.400 0.380 ;
        RECT  0.450 -0.380 0.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.010 4.480 2.410 5.420 ;
        RECT  9.500 4.480 9.900 5.420 ;
        RECT  11.120 4.260 11.520 5.420 ;
        RECT  0.000 4.660 12.400 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.720 0.830 7.960 3.300 ;
        RECT  10.000 2.030 10.360 2.430 ;
        RECT  10.000 0.830 10.240 2.430 ;
        RECT  7.720 0.830 10.240 1.070 ;
        RECT  8.920 3.400 9.480 3.640 ;
        RECT  8.920 1.870 9.160 3.640 ;
        RECT  8.920 1.870 9.210 2.340 ;
        RECT  9.000 1.330 9.240 2.110 ;
        RECT  9.000 1.330 9.480 1.570 ;
        RECT  4.910 4.180 8.680 4.420 ;
        RECT  8.440 1.330 8.680 4.420 ;
        RECT  4.910 1.100 5.150 4.420 ;
        RECT  3.500 2.910 3.930 3.150 ;
        RECT  3.690 1.100 3.930 3.150 ;
        RECT  3.510 1.580 3.930 1.820 ;
        RECT  8.360 1.330 8.760 1.570 ;
        RECT  3.690 1.100 5.150 1.340 ;
        RECT  5.390 3.470 7.240 3.710 ;
        RECT  7.000 1.250 7.240 3.710 ;
        RECT  5.390 1.500 5.630 3.710 ;
        RECT  6.180 0.620 6.420 3.230 ;
        RECT  2.790 2.830 3.210 3.230 ;
        RECT  2.970 0.620 3.210 3.230 ;
        RECT  6.100 1.580 6.500 1.820 ;
        RECT  2.720 1.480 3.210 1.720 ;
        RECT  2.970 0.620 6.420 0.860 ;
        RECT  2.090 3.470 4.670 3.710 ;
        RECT  4.430 1.580 4.670 3.710 ;
        RECT  1.390 3.250 1.630 3.650 ;
        RECT  1.390 3.250 2.330 3.490 ;
        RECT  2.090 1.480 2.330 3.710 ;
        RECT  4.270 2.910 4.670 3.150 ;
        RECT  2.090 2.150 2.730 2.550 ;
        RECT  4.270 1.580 4.670 1.820 ;
        RECT  1.340 1.480 2.330 1.720 ;
        RECT  0.820 4.000 3.600 4.240 ;
        RECT  0.450 3.760 1.060 4.000 ;
        RECT  0.820 1.280 1.060 4.240 ;
        RECT  0.600 1.280 1.060 1.520 ;
    END
END XOR3T

MACRO XOR4
    CLASS CORE ;
    FOREIGN XOR4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.460 2.810 9.750 3.210 ;
        RECT  9.470 0.620 9.750 3.300 ;
        RECT  9.440 1.250 9.750 1.650 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.450 2.740 ;
        RECT  0.120 2.280 0.580 2.740 ;
        RECT  0.120 3.910 2.910 4.150 ;
        RECT  4.030 3.910 4.430 4.320 ;
        RECT  2.670 4.080 4.430 4.320 ;
        RECT  0.120 2.280 0.360 4.150 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.940 1.690 2.740 ;
        RECT  1.300 1.940 1.690 2.340 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 2.130 14.760 2.740 ;
        RECT  14.300 2.280 14.760 2.740 ;
        RECT  14.520 2.130 14.760 4.240 ;
        RECT  11.850 4.000 14.760 4.240 ;
        RECT  11.850 4.000 12.090 4.420 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.940 13.580 2.340 ;
        RECT  13.190 1.940 13.470 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 0.560 ;
        RECT  7.840 -0.380 8.800 0.560 ;
        RECT  12.370 -0.380 12.770 0.560 ;
        RECT  14.030 -0.380 14.430 0.560 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  0.440 -0.380 0.840 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 4.480 2.060 5.420 ;
        RECT  7.280 4.200 7.680 5.420 ;
        RECT  8.820 4.150 9.220 5.420 ;
        RECT  12.480 4.480 12.880 5.420 ;
        RECT  13.790 4.480 14.190 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.820 3.130 14.280 3.530 ;
        RECT  13.820 1.760 14.060 3.530 ;
        RECT  13.890 0.800 14.130 2.000 ;
        RECT  13.890 1.200 14.360 1.600 ;
        RECT  11.460 0.800 14.130 1.040 ;
        RECT  11.460 0.620 11.860 1.040 ;
        RECT  10.490 3.430 12.950 3.670 ;
        RECT  12.710 1.280 12.950 3.670 ;
        RECT  10.490 1.200 10.730 3.670 ;
        RECT  13.320 2.980 13.560 3.380 ;
        RECT  12.710 3.060 13.560 3.300 ;
        RECT  10.480 2.670 10.730 3.070 ;
        RECT  12.310 1.760 12.950 2.160 ;
        RECT  12.710 1.280 13.650 1.520 ;
        RECT  11.920 2.380 12.160 3.070 ;
        RECT  11.830 1.280 12.070 2.620 ;
        RECT  11.830 1.280 12.250 1.520 ;
        RECT  8.720 3.660 10.230 3.900 ;
        RECT  9.990 0.620 10.230 3.900 ;
        RECT  8.720 2.610 8.960 3.900 ;
        RECT  8.300 2.610 8.960 3.010 ;
        RECT  10.970 2.750 11.520 2.990 ;
        RECT  10.970 0.620 11.210 2.990 ;
        RECT  10.970 1.280 11.530 1.520 ;
        RECT  9.990 0.620 11.210 0.860 ;
        RECT  5.960 2.740 6.360 2.980 ;
        RECT  6.040 0.740 6.280 2.980 ;
        RECT  8.790 0.800 9.030 2.330 ;
        RECT  7.320 0.800 9.030 1.040 ;
        RECT  6.040 0.740 7.560 0.980 ;
        RECT  5.730 3.700 8.040 3.940 ;
        RECT  7.800 1.280 8.040 3.940 ;
        RECT  7.800 3.300 8.480 3.540 ;
        RECT  7.800 1.280 8.460 1.520 ;
        RECT  5.320 0.620 5.560 3.480 ;
        RECT  5.320 3.220 7.560 3.460 ;
        RECT  7.320 1.870 7.560 3.460 ;
        RECT  3.340 2.630 3.920 2.870 ;
        RECT  3.680 0.620 3.920 2.870 ;
        RECT  7.230 1.870 7.560 2.270 ;
        RECT  3.350 1.180 3.920 1.420 ;
        RECT  3.680 0.620 5.560 0.860 ;
        RECT  6.680 2.740 7.080 2.980 ;
        RECT  6.750 1.220 6.990 2.980 ;
        RECT  6.680 1.220 7.080 1.460 ;
        RECT  4.840 4.180 6.850 4.420 ;
        RECT  4.840 1.100 5.080 4.420 ;
        RECT  4.780 1.100 5.080 1.500 ;
        RECT  1.930 3.430 4.520 3.670 ;
        RECT  4.280 1.100 4.520 3.670 ;
        RECT  1.930 1.280 2.170 3.670 ;
        RECT  1.320 2.980 1.560 3.380 ;
        RECT  1.320 2.980 2.170 3.220 ;
        RECT  1.930 1.850 2.570 2.250 ;
        RECT  1.320 1.280 2.170 1.520 ;
        RECT  4.240 1.100 4.520 1.500 ;
        RECT  0.600 2.980 1.060 3.380 ;
        RECT  0.820 0.800 1.060 3.380 ;
        RECT  0.680 1.200 1.060 1.600 ;
        RECT  0.820 0.800 2.980 1.040 ;
        RECT  2.740 0.620 3.440 0.860 ;
        RECT  2.560 2.790 3.050 3.190 ;
        RECT  2.810 1.280 3.050 3.190 ;
        RECT  2.560 1.280 3.050 1.520 ;
    END
END XOR4

MACRO XOR4P
    CLASS CORE ;
    FOREIGN XOR4P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.500 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.470 1.250 9.880 1.650 ;
        RECT  9.470 2.810 9.890 3.210 ;
        RECT  9.470 0.620 9.750 3.300 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.450 2.740 ;
        RECT  0.120 2.280 0.580 2.740 ;
        RECT  0.120 3.910 2.910 4.150 ;
        RECT  4.250 3.910 4.650 4.320 ;
        RECT  2.670 4.080 4.650 4.320 ;
        RECT  0.120 2.280 0.360 4.150 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.940 1.690 2.740 ;
        RECT  1.300 1.940 1.690 2.340 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.050 2.130 15.380 2.740 ;
        RECT  14.920 2.280 15.380 2.740 ;
        RECT  15.140 2.130 15.380 4.240 ;
        RECT  12.470 4.000 15.380 4.240 ;
        RECT  12.470 4.000 12.710 4.420 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.810 1.940 14.200 2.340 ;
        RECT  13.810 1.940 14.090 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 0.560 ;
        RECT  8.040 -0.380 9.000 0.560 ;
        RECT  10.450 -0.380 10.850 0.560 ;
        RECT  12.990 -0.380 13.390 0.560 ;
        RECT  14.650 -0.380 15.050 0.560 ;
        RECT  0.000 -0.380 15.500 0.380 ;
        RECT  0.440 -0.380 0.840 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 4.480 2.060 5.420 ;
        RECT  7.480 4.200 7.880 5.420 ;
        RECT  8.960 4.150 9.360 5.420 ;
        RECT  10.270 4.390 10.670 5.420 ;
        RECT  13.100 4.480 13.500 5.420 ;
        RECT  14.410 4.480 14.810 5.420 ;
        RECT  0.000 4.660 15.500 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  14.440 3.130 14.900 3.530 ;
        RECT  14.440 1.760 14.680 3.530 ;
        RECT  14.510 0.800 14.750 2.000 ;
        RECT  14.510 1.200 14.980 1.600 ;
        RECT  12.150 0.800 14.750 1.040 ;
        RECT  12.150 0.620 12.550 1.040 ;
        RECT  11.110 3.430 13.570 3.670 ;
        RECT  13.330 1.280 13.570 3.670 ;
        RECT  11.110 1.280 11.350 3.670 ;
        RECT  13.940 2.980 14.180 3.380 ;
        RECT  13.330 3.060 14.180 3.300 ;
        RECT  11.100 2.670 11.350 3.070 ;
        RECT  12.930 1.760 13.570 2.160 ;
        RECT  13.330 1.280 14.270 1.520 ;
        RECT  11.030 1.280 11.430 1.520 ;
        RECT  12.540 2.380 12.780 3.070 ;
        RECT  12.450 1.280 12.690 2.620 ;
        RECT  12.450 1.280 12.870 1.520 ;
        RECT  8.920 3.660 10.790 3.900 ;
        RECT  10.550 0.800 10.790 3.900 ;
        RECT  8.920 2.610 9.160 3.900 ;
        RECT  8.490 2.610 9.160 3.010 ;
        RECT  11.670 2.750 12.140 2.990 ;
        RECT  11.670 0.800 11.910 2.990 ;
        RECT  11.670 1.280 12.150 1.520 ;
        RECT  10.550 0.800 11.910 1.040 ;
        RECT  6.160 2.740 6.560 2.980 ;
        RECT  6.240 0.740 6.480 2.980 ;
        RECT  8.990 0.800 9.230 2.330 ;
        RECT  7.520 0.800 9.230 1.040 ;
        RECT  6.240 0.740 7.760 0.980 ;
        RECT  5.930 3.700 8.240 3.940 ;
        RECT  8.000 1.280 8.240 3.940 ;
        RECT  8.000 3.300 8.670 3.540 ;
        RECT  8.000 1.280 8.660 1.520 ;
        RECT  5.520 2.320 5.760 3.480 ;
        RECT  5.520 3.220 7.760 3.460 ;
        RECT  7.520 1.870 7.760 3.460 ;
        RECT  3.340 2.630 3.920 2.870 ;
        RECT  3.680 0.620 3.920 2.870 ;
        RECT  5.760 1.220 6.000 2.560 ;
        RECT  7.430 1.870 7.760 2.270 ;
        RECT  5.440 1.220 6.000 1.460 ;
        RECT  3.350 1.180 3.920 1.420 ;
        RECT  5.440 0.620 5.680 1.460 ;
        RECT  3.680 0.620 5.680 0.860 ;
        RECT  6.880 2.740 7.280 2.980 ;
        RECT  6.950 1.220 7.190 2.980 ;
        RECT  6.880 1.220 7.280 1.460 ;
        RECT  5.040 4.180 7.050 4.420 ;
        RECT  5.040 1.760 5.280 4.420 ;
        RECT  5.040 1.760 5.520 2.000 ;
        RECT  1.930 3.430 4.650 3.670 ;
        RECT  4.410 1.180 4.650 3.670 ;
        RECT  1.930 1.280 2.170 3.670 ;
        RECT  1.320 2.980 1.560 3.380 ;
        RECT  1.320 2.980 2.170 3.220 ;
        RECT  4.200 2.630 4.650 2.870 ;
        RECT  1.930 1.850 2.570 2.250 ;
        RECT  1.320 1.280 2.170 1.520 ;
        RECT  4.160 1.180 4.650 1.420 ;
        RECT  0.600 2.980 1.060 3.380 ;
        RECT  0.820 0.800 1.060 3.380 ;
        RECT  0.680 1.200 1.060 1.600 ;
        RECT  0.820 0.800 2.980 1.040 ;
        RECT  2.740 0.620 3.440 0.860 ;
        RECT  2.560 2.790 3.050 3.190 ;
        RECT  2.810 1.280 3.050 3.190 ;
        RECT  2.560 1.280 3.050 1.520 ;
    END
END XOR4P

MACRO XOR4S
    CLASS CORE ;
    FOREIGN XOR4S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.880 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.460 2.810 9.750 3.210 ;
        RECT  9.470 0.620 9.750 3.300 ;
        RECT  9.440 0.910 9.750 1.310 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.450 2.740 ;
        RECT  0.120 2.280 0.580 2.740 ;
        RECT  0.120 3.910 2.910 4.150 ;
        RECT  3.920 3.910 4.320 4.320 ;
        RECT  2.670 4.080 4.320 4.320 ;
        RECT  0.120 2.280 0.360 4.150 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.940 1.690 2.740 ;
        RECT  1.300 1.940 1.690 2.340 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 2.130 14.760 2.740 ;
        RECT  14.300 2.280 14.760 2.740 ;
        RECT  14.520 2.130 14.760 4.240 ;
        RECT  11.850 4.000 14.760 4.240 ;
        RECT  11.850 4.000 12.090 4.420 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.190 1.940 13.580 2.340 ;
        RECT  13.190 1.940 13.470 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 0.560 ;
        RECT  7.840 -0.380 8.800 0.560 ;
        RECT  12.370 -0.380 12.770 0.560 ;
        RECT  14.030 -0.380 14.430 0.560 ;
        RECT  0.000 -0.380 14.880 0.380 ;
        RECT  0.440 -0.380 0.840 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 4.480 2.060 5.420 ;
        RECT  7.280 4.200 7.680 5.420 ;
        RECT  8.820 4.150 9.220 5.420 ;
        RECT  12.480 4.480 12.880 5.420 ;
        RECT  13.790 4.480 14.190 5.420 ;
        RECT  0.000 4.660 14.880 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.820 3.130 14.280 3.530 ;
        RECT  13.820 1.760 14.060 3.530 ;
        RECT  13.890 0.800 14.130 2.000 ;
        RECT  13.890 1.200 14.360 1.600 ;
        RECT  11.460 0.800 14.130 1.040 ;
        RECT  11.460 0.620 11.860 1.040 ;
        RECT  10.490 3.430 12.950 3.670 ;
        RECT  12.710 1.280 12.950 3.670 ;
        RECT  10.490 1.200 10.730 3.670 ;
        RECT  13.320 2.980 13.560 3.380 ;
        RECT  12.710 3.060 13.560 3.300 ;
        RECT  10.480 2.670 10.730 3.070 ;
        RECT  12.310 1.760 12.950 2.160 ;
        RECT  12.710 1.280 13.650 1.520 ;
        RECT  11.920 2.380 12.160 3.070 ;
        RECT  11.830 1.280 12.070 2.620 ;
        RECT  11.830 1.280 12.250 1.520 ;
        RECT  8.720 3.660 10.230 3.900 ;
        RECT  9.990 0.640 10.230 3.900 ;
        RECT  8.720 2.420 8.960 3.900 ;
        RECT  10.970 2.750 11.520 2.990 ;
        RECT  8.300 2.420 8.960 2.820 ;
        RECT  10.970 0.640 11.210 2.990 ;
        RECT  10.970 1.280 11.530 1.520 ;
        RECT  9.990 0.640 11.210 0.880 ;
        RECT  5.960 2.740 6.360 2.980 ;
        RECT  6.040 0.740 6.280 2.980 ;
        RECT  8.790 0.800 9.030 2.050 ;
        RECT  7.320 0.800 9.030 1.040 ;
        RECT  6.040 0.740 7.560 0.980 ;
        RECT  5.730 3.700 8.040 3.940 ;
        RECT  7.800 1.280 8.040 3.940 ;
        RECT  7.800 3.300 8.470 3.540 ;
        RECT  7.800 1.280 8.460 1.520 ;
        RECT  5.320 0.620 5.560 3.480 ;
        RECT  5.320 3.220 7.560 3.460 ;
        RECT  7.320 1.870 7.560 3.460 ;
        RECT  3.340 2.630 3.920 2.870 ;
        RECT  3.680 0.620 3.920 2.870 ;
        RECT  7.230 1.870 7.560 2.270 ;
        RECT  3.350 1.180 3.920 1.420 ;
        RECT  3.680 0.620 5.560 0.860 ;
        RECT  6.680 2.740 7.080 2.980 ;
        RECT  6.750 1.220 6.990 2.980 ;
        RECT  6.680 1.220 7.080 1.460 ;
        RECT  4.780 4.180 6.850 4.420 ;
        RECT  4.780 1.100 5.020 4.420 ;
        RECT  1.930 3.430 4.480 3.670 ;
        RECT  4.240 1.100 4.480 3.670 ;
        RECT  1.930 1.280 2.170 3.670 ;
        RECT  1.320 2.980 1.560 3.380 ;
        RECT  1.320 2.980 2.170 3.220 ;
        RECT  4.240 2.550 4.520 2.950 ;
        RECT  1.930 1.850 2.570 2.250 ;
        RECT  1.320 1.280 2.170 1.520 ;
        RECT  0.600 2.980 1.060 3.380 ;
        RECT  0.820 0.800 1.060 3.380 ;
        RECT  0.680 1.200 1.060 1.600 ;
        RECT  0.820 0.800 2.980 1.040 ;
        RECT  2.740 0.620 3.440 0.860 ;
        RECT  2.560 2.790 3.050 3.190 ;
        RECT  2.810 1.280 3.050 3.190 ;
        RECT  2.560 1.280 3.050 1.520 ;
    END
END XOR4S

MACRO XOR4T
    CLASS CORE ;
    FOREIGN XOR4T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.120 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.330 2.820 10.940 3.060 ;
        RECT  9.320 1.330 10.950 1.570 ;
        RECT  10.700 2.740 10.940 3.140 ;
        RECT  10.710 1.250 10.950 1.650 ;
        RECT  10.090 1.330 10.370 3.060 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.740 0.450 2.740 ;
        RECT  0.120 2.280 0.580 2.740 ;
        RECT  0.120 3.910 2.910 4.150 ;
        RECT  4.010 3.910 4.410 4.320 ;
        RECT  2.670 4.080 4.410 4.320 ;
        RECT  0.120 2.280 0.360 4.150 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.940 1.690 2.740 ;
        RECT  1.300 1.940 1.690 2.340 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.670 2.080 16.000 2.740 ;
        RECT  15.540 2.280 16.000 2.740 ;
        RECT  15.760 2.080 16.000 4.240 ;
        RECT  13.090 4.000 16.000 4.240 ;
        RECT  13.090 4.000 13.330 4.420 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.430 1.940 14.820 2.340 ;
        RECT  14.430 1.940 14.710 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.900 -0.380 2.300 0.560 ;
        RECT  7.840 -0.380 8.800 0.560 ;
        RECT  9.970 -0.380 10.370 0.780 ;
        RECT  13.610 -0.380 14.010 0.560 ;
        RECT  15.270 -0.380 15.670 0.560 ;
        RECT  0.000 -0.380 16.120 0.380 ;
        RECT  0.440 -0.380 0.840 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 4.480 2.060 5.420 ;
        RECT  7.280 4.200 7.680 5.420 ;
        RECT  8.710 4.150 9.110 5.420 ;
        RECT  9.980 4.150 10.380 5.420 ;
        RECT  13.720 4.480 14.120 5.420 ;
        RECT  15.030 4.480 15.430 5.420 ;
        RECT  0.000 4.660 16.120 5.420 ;
        RECT  0.440 4.480 0.840 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  15.060 3.110 15.520 3.510 ;
        RECT  15.060 1.760 15.300 3.510 ;
        RECT  15.130 0.800 15.370 2.000 ;
        RECT  15.130 1.200 15.600 1.600 ;
        RECT  12.700 0.800 15.370 1.040 ;
        RECT  12.700 0.620 13.100 1.040 ;
        RECT  11.730 3.430 14.190 3.670 ;
        RECT  13.950 1.280 14.190 3.670 ;
        RECT  11.730 1.200 11.970 3.670 ;
        RECT  14.560 2.980 14.800 3.380 ;
        RECT  13.950 3.060 14.800 3.300 ;
        RECT  11.720 2.670 11.970 3.070 ;
        RECT  13.550 1.760 14.190 2.160 ;
        RECT  13.950 1.280 14.890 1.520 ;
        RECT  13.160 2.380 13.400 3.070 ;
        RECT  13.070 1.280 13.310 2.620 ;
        RECT  13.070 1.280 13.490 1.520 ;
        RECT  8.720 3.660 11.430 3.900 ;
        RECT  11.190 0.620 11.430 3.900 ;
        RECT  8.720 2.610 8.960 3.900 ;
        RECT  8.290 2.610 8.960 3.010 ;
        RECT  12.210 2.750 12.760 2.990 ;
        RECT  12.210 0.620 12.450 2.990 ;
        RECT  12.210 1.280 12.770 1.520 ;
        RECT  11.190 0.620 12.450 0.860 ;
        RECT  5.960 2.740 6.360 2.980 ;
        RECT  6.040 0.740 6.280 2.980 ;
        RECT  8.790 0.800 9.030 2.330 ;
        RECT  7.320 0.800 9.030 1.040 ;
        RECT  6.040 0.740 7.560 0.980 ;
        RECT  5.730 3.700 8.040 3.940 ;
        RECT  7.800 1.280 8.040 3.940 ;
        RECT  7.800 3.300 8.470 3.540 ;
        RECT  7.800 1.280 8.460 1.520 ;
        RECT  5.320 3.220 7.560 3.460 ;
        RECT  7.320 1.870 7.560 3.460 ;
        RECT  5.320 0.620 5.560 3.460 ;
        RECT  3.340 2.630 3.920 2.870 ;
        RECT  3.680 0.620 3.920 2.870 ;
        RECT  7.230 1.870 7.560 2.270 ;
        RECT  3.350 1.180 3.920 1.420 ;
        RECT  3.680 0.620 5.560 0.860 ;
        RECT  6.680 2.740 7.080 2.980 ;
        RECT  6.750 1.220 6.990 2.980 ;
        RECT  6.680 1.220 7.080 1.460 ;
        RECT  4.780 4.180 6.850 4.420 ;
        RECT  4.780 1.100 5.020 4.420 ;
        RECT  1.930 3.430 4.480 3.670 ;
        RECT  4.240 1.100 4.480 3.670 ;
        RECT  1.930 1.280 2.170 3.670 ;
        RECT  1.320 2.980 1.560 3.380 ;
        RECT  1.320 2.980 2.170 3.220 ;
        RECT  4.240 2.550 4.520 2.950 ;
        RECT  1.930 1.850 2.570 2.250 ;
        RECT  1.320 1.280 2.170 1.520 ;
        RECT  0.600 2.980 1.060 3.380 ;
        RECT  0.820 0.800 1.060 3.380 ;
        RECT  0.680 1.200 1.060 1.600 ;
        RECT  0.820 0.800 2.980 1.040 ;
        RECT  2.740 0.620 3.440 0.860 ;
        RECT  2.560 2.790 3.050 3.190 ;
        RECT  2.810 1.280 3.050 3.190 ;
        RECT  2.560 1.280 3.050 1.520 ;
    END
END XOR4T

END LIBRARY
