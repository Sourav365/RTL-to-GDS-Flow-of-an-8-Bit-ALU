VERSION 5.5 ;
NAMESCASESENSITIVE ON ;





LAYER metal1  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal1

LAYER metal2
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal2

LAYER metal3
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal3

LAYER metal4  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal4

LAYER metal5  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal5

LAYER metal6
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal6


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:03 CST 2007
#
#**********************************************************************




MACRO AN2
  PIN I1
   AntennaPartialMetalArea                    0.201400 LAYER metal1 ;
   AntennaGateArea                            0.167400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.274794 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.615836 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.092700 LAYER metal1 ;
  END O

END AN2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:06 CST 2007
#
#**********************************************************************




MACRO AN2B1
  PIN B1
   AntennaPartialMetalArea                    1.552000 LAYER metal1 ;
   AntennaGateArea                            0.774000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.256852 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.207200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.082262 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.058400 LAYER metal1 ;
   AntennaDiffArea                            1.722000 LAYER metal1 ;
  END O

END AN2B1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:11 CST 2007
#
#**********************************************************************




MACRO AN2B1P
  PIN B1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.972227 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.361110 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.931200 LAYER metal1 ;
   AntennaDiffArea                            2.119600 LAYER metal1 ;
  END O

END AN2B1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:14 CST 2007
#
#**********************************************************************




MACRO AN2B1S
  PIN B1
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.208584 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.207200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.858589 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.911600 LAYER metal1 ;
   AntennaDiffArea                            1.192000 LAYER metal1 ;
  END O

END AN2B1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:17 CST 2007
#
#**********************************************************************




MACRO AN2B1T
  PIN B1
   AntennaPartialMetalArea                    0.286000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.381314 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.307200 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.069692 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    2.904400 LAYER metal1 ;
   AntennaDiffArea                            2.865400 LAYER metal1 ;
  END O

END AN2B1T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:20 CST 2007
#
#**********************************************************************




MACRO AN2P
  PIN I1
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.534185 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.199200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.111107 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.697600 LAYER metal1 ;
   AntennaDiffArea                            1.846700 LAYER metal1 ;
  END O

END AN2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:22 CST 2007
#
#**********************************************************************




MACRO AN2S
  PIN I1
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.144206 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.212800 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.569737 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.612000 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END AN2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:25 CST 2007
#
#**********************************************************************




MACRO AN2T
  PIN I1
   AntennaPartialMetalArea                    0.244800 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.261618 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.303600 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.061613 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    2.816400 LAYER metal1 ;
   AntennaDiffArea                            2.899000 LAYER metal1 ;
  END O

END AN2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:27 CST 2007
#
#**********************************************************************




MACRO AN3
  PIN I1
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.718673 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.250588 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.250588 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END O

END AN3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:30 CST 2007
#
#**********************************************************************




MACRO AN3B1
  PIN B1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.642677 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.569738 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.621748 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END O

END AN3B1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:33 CST 2007
#
#**********************************************************************




MACRO AN3B1P
  PIN B1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.699497 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.484638 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.484638 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.641600 LAYER metal1 ;
   AntennaDiffArea                            1.677500 LAYER metal1 ;
  END O

END AN3B1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:35 CST 2007
#
#**********************************************************************




MACRO AN3B1S
  PIN B1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.290407 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.438127 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.460857 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.766000 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END AN3B1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:38 CST 2007
#
#**********************************************************************




MACRO AN3B1T
  PIN B1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.790407 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.637036 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.267600 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.637039 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.232400 LAYER metal1 ;
   AntennaDiffArea                            2.739000 LAYER metal1 ;
  END O

END AN3B1T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:41 CST 2007
#
#**********************************************************************




MACRO AN3B2
  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.449497 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.654037 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.350400 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.718678 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.316500 LAYER metal1 ;
  END O

END AN3B2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:44 CST 2007
#
#**********************************************************************




MACRO AN3B2P
  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.255047 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.654037 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.252800 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.718680 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.329000 LAYER metal1 ;
  END O

END AN3B2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:47 CST 2007
#
#**********************************************************************




MACRO AN3B2S
  PIN B1
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.419400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.015263 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.419400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.041013 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.207200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.918802 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.092400 LAYER metal1 ;
   AntennaDiffArea                            1.411700 LAYER metal1 ;
  END O

END AN3B2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:50 CST 2007
#
#**********************************************************************




MACRO AN3B2T
  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.255047 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.239200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.654039 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.252800 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.943704 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.122400 LAYER metal1 ;
   AntennaDiffArea                            2.664500 LAYER metal1 ;
  END O

END AN3B2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:52 CST 2007
#
#**********************************************************************




MACRO AN3P
  PIN I1
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.718673 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.302598 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.199200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.303785 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.697600 LAYER metal1 ;
   AntennaDiffArea                            1.721500 LAYER metal1 ;
  END O

END AN3P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:55 CST 2007
#
#**********************************************************************




MACRO AN3S
  PIN I1
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.984852 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.540407 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.540407 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.928400 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END AN3S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:58 CST 2007
#
#**********************************************************************




MACRO AN3T
  PIN I1
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.271800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.937458 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.271800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.678442 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.271800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.646065 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.218400 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END O

END AN3T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:02 CST 2007
#
#**********************************************************************




MACRO AN4
  PIN I1
   AntennaPartialMetalArea                    0.235600 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.325556 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.255200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.211671 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.267778 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.255600 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.267780 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.846400 LAYER metal1 ;
   AntennaDiffArea                            1.657800 LAYER metal1 ;
  END O

END AN4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:04 CST 2007
#
#**********************************************************************




MACRO AN4B1
  PIN B1
   AntennaPartialMetalArea                    1.427600 LAYER metal1 ;
   AntennaGateArea                            0.879600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.070460 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.439800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.947702 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.298400 LAYER metal1 ;
   AntennaGateArea                            0.438600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.010483 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.438600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.301418 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.732400 LAYER metal1 ;
   AntennaDiffArea                            1.927000 LAYER metal1 ;
  END O

END AN4B1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:07 CST 2007
#
#**********************************************************************




MACRO AN4B1P
  PIN B1
   AntennaPartialMetalArea                    1.127200 LAYER metal1 ;
   AntennaGateArea                            1.749600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.087598 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.215200 LAYER metal1 ;
   AntennaGateArea                            0.542400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.707595 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.249200 LAYER metal1 ;
   AntennaGateArea                            0.537600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.664808 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.547200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.998905 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    2.469600 LAYER metal1 ;
   AntennaDiffArea                            3.692400 LAYER metal1 ;
  END O

END AN4B1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:10 CST 2007
#
#**********************************************************************




MACRO AN4B1S
  PIN B1
   AntennaPartialMetalArea                    0.221600 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.859647 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.119952 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.228000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.483586 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.758842 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.372800 LAYER metal1 ;
   AntennaDiffArea                            1.211000 LAYER metal1 ;
  END O

END AN4B1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:13 CST 2007
#
#**********************************************************************




MACRO AN4B1T
  PIN B1
   AntennaPartialMetalArea                    2.572000 LAYER metal1 ;
   AntennaGateArea                            2.649600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.078347 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.527400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.660601 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.223200 LAYER metal1 ;
   AntennaGateArea                            0.527400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.660602 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.527400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.660596 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    3.200000 LAYER metal1 ;
   AntennaDiffArea                            5.811600 LAYER metal1 ;
  END O

END AN4B1T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:16 CST 2007
#
#**********************************************************************




MACRO AN4P
  PIN I1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.513600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.873052 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.504000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.814679 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.750199 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.223200 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785367 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    2.971600 LAYER metal1 ;
   AntennaDiffArea                            3.747950 LAYER metal1 ;
  END O

END AN4P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:18 CST 2007
#
#**********************************************************************




MACRO AN4S
  PIN I1
   AntennaPartialMetalArea                    0.199200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.450754 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.237200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.108585 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.040403 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.202400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.753792 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    1.102800 LAYER metal1 ;
   AntennaDiffArea                            0.956000 LAYER metal1 ;
  END O

END AN4S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:21 CST 2007
#
#**********************************************************************




MACRO AN4T
  PIN I1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.513600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.873052 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.504000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.814679 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.750199 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.223200 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785367 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    3.324800 LAYER metal1 ;
   AntennaDiffArea                            5.811600 LAYER metal1 ;
  END O

END AN4T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:24 CST 2007
#
#**********************************************************************




MACRO ANTENNA
  PIN A
   AntennaPartialMetalArea                    0.396000 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
  END A

END ANTENNA


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:27 CST 2007
#
#**********************************************************************




MACRO AO112
  PIN A1
   AntennaPartialMetalArea                    0.198000 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.667823 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.202400 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.591432 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.202000 LAYER metal1 ;
   AntennaGateArea                            0.385200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.286087 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.385200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.303218 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.553200 LAYER metal1 ;
   AntennaDiffArea                            1.363750 LAYER metal1 ;
  END O

END AO112


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:29 CST 2007
#
#**********************************************************************




MACRO AO112P
  PIN A1
   AntennaPartialMetalArea                    0.276400 LAYER metal1 ;
   AntennaGateArea                            0.437400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.017834 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.304400 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.608469 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.263200 LAYER metal1 ;
   AntennaGateArea                            0.473400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.735952 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.295200 LAYER metal1 ;
   AntennaGateArea                            0.473400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758766 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.902000 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END O

END AO112P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:32 CST 2007
#
#**********************************************************************




MACRO AO112S
  PIN A1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.774462 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.186000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.847426 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.362359 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.481759 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.853600 LAYER metal1 ;
   AntennaDiffArea                            0.661000 LAYER metal1 ;
  END O

END AO112S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:35 CST 2007
#
#**********************************************************************




MACRO AO112T
  PIN A1
   AntennaPartialMetalArea                    0.276400 LAYER metal1 ;
   AntennaGateArea                            0.437400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.017834 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.307200 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.526982 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.291200 LAYER metal1 ;
   AntennaGateArea                            0.473400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.735955 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.267200 LAYER metal1 ;
   AntennaGateArea                            0.473400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.791722 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.252400 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END O

END AO112T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:38 CST 2007
#
#**********************************************************************




MACRO AO12
  PIN A1
   AntennaPartialMetalArea                    0.225200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.377285 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.261200 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.065923 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.245600 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.505930 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.799600 LAYER metal1 ;
   AntennaDiffArea                            1.556300 LAYER metal1 ;
  END O

END AO12


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:41 CST 2007
#
#**********************************************************************




MACRO AO12P
  PIN A1
   AntennaPartialMetalArea                    0.225200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.503088 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.261200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.299444 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.629448 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.682800 LAYER metal1 ;
   AntennaDiffArea                            1.672400 LAYER metal1 ;
  END O

END AO12P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:44 CST 2007
#
#**********************************************************************




MACRO AO12S
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.095959 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.223600 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.358587 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.209200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.780804 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.852800 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END AO12S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:47 CST 2007
#
#**********************************************************************




MACRO AO12T
  PIN A1
   AntennaPartialMetalArea                    0.225200 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.683941 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.261200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.680866 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.251200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.790206 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.293200 LAYER metal1 ;
   AntennaDiffArea                            2.973700 LAYER metal1 ;
  END O

END AO12T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:49 CST 2007
#
#**********************************************************************




MACRO AO13
  PIN A1
   AntennaPartialMetalArea                    0.190400 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.795054 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.197200 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052530 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052525 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.252000 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.374746 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.718400 LAYER metal1 ;
   AntennaDiffArea                            1.636950 LAYER metal1 ;
  END O

END AO13


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:52 CST 2007
#
#**********************************************************************




MACRO AO13P
  PIN A1
   AntennaPartialMetalArea                    0.225200 LAYER metal1 ;
   AntennaGateArea                            0.455400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.021520 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.234600 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.618390 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.618389 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.252000 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.790206 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.900800 LAYER metal1 ;
   AntennaDiffArea                            1.739600 LAYER metal1 ;
  END O

END AO13P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:55 CST 2007
#
#**********************************************************************




MACRO AO13S
  PIN A1
   AntennaPartialMetalArea                    0.185600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.233583 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.209200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.830129 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.202400 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.736113 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.186000 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.300210 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.960400 LAYER metal1 ;
   AntennaDiffArea                            0.614200 LAYER metal1 ;
  END O

END AO13S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:57 CST 2007
#
#**********************************************************************




MACRO AO13T
  PIN A1
   AntennaPartialMetalArea                    0.281200 LAYER metal1 ;
   AntennaGateArea                            0.455400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.021521 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.302600 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.618384 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.249200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.618385 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.279000 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.790202 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    1.198400 LAYER metal1 ;
   AntennaDiffArea                            3.063950 LAYER metal1 ;
  END O

END AO13T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:00 CST 2007
#
#**********************************************************************




MACRO AO22
  PIN A1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.327000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.533335 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.190000 LAYER metal1 ;
   AntennaGateArea                            0.327000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.555350 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.322200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.533833 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.209600 LAYER metal1 ;
   AntennaGateArea                            0.322200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.902542 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.500000 LAYER metal1 ;
   AntennaDiffArea                            1.280450 LAYER metal1 ;
  END O

END AO22


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:03 CST 2007
#
#**********************************************************************




MACRO AO222
  PIN A1
   AntennaPartialMetalArea                    0.251600 LAYER metal1 ;
   AntennaGateArea                            0.384600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.188244 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.384600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.149251 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.272000 LAYER metal1 ;
   AntennaGateArea                            0.386400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.178056 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.382800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.281083 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.214000 LAYER metal1 ;
   AntennaGateArea                            0.390000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.437952 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.240000 LAYER metal1 ;
   AntennaGateArea                            0.390000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.133335 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.550400 LAYER metal1 ;
   AntennaDiffArea                            1.254950 LAYER metal1 ;
  END O

END AO222


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:06 CST 2007
#
#**********************************************************************




MACRO AO222P
  PIN A1
   AntennaPartialMetalArea                    0.199600 LAYER metal1 ;
   AntennaGateArea                            0.463800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.914192 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.455400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.022619 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.212000 LAYER metal1 ;
   AntennaGateArea                            0.459600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.981289 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.453600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.934741 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.214000 LAYER metal1 ;
   AntennaGateArea                            0.458400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.184119 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.244000 LAYER metal1 ;
   AntennaGateArea                            0.458400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.924954 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.854000 LAYER metal1 ;
   AntennaDiffArea                            1.606500 LAYER metal1 ;
  END O

END AO222P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:09 CST 2007
#
#**********************************************************************




MACRO AO222S
  PIN A1
   AntennaPartialMetalArea                    0.191600 LAYER metal1 ;
   AntennaGateArea                            0.309000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.680905 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.765584 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.307200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.690759 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.759483 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.214000 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.161928 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.240000 LAYER metal1 ;
   AntennaGateArea                            0.304800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.704068 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.796800 LAYER metal1 ;
   AntennaDiffArea                            0.603000 LAYER metal1 ;
  END O

END AO222S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:12 CST 2007
#
#**********************************************************************




MACRO AO222T
  PIN A1
   AntennaPartialMetalArea                    0.227600 LAYER metal1 ;
   AntennaGateArea                            0.517800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.730008 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.248400 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.789167 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.248400 LAYER metal1 ;
   AntennaGateArea                            0.519000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.764937 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.516600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.716226 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.214000 LAYER metal1 ;
   AntennaGateArea                            0.517800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.943993 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.280400 LAYER metal1 ;
   AntennaGateArea                            0.517800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.714558 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.246000 LAYER metal1 ;
   AntennaDiffArea                            2.747450 LAYER metal1 ;
  END O

END AO222T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:15 CST 2007
#
#**********************************************************************




MACRO AO22P
  PIN A1
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.489000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.797140 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.177600 LAYER metal1 ;
   AntennaGateArea                            0.489000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.833130 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.494400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784791 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.206400 LAYER metal1 ;
   AntennaGateArea                            0.494400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.042884 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.640000 LAYER metal1 ;
   AntennaDiffArea                            1.799850 LAYER metal1 ;
  END O

END AO22P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:19 CST 2007
#
#**********************************************************************




MACRO AO22S
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.198178 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.204400 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.198180 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.522388 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.923713 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.799600 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END AO22S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:21 CST 2007
#
#**********************************************************************




MACRO AO22T
  PIN A1
   AntennaPartialMetalArea                    0.233600 LAYER metal1 ;
   AntennaGateArea                            0.561000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.624241 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.193600 LAYER metal1 ;
   AntennaGateArea                            0.561000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.655612 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.567600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.613812 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.224400 LAYER metal1 ;
   AntennaGateArea                            0.566400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.832624 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.205600 LAYER metal1 ;
   AntennaDiffArea                            2.998400 LAYER metal1 ;
  END O

END AO22T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:24 CST 2007
#
#**********************************************************************




MACRO AOI112H
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.528200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.770318 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.528200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.770318 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            1.690200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.696485 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.690200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.696486 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    2.613200 LAYER metal1 ;
   AntennaDiffArea                            4.809500 LAYER metal1 ;
  END O

END AOI112H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:28 CST 2007
#
#**********************************************************************




MACRO AOI112HP
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.056400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.848057 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.056400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.848057 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    4.492000 LAYER metal1 ;
   AntennaDiffArea                            8.310600 LAYER metal1 ;
  END O

END AOI112HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:31 CST 2007
#
#**********************************************************************




MACRO AOI112HS
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.018800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.692580 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            1.018800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.692579 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.666800 LAYER metal1 ;
   AntennaDiffArea                            2.770200 LAYER metal1 ;
  END O

END AOI112HS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:34 CST 2007
#
#**********************************************************************




MACRO AOI112HT
  PIN A1
   AntennaPartialMetalArea                    0.207200 LAYER metal1 ;
   AntennaGateArea                            4.584600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.873969 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.207200 LAYER metal1 ;
   AntennaGateArea                            4.584600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.873969 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            5.070600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.790202 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            5.070600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.790202 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    6.959600 LAYER metal1 ;
   AntennaDiffArea                           13.140900 LAYER metal1 ;
  END O

END AOI112HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:37 CST 2007
#
#**********************************************************************




MACRO AOI12H
  PIN A1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            1.072800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.678225 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    2.042800 LAYER metal1 ;
   AntennaDiffArea                            3.630200 LAYER metal1 ;
  END O

END AOI12H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:40 CST 2007
#
#**********************************************************************




MACRO AOI12HP
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.145600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.815622 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    3.354400 LAYER metal1 ;
   AntennaDiffArea                            5.960600 LAYER metal1 ;
  END O

END AOI12HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:42 CST 2007
#
#**********************************************************************




MACRO AOI12HS
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.536400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.649515 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.618388 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.223600 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.821444 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.239200 LAYER metal1 ;
   AntennaDiffArea                            2.328000 LAYER metal1 ;
  END O

END AOI12HS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:46 CST 2007
#
#**********************************************************************




MACRO AOI12HT
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.218400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.840915 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    4.453600 LAYER metal1 ;
   AntennaDiffArea                            8.308400 LAYER metal1 ;
  END O

END AOI12HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:49 CST 2007
#
#**********************************************************************




MACRO AOI13H
  PIN A1
   AntennaPartialMetalArea                    0.234000 LAYER metal1 ;
   AntennaGateArea                            1.018800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.692579 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.261800 LAYER metal1 ;
   AntennaGateArea                            1.067400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.718756 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.223600 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.252000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    1.562400 LAYER metal1 ;
   AntennaDiffArea                            2.739200 LAYER metal1 ;
  END O

END AOI13H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:53 CST 2007
#
#**********************************************************************




MACRO AOI13HP
  PIN A1
   AntennaPartialMetalArea                    0.234000 LAYER metal1 ;
   AntennaGateArea                            2.001600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.823741 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.261800 LAYER metal1 ;
   AntennaGateArea                            2.194200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.751435 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.223600 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.252000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    2.517600 LAYER metal1 ;
   AntennaDiffArea                            4.904900 LAYER metal1 ;
  END O

END AOI13HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:56 CST 2007
#
#**********************************************************************




MACRO AOI13HS
  PIN A1
   AntennaPartialMetalArea                    0.331600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.683938 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.363800 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.712108 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.347600 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.618392 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.252000 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.889693 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    1.564800 LAYER metal1 ;
   AntennaDiffArea                            1.840700 LAYER metal1 ;
  END O

END AOI13HS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:59 CST 2007
#
#**********************************************************************




MACRO AOI13HT
  PIN A1
   AntennaPartialMetalArea                    0.234000 LAYER metal1 ;
   AntennaGateArea                            2.957400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.876445 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.255000 LAYER metal1 ;
   AntennaGateArea                            3.317400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.781335 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.210000 LAYER metal1 ;
   AntennaGateArea                            3.285000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.789041 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.240000 LAYER metal1 ;
   AntennaGateArea                            3.285000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.789041 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    3.508800 LAYER metal1 ;
   AntennaDiffArea                            6.996900 LAYER metal1 ;
  END O

END AOI13HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:02 CST 2007
#
#**********************************************************************




MACRO AOI222H
  PIN A1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            1.690200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.696485 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            1.690200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.696485 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.690200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.696486 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.690200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.696486 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.690200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.696486 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.690200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.696486 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    4.006400 LAYER metal1 ;
   AntennaDiffArea                            6.901800 LAYER metal1 ;
  END O

END AOI222H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:07 CST 2007
#
#**********************************************************************




MACRO AOI222HP
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.181600 LAYER metal1 ;
   AntennaGateArea                            3.292200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.788105 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    6.612800 LAYER metal1 ;
   AntennaDiffArea                           12.188400 LAYER metal1 ;
  END O

END AOI222HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:10 CST 2007
#
#**********************************************************************




MACRO AOI222HS
  PIN A1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.235200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    2.861600 LAYER metal1 ;
   AntennaDiffArea                            4.082400 LAYER metal1 ;
  END O

END AOI222HS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:13 CST 2007
#
#**********************************************************************




MACRO AOI22H
  PIN A1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            1.103400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.639478 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.575200 LAYER metal1 ;
   AntennaDiffArea                            3.364800 LAYER metal1 ;
  END O

END AOI22H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:17 CST 2007
#
#**********************************************************************




MACRO AOI22HP
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.165400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.761430 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    2.842400 LAYER metal1 ;
   AntennaDiffArea                            6.741600 LAYER metal1 ;
  END O

END AOI22HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:19 CST 2007
#
#**********************************************************************




MACRO AOI22HT
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    4.330400 LAYER metal1 ;
   AntennaDiffArea                           10.141200 LAYER metal1 ;
  END O

END AOI22HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:22 CST 2007
#
#**********************************************************************




MACRO AOI22S
  PIN A1
   AntennaPartialMetalArea                    0.197600 LAYER metal1 ;
   AntennaGateArea                            0.562200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.752404 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.186800 LAYER metal1 ;
   AntennaGateArea                            0.565200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.699218 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.289200 LAYER metal1 ;
   AntennaGateArea                            0.541800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.821334 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.571800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.710039 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.830400 LAYER metal1 ;
   AntennaDiffArea                            1.368000 LAYER metal1 ;
  END O

END AOI22S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:25 CST 2007
#
#**********************************************************************




MACRO BHD1
  PIN H
   AntennaPartialMetalArea                    1.425300 LAYER metal1 ;
   AntennaGateArea                            0.349200 LAYER metal1 ;
   AntennaDiffArea                            0.492800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.243415 LAYER metal1 ; 
  END H

END BHD1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:28 CST 2007
#
#**********************************************************************




MACRO BUF1
  PIN I
   AntennaPartialMetalArea                    0.199200 LAYER metal1 ;
   AntennaGateArea                            0.196200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.941899 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.586800 LAYER metal1 ;
   AntennaDiffArea                            1.538600 LAYER metal1 ;
  END O

END BUF1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:31 CST 2007
#
#**********************************************************************




MACRO BUF12CK
  PIN I
   AntennaPartialMetalArea                    0.277200 LAYER metal1 ;
   AntennaGateArea                            2.257200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.944973 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                   16.699200 LAYER metal1 ;
   AntennaDiffArea                            9.072000 LAYER metal1 ;
  END O

END BUF12CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:34 CST 2007
#
#**********************************************************************




MACRO BUF1CK
  PIN I
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.313200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.553639 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.152000 LAYER metal1 ;
   AntennaDiffArea                            1.288700 LAYER metal1 ;
  END O

END BUF1CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:36 CST 2007
#
#**********************************************************************




MACRO BUF1S
  PIN I
   AntennaPartialMetalArea                    0.334000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.477274 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.844000 LAYER metal1 ;
   AntennaDiffArea                            0.568400 LAYER metal1 ;
  END O

END BUF1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:39 CST 2007
#
#**********************************************************************




MACRO BUF2
  PIN I
   AntennaPartialMetalArea                    0.222400 LAYER metal1 ;
   AntennaGateArea                            0.369000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.217340 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.948600 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END O

END BUF2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:42 CST 2007
#
#**********************************************************************




MACRO BUF2CK
  PIN I
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.361800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.251519 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.066800 LAYER metal1 ;
   AntennaDiffArea                            1.420200 LAYER metal1 ;
  END O

END BUF2CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:44 CST 2007
#
#**********************************************************************




MACRO BUF3
  PIN I
   AntennaPartialMetalArea                    0.344000 LAYER metal1 ;
   AntennaGateArea                            0.567000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.844798 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.576800 LAYER metal1 ;
   AntennaDiffArea                            2.948150 LAYER metal1 ;
  END O

END BUF3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:47 CST 2007
#
#**********************************************************************




MACRO BUF3CK
  PIN I
   AntennaPartialMetalArea                    0.193200 LAYER metal1 ;
   AntennaGateArea                            0.565200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.675164 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    3.168400 LAYER metal1 ;
   AntennaDiffArea                            2.708900 LAYER metal1 ;
  END O

END BUF3CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:50 CST 2007
#
#**********************************************************************




MACRO BUF4
  PIN I
   AntennaPartialMetalArea                    0.199600 LAYER metal1 ;
   AntennaGateArea                            0.594000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.756903 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    2.354500 LAYER metal1 ;
   AntennaDiffArea                            2.794700 LAYER metal1 ;
  END O

END BUF4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:52 CST 2007
#
#**********************************************************************




MACRO BUF4CK
  PIN I
   AntennaPartialMetalArea                    0.193200 LAYER metal1 ;
   AntennaGateArea                            0.752400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.055022 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    3.168400 LAYER metal1 ;
   AntennaDiffArea                            3.104200 LAYER metal1 ;
  END O

END BUF4CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:55 CST 2007
#
#**********************************************************************




MACRO BUF6
  PIN I
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.080000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.491484 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    6.915600 LAYER metal1 ;
   AntennaDiffArea                            5.119200 LAYER metal1 ;
  END O

END BUF6


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:37:57 CST 2007
#
#**********************************************************************




MACRO BUF6CK
  PIN I
   AntennaPartialMetalArea                    0.193200 LAYER metal1 ;
   AntennaGateArea                            1.130400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.310507 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    5.661600 LAYER metal1 ;
   AntennaDiffArea                            4.471800 LAYER metal1 ;
  END O

END BUF6CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:00 CST 2007
#
#**********************************************************************




MACRO BUF8
  PIN I
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            1.225200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.735635 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    7.238000 LAYER metal1 ;
   AntennaDiffArea                            6.613550 LAYER metal1 ;
  END O

END BUF8


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:04 CST 2007
#
#**********************************************************************




MACRO BUF8CK
  PIN I
   AntennaPartialMetalArea                    0.193200 LAYER metal1 ;
   AntennaGateArea                            1.504800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.222491 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    7.879200 LAYER metal1 ;
   AntennaDiffArea                            6.288500 LAYER metal1 ;
  END O

END BUF8CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:06 CST 2007
#
#**********************************************************************




MACRO BUFB1
  PIN EB
   AntennaPartialMetalArea                    0.840600 LAYER metal1 ;
   AntennaGateArea                            0.871800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.938478 LAYER metal1 ; 
  END EB

  PIN I
   AntennaPartialMetalArea                    0.292000 LAYER metal1 ;
   AntennaGateArea                            0.375600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.642707 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.012800 LAYER metal1 ;
   AntennaDiffArea                            1.426850 LAYER metal1 ;
  END O

END BUFB1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:09 CST 2007
#
#**********************************************************************




MACRO BUFB2
  PIN EB
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.446400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.947135 LAYER metal1 ; 
  END EB

  PIN I
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.547200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.585525 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.936000 LAYER metal1 ;
   AntennaDiffArea                            1.698500 LAYER metal1 ;
  END O

END BUFB2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:12 CST 2007
#
#**********************************************************************




MACRO BUFB3
  PIN EB
   AntennaPartialMetalArea                    0.210800 LAYER metal1 ;
   AntennaGateArea                            0.529200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.366403 LAYER metal1 ; 
  END EB

  PIN I
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.658800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.049180 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.535400 LAYER metal1 ;
   AntennaDiffArea                            2.998300 LAYER metal1 ;
  END O

END BUFB3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:14 CST 2007
#
#**********************************************************************




MACRO BUFT1
  PIN E
   AntennaPartialMetalArea                    1.188400 LAYER metal1 ;
   AntennaGateArea                            0.693000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.938477 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.292000 LAYER metal1 ;
   AntennaGateArea                            0.375600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.642707 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.012800 LAYER metal1 ;
   AntennaDiffArea                            1.425050 LAYER metal1 ;
  END O

END BUFT1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:17 CST 2007
#
#**********************************************************************




MACRO BUFT2
  PIN E
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.477000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.883649 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.549000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.086698 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.022400 LAYER metal1 ;
   AntennaDiffArea                            1.512550 LAYER metal1 ;
  END O

END BUFT2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:20 CST 2007
#
#**********************************************************************




MACRO BUFT3
  PIN E
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.511200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.804582 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.191400 LAYER metal1 ;
   AntennaGateArea                            0.673200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.460786 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.442400 LAYER metal1 ;
   AntennaDiffArea                            2.790450 LAYER metal1 ;
  END O

END BUFT3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:23 CST 2007
#
#**********************************************************************




MACRO BUFT4
  PIN E
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.619200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.498544 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.905400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.601506 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.473000 LAYER metal1 ;
   AntennaDiffArea                            2.999250 LAYER metal1 ;
  END O

END BUFT4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:28 CST 2007
#
#**********************************************************************




MACRO CMPE4
  PIN A0
   AntennaPartialMetalArea                    0.224400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.472223 LAYER metal1 ; 
  END A0

  PIN A1
   AntennaPartialMetalArea                    0.300400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.404045 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.300400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.404045 LAYER metal1 ; 
  END A2

  PIN A3
   AntennaPartialMetalArea                    0.372400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.472220 LAYER metal1 ; 
  END A3

  PIN B0
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.809347 LAYER metal1 ; 
  END B0

  PIN B1
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.896463 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.877521 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.215600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.816284 LAYER metal1 ; 
  END B3

  PIN OEQ
   AntennaPartialMetalArea                    1.596000 LAYER metal1 ;
   AntennaDiffArea                            1.794600 LAYER metal1 ;
  END OEQ

END CMPE4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:32 CST 2007
#
#**********************************************************************




MACRO CMPE4S
  PIN A0
   AntennaPartialMetalArea                    0.224400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.756313 LAYER metal1 ; 
  END A0

  PIN A1
   AntennaPartialMetalArea                    0.311600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.404038 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.404038 LAYER metal1 ; 
  END A2

  PIN A3
   AntennaPartialMetalArea                    0.246400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.938134 LAYER metal1 ; 
  END A3

  PIN B0
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          8.166667 LAYER metal1 ; 
  END B0

  PIN B1
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.697603 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.843431 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.215600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          8.215274 LAYER metal1 ; 
  END B3

  PIN OEQ
   AntennaPartialMetalArea                    1.545600 LAYER metal1 ;
   AntennaDiffArea                            1.454000 LAYER metal1 ;
  END OEQ

END CMPE4S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:37 CST 2007
#
#**********************************************************************




MACRO DBFRBN
  PIN CKB
   AntennaPartialMetalArea                    0.209600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.977278 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.778958 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.628000 LAYER metal1 ;
   AntennaDiffArea                            1.218700 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.759200 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.193997 LAYER metal1 ; 
  END RB

END DBFRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:40 CST 2007
#
#**********************************************************************




MACRO DBFRSBN
  PIN CKB
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.392680 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.604000 LAYER metal1 ;
   AntennaDiffArea                            1.218700 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.735200 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.455600 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.212616 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    1.566000 LAYER metal1 ;
   AntennaGateArea                            0.504000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.216307 LAYER metal1 ; 
  END SB

END DBFRSBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:43 CST 2007
#
#**********************************************************************




MACRO DBHRBN
  PIN CKB
   AntennaPartialMetalArea                    0.494200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.790401 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.306800 LAYER metal1 ;
   AntennaGateArea                            0.268200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.536168 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.709600 LAYER metal1 ;
   AntennaDiffArea                            1.165500 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.589600 LAYER metal1 ;
   AntennaDiffArea                            1.172500 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.323200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.230859 LAYER metal1 ; 
  END RB

END DBHRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:46 CST 2007
#
#**********************************************************************




MACRO DBHRBS
  PIN CKB
   AntennaPartialMetalArea                    0.494200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.790401 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.306800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.601011 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.709600 LAYER metal1 ;
   AntennaDiffArea                            0.784000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.589600 LAYER metal1 ;
   AntennaDiffArea                            0.784000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.323200 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.350949 LAYER metal1 ; 
  END RB

END DBHRBS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:49 CST 2007
#
#**********************************************************************




MACRO DBZRBN
  PIN CKB
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.506313 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.628000 LAYER metal1 ;
   AntennaDiffArea                            1.218700 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.759200 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.193997 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227899 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DBZRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:52 CST 2007
#
#**********************************************************************




MACRO DBZRSBN
  PIN CKB
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.506313 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.604000 LAYER metal1 ;
   AntennaDiffArea                            1.218700 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.735200 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.455600 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.212616 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    1.566000 LAYER metal1 ;
   AntennaGateArea                            0.504000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.216307 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227899 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DBZRSBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:55 CST 2007
#
#**********************************************************************




MACRO DELA
  PIN I
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.281569 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.841600 LAYER metal1 ;
   AntennaDiffArea                            1.460200 LAYER metal1 ;
  END O

END DELA


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:38:58 CST 2007
#
#**********************************************************************




MACRO DELB
  PIN I
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.281569 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.841600 LAYER metal1 ;
   AntennaDiffArea                            1.460200 LAYER metal1 ;
  END O

END DELB


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:00 CST 2007
#
#**********************************************************************




MACRO DELC
  PIN I
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.281569 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.841600 LAYER metal1 ;
   AntennaDiffArea                            1.470000 LAYER metal1 ;
  END O

END DELC


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:07 CST 2007
#
#**********************************************************************




MACRO DFCLRBN
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.443183 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.672701 LAYER metal1 ; 
  END D

  PIN LD
   AntennaPartialMetalArea                    1.648800 LAYER metal1 ;
   AntennaGateArea                            0.716400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.967172 LAYER metal1 ; 
  END LD

  PIN Q
   AntennaPartialMetalArea                    0.927600 LAYER metal1 ;
   AntennaDiffArea                            1.073800 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.654800 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.260000 LAYER metal1 ;
   AntennaGateArea                            0.487800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.776955 LAYER metal1 ; 
  END RB

END DFCLRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:09 CST 2007
#
#**********************************************************************




MACRO DFCRBN
  PIN CK
   AntennaPartialMetalArea                    0.297600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.164142 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.297600 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.688318 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.876000 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.677200 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755556 LAYER metal1 ; 
  END RB

END DFCRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:12 CST 2007
#
#**********************************************************************




MACRO DFFN
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.517678 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.285600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.890850 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.893200 LAYER metal1 ;
   AntennaDiffArea                            1.063300 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.505600 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

END DFFN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:15 CST 2007
#
#**********************************************************************




MACRO DFFP
  PIN CK
   AntennaPartialMetalArea                    0.297600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.704542 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.959957 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.878400 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    1.204000 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QB

END DFFP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:17 CST 2007
#
#**********************************************************************




MACRO DFFRBN
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.977273 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.778958 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.628000 LAYER metal1 ;
   AntennaDiffArea                            1.218700 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.759200 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.662400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.233096 LAYER metal1 ; 
  END RB

END DFFRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:20 CST 2007
#
#**********************************************************************




MACRO DFFRBP
  PIN CK
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.404040 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.770320 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.840000 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.746400 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.898200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.793361 LAYER metal1 ; 
  END RB

END DFFRBP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:23 CST 2007
#
#**********************************************************************




MACRO DFFRBS
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.977273 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.778958 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.501200 LAYER metal1 ;
   AntennaDiffArea                            0.624400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    1.014000 LAYER metal1 ;
   AntennaDiffArea                            0.769300 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.608400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.357333 LAYER metal1 ; 
  END RB

END DFFRBS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:26 CST 2007
#
#**********************************************************************




MACRO DFFRBT
  PIN CK
   AntennaPartialMetalArea                    0.249600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.472222 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    1.616000 LAYER metal1 ;
   AntennaDiffArea                            2.917300 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    2.069600 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.898200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.791361 LAYER metal1 ; 
  END RB

END DFFRBT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:29 CST 2007
#
#**********************************************************************




MACRO DFFRSBN
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.279043 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.604000 LAYER metal1 ;
   AntennaDiffArea                            1.218700 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.735200 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.455600 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.212616 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    1.558800 LAYER metal1 ;
   AntennaGateArea                            0.525600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.795597 LAYER metal1 ; 
  END SB

END DFFRSBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:32 CST 2007
#
#**********************************************************************




MACRO DFFS
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.517678 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.285600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.890850 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.893200 LAYER metal1 ;
   AntennaDiffArea                            0.626500 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.687600 LAYER metal1 ;
   AntennaDiffArea                            0.769300 LAYER metal1 ;
  END QB

END DFFS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:34 CST 2007
#
#**********************************************************************




MACRO DFFSBN
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.279043 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.684000 LAYER metal1 ;
   AntennaDiffArea                            1.061200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.500000 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN SB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.793800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.959691 LAYER metal1 ; 
  END SB

END DFFSBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:37 CST 2007
#
#**********************************************************************




MACRO DFTRBN
  PIN CK
   AntennaPartialMetalArea                    0.245600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.347225 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.778958 LAYER metal1 ; 
  END D

  PIN E
   AntennaPartialMetalArea                    0.292800 LAYER metal1 ;
   AntennaGateArea                            0.756000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.520368 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.906800 LAYER metal1 ;
   AntennaDiffArea                            1.126300 LAYER metal1 ;
  END Q

  PIN QZ
   AntennaPartialMetalArea                    0.822800 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QZ

  PIN RB
   AntennaPartialMetalArea                    0.293900 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.253759 LAYER metal1 ; 
  END RB

END DFTRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:40 CST 2007
#
#**********************************************************************




MACRO DFTRBS
  PIN CK
   AntennaPartialMetalArea                    0.245600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.347225 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.778958 LAYER metal1 ; 
  END D

  PIN E
   AntennaPartialMetalArea                    0.295600 LAYER metal1 ;
   AntennaGateArea                            0.522000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.463216 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.972000 LAYER metal1 ;
   AntennaDiffArea                            0.746200 LAYER metal1 ;
  END Q

  PIN QZ
   AntennaPartialMetalArea                    1.508000 LAYER metal1 ;
   AntennaDiffArea                            1.134400 LAYER metal1 ;
  END QZ

  PIN RB
   AntennaPartialMetalArea                    0.293900 LAYER metal1 ;
   AntennaGateArea                            0.615600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.394410 LAYER metal1 ; 
  END RB

END DFTRBS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:43 CST 2007
#
#**********************************************************************




MACRO DFZCLRBN
  PIN CK
   AntennaPartialMetalArea                    0.297600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.954542 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.238000 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.672705 LAYER metal1 ; 
  END D

  PIN LD
   AntennaPartialMetalArea                    1.508000 LAYER metal1 ;
   AntennaGateArea                            0.716400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.506311 LAYER metal1 ; 
  END LD

  PIN Q
   AntennaPartialMetalArea                    0.768000 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.666400 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.304800 LAYER metal1 ;
   AntennaGateArea                            0.487800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.776954 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    1.343200 LAYER metal1 ;
   AntennaGateArea                            0.721800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.662977 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.316800 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.703940 LAYER metal1 ; 
  END TD

END DFZCLRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:47 CST 2007
#
#**********************************************************************




MACRO DFZCRBN
  PIN CK
   AntennaPartialMetalArea                    0.233600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.688133 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.294400 LAYER metal1 ;
   AntennaGateArea                            0.561600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.701563 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.834000 LAYER metal1 ;
   AntennaDiffArea                            1.090600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.626000 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.330400 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.543858 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.435600 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.481636 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.283600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.631316 LAYER metal1 ; 
  END TD

END DFZCRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:50 CST 2007
#
#**********************************************************************




MACRO DFZN
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.517678 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.893200 LAYER metal1 ;
   AntennaDiffArea                            1.063300 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.505600 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277069 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:53 CST 2007
#
#**********************************************************************




MACRO DFZP
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.494948 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.905600 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    1.019200 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277069 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:39:57 CST 2007
#
#**********************************************************************




MACRO DFZRBN
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.506313 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.628000 LAYER metal1 ;
   AntennaDiffArea                            1.218700 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.759200 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.662400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.233096 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227899 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:00 CST 2007
#
#**********************************************************************




MACRO DFZRBP
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.494953 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.778400 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.658400 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.898200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.793368 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227899 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZRBP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:03 CST 2007
#
#**********************************************************************




MACRO DFZRBS
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.506313 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.517200 LAYER metal1 ;
   AntennaDiffArea                            0.720400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    1.014000 LAYER metal1 ;
   AntennaDiffArea                            0.769300 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.608400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.378043 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227899 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZRBS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:08 CST 2007
#
#**********************************************************************




MACRO DFZRBT
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.494948 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    1.618400 LAYER metal1 ;
   AntennaDiffArea                            2.917300 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    1.997600 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.209600 LAYER metal1 ;
   AntennaGateArea                            0.898200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.791364 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277069 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZRBT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:11 CST 2007
#
#**********************************************************************




MACRO DFZRSBN
  PIN CK
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.063133 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.517200 LAYER metal1 ;
   AntennaDiffArea                            1.061200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.990000 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.455600 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.212616 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    1.569200 LAYER metal1 ;
   AntennaGateArea                            0.525600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.795600 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.193384 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZRSBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:15 CST 2007
#
#**********************************************************************




MACRO DFZS
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.517678 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.893200 LAYER metal1 ;
   AntennaDiffArea                            0.626500 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.687600 LAYER metal1 ;
   AntennaDiffArea                            0.769300 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277069 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:18 CST 2007
#
#**********************************************************************




MACRO DFZSBN
  PIN CK
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.063133 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.660000 LAYER metal1 ;
   AntennaDiffArea                            1.061200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.500000 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN SB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.793800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.959691 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.193384 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZSBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:20 CST 2007
#
#**********************************************************************




MACRO DFZTRBN
  PIN CK
   AntennaPartialMetalArea                    0.245600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.506315 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN E
   AntennaPartialMetalArea                    0.292800 LAYER metal1 ;
   AntennaGateArea                            0.756000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.520368 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.855600 LAYER metal1 ;
   AntennaDiffArea                            1.162000 LAYER metal1 ;
  END Q

  PIN QZ
   AntennaPartialMetalArea                    0.755600 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QZ

  PIN RB
   AntennaPartialMetalArea                    0.293900 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.280779 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.243029 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZTRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:23 CST 2007
#
#**********************************************************************




MACRO DFZTRBS
  PIN CK
   AntennaPartialMetalArea                    0.245600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.506315 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN E
   AntennaPartialMetalArea                    0.295600 LAYER metal1 ;
   AntennaGateArea                            0.522000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.463216 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.972000 LAYER metal1 ;
   AntennaDiffArea                            0.746200 LAYER metal1 ;
  END Q

  PIN QZ
   AntennaPartialMetalArea                    1.508000 LAYER metal1 ;
   AntennaDiffArea                            1.134400 LAYER metal1 ;
  END QZ

  PIN RB
   AntennaPartialMetalArea                    0.293900 LAYER metal1 ;
   AntennaGateArea                            0.615600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.394410 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.243029 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END DFZTRBS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:26 CST 2007
#
#**********************************************************************




MACRO DLHN
  PIN CK
   AntennaPartialMetalArea                    0.310000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.338379 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.293600 LAYER metal1 ;
   AntennaGateArea                            0.253800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.424744 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.890400 LAYER metal1 ;
   AntennaDiffArea                            0.991200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.575600 LAYER metal1 ;
   AntennaDiffArea                            1.411200 LAYER metal1 ;
  END QB

END DLHN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:31 CST 2007
#
#**********************************************************************




MACRO DLHP
  PIN CK
   AntennaPartialMetalArea                    0.353200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.717172 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.388400 LAYER metal1 ;
   AntennaGateArea                            0.271800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.348048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.773600 LAYER metal1 ;
   AntennaDiffArea                            1.641600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.580000 LAYER metal1 ;
   AntennaDiffArea                            1.641600 LAYER metal1 ;
  END QB

END DLHP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:36 CST 2007
#
#**********************************************************************




MACRO DLHRBN
  PIN CK
   AntennaPartialMetalArea                    0.494200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.790401 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.306800 LAYER metal1 ;
   AntennaGateArea                            0.268200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.536168 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.709600 LAYER metal1 ;
   AntennaDiffArea                            1.165500 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.589600 LAYER metal1 ;
   AntennaDiffArea                            1.253000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.323200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.230859 LAYER metal1 ; 
  END RB

END DLHRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:39 CST 2007
#
#**********************************************************************




MACRO DLHRBP
  PIN CK
   AntennaPartialMetalArea                    0.494200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.790401 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.306800 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.204674 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.658800 LAYER metal1 ;
   AntennaDiffArea                            1.415600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.953200 LAYER metal1 ;
   AntennaDiffArea                            1.385650 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.323200 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.166081 LAYER metal1 ; 
  END RB

END DLHRBP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:42 CST 2007
#
#**********************************************************************




MACRO DLHRBS
  PIN CK
   AntennaPartialMetalArea                    0.494200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.790401 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.306800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.601011 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.709600 LAYER metal1 ;
   AntennaDiffArea                            0.793800 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.589600 LAYER metal1 ;
   AntennaDiffArea                            0.793800 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.323200 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.350949 LAYER metal1 ; 
  END RB

END DLHRBS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:45 CST 2007
#
#**********************************************************************




MACRO DLHS
  PIN CK
   AntennaPartialMetalArea                    0.310000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.338379 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.293600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.771465 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.851200 LAYER metal1 ;
   AntennaDiffArea                            0.632800 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.662400 LAYER metal1 ;
   AntennaDiffArea                            0.784000 LAYER metal1 ;
  END QB

END DLHS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:48 CST 2007
#
#**********************************************************************




MACRO FA1
  PIN A
   AntennaPartialMetalArea                    2.454400 LAYER metal1 ;
   AntennaGateArea                            0.554400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869952 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.726400 LAYER metal1 ;
   AntennaGateArea                            0.712800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.822840 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    4.092000 LAYER metal1 ;
   AntennaGateArea                            0.514800 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.493082 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    0.743600 LAYER metal1 ;
   AntennaDiffArea                            1.156400 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.774400 LAYER metal1 ;
   AntennaDiffArea                            1.131200 LAYER metal1 ;
  END S

END FA1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:51 CST 2007
#
#**********************************************************************




MACRO FA1P
  PIN A
   AntennaPartialMetalArea                    2.430400 LAYER metal1 ;
   AntennaGateArea                            0.554400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.858582 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.714400 LAYER metal1 ;
   AntennaGateArea                            0.712800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.844595 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    4.122000 LAYER metal1 ;
   AntennaGateArea                            0.514800 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.424207 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    1.103200 LAYER metal1 ;
   AntennaDiffArea                            1.343600 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.901600 LAYER metal1 ;
   AntennaDiffArea                            1.360350 LAYER metal1 ;
  END S

END FA1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:56 CST 2007
#
#**********************************************************************




MACRO FA1S
  PIN A
   AntennaPartialMetalArea                    4.154200 LAYER metal1 ;
   AntennaGateArea                            0.673200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.651514 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    2.636800 LAYER metal1 ;
   AntennaGateArea                            0.673200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.881315 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    2.795400 LAYER metal1 ;
   AntennaGateArea                            0.514800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.756310 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    0.491200 LAYER metal1 ;
   AntennaDiffArea                            0.623000 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.743600 LAYER metal1 ;
   AntennaDiffArea                            0.623000 LAYER metal1 ;
  END S

END FA1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:40:59 CST 2007
#
#**********************************************************************




MACRO FA1T
  PIN A
   AntennaPartialMetalArea                    2.443600 LAYER metal1 ;
   AntennaGateArea                            0.554400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.858582 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.726400 LAYER metal1 ;
   AntennaGateArea                            0.712800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.848100 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    4.282400 LAYER metal1 ;
   AntennaGateArea                            0.514800 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.424230 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    1.422400 LAYER metal1 ;
   AntennaDiffArea                            2.474550 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    1.316000 LAYER metal1 ;
   AntennaDiffArea                            2.806450 LAYER metal1 ;
  END S

END FA1T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:02 CST 2007
#
#**********************************************************************




MACRO FA2
  PIN A
   AntennaPartialMetalArea                    1.541800 LAYER metal1 ;
   AntennaGateArea                            0.568800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.840381 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    2.200800 LAYER metal1 ;
   AntennaGateArea                            0.729000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.633210 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    1.616700 LAYER metal1 ;
   AntennaGateArea                            1.486800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.257571 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    4.231200 LAYER metal1 ;
   AntennaDiffArea                            2.809300 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.774400 LAYER metal1 ;
   AntennaDiffArea                            1.108800 LAYER metal1 ;
  END S

END FA2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:04 CST 2007
#
#**********************************************************************




MACRO FA2P
  PIN A
   AntennaPartialMetalArea                    1.893600 LAYER metal1 ;
   AntennaGateArea                            0.568800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.891146 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    2.275200 LAYER metal1 ;
   AntennaGateArea                            0.729000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.593432 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    2.046600 LAYER metal1 ;
   AntennaGateArea                            2.656800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.357955 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    6.121400 LAYER metal1 ;
   AntennaDiffArea                            5.414700 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.662400 LAYER metal1 ;
   AntennaDiffArea                            1.564200 LAYER metal1 ;
  END S

END FA2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:10 CST 2007
#
#**********************************************************************




MACRO FA2S
  PIN A
   AntennaPartialMetalArea                    1.503800 LAYER metal1 ;
   AntennaGateArea                            0.568800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.789618 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    2.368800 LAYER metal1 ;
   AntennaGateArea                            0.729000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.633207 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    1.876800 LAYER metal1 ;
   AntennaGateArea                            0.802800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.156562 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    3.472000 LAYER metal1 ;
   AntennaDiffArea                            1.760200 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.774400 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END S

END FA2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:13 CST 2007
#
#**********************************************************************




MACRO FA3
  PIN A
   AntennaPartialMetalArea                    0.365600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.460859 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.437600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.354797 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    1.275800 LAYER metal1 ;
   AntennaGateArea                            1.486800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.378156 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    4.548000 LAYER metal1 ;
   AntennaDiffArea                            2.703700 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.774400 LAYER metal1 ;
   AntennaDiffArea                            1.146600 LAYER metal1 ;
  END S

END FA3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:16 CST 2007
#
#**********************************************************************




MACRO FA3P
  PIN A
   AntennaPartialMetalArea                    0.341600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.460854 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.409600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.354801 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    2.116300 LAYER metal1 ;
   AntennaGateArea                            2.656800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.595330 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    6.212500 LAYER metal1 ;
   AntennaDiffArea                            5.414700 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.662400 LAYER metal1 ;
   AntennaDiffArea                            1.564200 LAYER metal1 ;
  END S

END FA3P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:19 CST 2007
#
#**********************************************************************




MACRO FA3S
  PIN A
   AntennaPartialMetalArea                    0.384800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.460857 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.385600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.202018 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    1.870200 LAYER metal1 ;
   AntennaGateArea                            0.802800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.702024 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    3.703800 LAYER metal1 ;
   AntennaDiffArea                            1.821800 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.774400 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END S

END FA3S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:23 CST 2007
#
#**********************************************************************




MACRO FACS1
  PIN A
   AntennaPartialMetalArea                   14.433400 LAYER metal1 ;
   AntennaGateArea                            1.458000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.040449 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                   14.132800 LAYER metal1 ;
   AntennaGateArea                            1.774800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656562 LAYER metal1 ; 
  END B

  PIN CI0
   AntennaPartialMetalArea                    2.452800 LAYER metal1 ;
   AntennaGateArea                            1.342800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.662249 LAYER metal1 ; 
  END CI0

  PIN CI1
   AntennaPartialMetalArea                    2.472000 LAYER metal1 ;
   AntennaGateArea                            1.342800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656571 LAYER metal1 ; 
  END CI1

  PIN CO0
   AntennaPartialMetalArea                    2.814400 LAYER metal1 ;
   AntennaDiffArea                            2.423750 LAYER metal1 ;
  END CO0

  PIN CO1
   AntennaPartialMetalArea                    2.745600 LAYER metal1 ;
   AntennaDiffArea                            2.423450 LAYER metal1 ;
  END CO1

  PIN CS
   AntennaPartialMetalArea                    0.231200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.406562 LAYER metal1 ; 
  END CS

  PIN S
   AntennaPartialMetalArea                    0.515200 LAYER metal1 ;
   AntennaDiffArea                            1.023050 LAYER metal1 ;
  END S

END FACS1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:26 CST 2007
#
#**********************************************************************




MACRO FACS1P
  PIN A
   AntennaPartialMetalArea                   17.404000 LAYER metal1 ;
   AntennaGateArea                            1.458000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.040400 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                   17.108800 LAYER metal1 ;
   AntennaGateArea                            1.774800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656553 LAYER metal1 ; 
  END B

  PIN CI0
   AntennaPartialMetalArea                    3.315200 LAYER metal1 ;
   AntennaGateArea                            2.368800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.662243 LAYER metal1 ; 
  END CI0

  PIN CI1
   AntennaPartialMetalArea                    3.243000 LAYER metal1 ;
   AntennaGateArea                            2.368800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656562 LAYER metal1 ; 
  END CI1

  PIN CO0
   AntennaPartialMetalArea                    4.413600 LAYER metal1 ;
   AntennaDiffArea                            4.749700 LAYER metal1 ;
  END CO0

  PIN CO1
   AntennaPartialMetalArea                    4.464000 LAYER metal1 ;
   AntennaDiffArea                            4.753900 LAYER metal1 ;
  END CO1

  PIN CS
   AntennaPartialMetalArea                    0.303200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.406569 LAYER metal1 ; 
  END CS

  PIN S
   AntennaPartialMetalArea                    0.608000 LAYER metal1 ;
   AntennaDiffArea                            1.378400 LAYER metal1 ;
  END S

END FACS1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:29 CST 2007
#
#**********************************************************************




MACRO FACS1S
  PIN A
   AntennaPartialMetalArea                   13.172000 LAYER metal1 ;
   AntennaGateArea                            1.458000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.040406 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                   12.138400 LAYER metal1 ;
   AntennaGateArea                            1.774800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656594 LAYER metal1 ; 
  END B

  PIN CI0
   AntennaPartialMetalArea                    2.136000 LAYER metal1 ;
   AntennaGateArea                            0.824400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.662245 LAYER metal1 ; 
  END CI0

  PIN CI1
   AntennaPartialMetalArea                    2.290400 LAYER metal1 ;
   AntennaGateArea                            0.824400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656567 LAYER metal1 ; 
  END CI1

  PIN CO0
   AntennaPartialMetalArea                    1.897600 LAYER metal1 ;
   AntennaDiffArea                            1.923500 LAYER metal1 ;
  END CO0

  PIN CO1
   AntennaPartialMetalArea                    1.869600 LAYER metal1 ;
   AntennaDiffArea                            1.923500 LAYER metal1 ;
  END CO1

  PIN CS
   AntennaPartialMetalArea                    0.234800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.179288 LAYER metal1 ; 
  END CS

  PIN S
   AntennaPartialMetalArea                    0.572000 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END S

END FACS1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:32 CST 2007
#
#**********************************************************************




MACRO FACS2
  PIN A
   AntennaPartialMetalArea                    8.521200 LAYER metal1 ;
   AntennaGateArea                            0.633600 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.040436 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    7.101600 LAYER metal1 ;
   AntennaGateArea                            0.950400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656578 LAYER metal1 ; 
  END B

  PIN CI0
   AntennaPartialMetalArea                    2.966400 LAYER metal1 ;
   AntennaGateArea                            1.342800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.662245 LAYER metal1 ; 
  END CI0

  PIN CI1
   AntennaPartialMetalArea                    2.985600 LAYER metal1 ;
   AntennaGateArea                            1.342800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656566 LAYER metal1 ; 
  END CI1

  PIN CO0
   AntennaPartialMetalArea                    2.790400 LAYER metal1 ;
   AntennaDiffArea                            2.423750 LAYER metal1 ;
  END CO0

  PIN CO1
   AntennaPartialMetalArea                    2.745600 LAYER metal1 ;
   AntennaDiffArea                            2.423450 LAYER metal1 ;
  END CO1

  PIN CS
   AntennaPartialMetalArea                    0.279200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.406567 LAYER metal1 ; 
  END CS

  PIN S
   AntennaPartialMetalArea                    0.556800 LAYER metal1 ;
   AntennaDiffArea                            1.051450 LAYER metal1 ;
  END S

END FACS2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:36 CST 2007
#
#**********************************************************************




MACRO FACS2P
  PIN A
   AntennaPartialMetalArea                    8.648800 LAYER metal1 ;
   AntennaGateArea                            0.633600 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.040447 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    7.316000 LAYER metal1 ;
   AntennaGateArea                            0.950400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656589 LAYER metal1 ; 
  END B

  PIN CI0
   AntennaPartialMetalArea                    3.983400 LAYER metal1 ;
   AntennaGateArea                            2.368800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.662249 LAYER metal1 ; 
  END CI0

  PIN CI1
   AntennaPartialMetalArea                    3.763200 LAYER metal1 ;
   AntennaGateArea                            2.368800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656568 LAYER metal1 ; 
  END CI1

  PIN CO0
   AntennaPartialMetalArea                    4.428000 LAYER metal1 ;
   AntennaDiffArea                            4.749700 LAYER metal1 ;
  END CO0

  PIN CO1
   AntennaPartialMetalArea                    4.444800 LAYER metal1 ;
   AntennaDiffArea                            4.753900 LAYER metal1 ;
  END CO1

  PIN CS
   AntennaPartialMetalArea                    0.231200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.406562 LAYER metal1 ; 
  END CS

  PIN S
   AntennaPartialMetalArea                    0.845600 LAYER metal1 ;
   AntennaDiffArea                            1.378400 LAYER metal1 ;
  END S

END FACS2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:39 CST 2007
#
#**********************************************************************




MACRO FACS2S
  PIN A
   AntennaPartialMetalArea                    8.574000 LAYER metal1 ;
   AntennaGateArea                            0.633600 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.040403 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    7.490800 LAYER metal1 ;
   AntennaGateArea                            0.950400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.866166 LAYER metal1 ; 
  END B

  PIN CI0
   AntennaPartialMetalArea                    2.694400 LAYER metal1 ;
   AntennaGateArea                            0.824400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.662244 LAYER metal1 ; 
  END CI0

  PIN CI1
   AntennaPartialMetalArea                    2.787200 LAYER metal1 ;
   AntennaGateArea                            0.824400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.656567 LAYER metal1 ; 
  END CI1

  PIN CO0
   AntennaPartialMetalArea                    1.910400 LAYER metal1 ;
   AntennaDiffArea                            1.923500 LAYER metal1 ;
  END CO0

  PIN CO1
   AntennaPartialMetalArea                    1.856800 LAYER metal1 ;
   AntennaDiffArea                            1.923500 LAYER metal1 ;
  END CO1

  PIN CS
   AntennaPartialMetalArea                    0.449600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.179288 LAYER metal1 ; 
  END CS

  PIN S
   AntennaPartialMetalArea                    0.612800 LAYER metal1 ;
   AntennaDiffArea                            0.660000 LAYER metal1 ;
  END S

END FACS2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:43 CST 2007
#
#**********************************************************************




MACRO GCKETF
  PIN CK
   AntennaPartialMetalArea                    1.264800 LAYER metal1 ;
   AntennaGateArea                            1.027800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.055560 LAYER metal1 ; 
  END CK

  PIN E
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.198827 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    2.235400 LAYER metal1 ;
   AntennaDiffArea                            3.118400 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.194400 LAYER metal1 ;
   AntennaGateArea                            0.658800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.205528 LAYER metal1 ; 
  END TE

END GCKETF


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:46 CST 2007
#
#**********************************************************************




MACRO GCKETN
  PIN CK
   AntennaPartialMetalArea                    0.984000 LAYER metal1 ;
   AntennaGateArea                            0.518400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.756312 LAYER metal1 ; 
  END CK

  PIN E
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.252000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.977776 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.741400 LAYER metal1 ;
   AntennaDiffArea                            1.367100 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.216000 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.482780 LAYER metal1 ; 
  END TE

END GCKETN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:49 CST 2007
#
#**********************************************************************




MACRO GCKETP
  PIN CK
   AntennaPartialMetalArea                    1.082400 LAYER metal1 ;
   AntennaGateArea                            0.599400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.756314 LAYER metal1 ; 
  END CK

  PIN E
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.668059 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.825000 LAYER metal1 ;
   AntennaDiffArea                            1.506600 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.188000 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.197636 LAYER metal1 ; 
  END TE

END GCKETP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:51 CST 2007
#
#**********************************************************************




MACRO GCKETT
  PIN CK
   AntennaPartialMetalArea                    1.269600 LAYER metal1 ;
   AntennaGateArea                            0.775800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.666666 LAYER metal1 ; 
  END CK

  PIN E
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.313200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.309070 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    1.684600 LAYER metal1 ;
   AntennaDiffArea                            3.166100 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.230400 LAYER metal1 ;
   AntennaGateArea                            0.612000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227449 LAYER metal1 ; 
  END TE

END GCKETT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:54 CST 2007
#
#**********************************************************************




MACRO HA1
  PIN A
   AntennaPartialMetalArea                    1.037200 LAYER metal1 ;
   AntennaGateArea                            0.439200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.219514 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    2.824800 LAYER metal1 ;
   AntennaGateArea                            0.536400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.346991 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.741600 LAYER metal1 ;
   AntennaDiffArea                            1.395300 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.768400 LAYER metal1 ;
   AntennaDiffArea                            1.402200 LAYER metal1 ;
  END S

END HA1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:41:57 CST 2007
#
#**********************************************************************




MACRO HA1P
  PIN A
   AntennaPartialMetalArea                    0.308000 LAYER metal1 ;
   AntennaGateArea                            0.585000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.928884 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    1.855600 LAYER metal1 ;
   AntennaGateArea                            0.682800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.239897 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.774400 LAYER metal1 ;
   AntennaDiffArea                            1.391000 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.981600 LAYER metal1 ;
   AntennaDiffArea                            1.407000 LAYER metal1 ;
  END S

END HA1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:00 CST 2007
#
#**********************************************************************




MACRO HA1S
  PIN A
   AntennaPartialMetalArea                    1.062800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.165402 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    2.708800 LAYER metal1 ;
   AntennaGateArea                            0.475200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.231063 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.816800 LAYER metal1 ;
   AntennaDiffArea                            0.590000 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.874000 LAYER metal1 ;
   AntennaDiffArea                            0.598100 LAYER metal1 ;
  END S

END HA1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:03 CST 2007
#
#**********************************************************************




MACRO HA1T
  PIN A
   AntennaPartialMetalArea                    0.328000 LAYER metal1 ;
   AntennaGateArea                            0.585000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.951966 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    1.859400 LAYER metal1 ;
   AntennaGateArea                            0.682800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.239901 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    1.403200 LAYER metal1 ;
   AntennaDiffArea                            2.461500 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    1.293600 LAYER metal1 ;
   AntennaDiffArea                            2.637500 LAYER metal1 ;
  END S

END HA1T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:05 CST 2007
#
#**********************************************************************




MACRO HA2
  PIN A
   AntennaPartialMetalArea                    1.167600 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.258067 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    1.742800 LAYER metal1 ;
   AntennaGateArea                            1.237200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.944445 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    1.213600 LAYER metal1 ;
   AntennaDiffArea                            1.531600 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.768400 LAYER metal1 ;
   AntennaDiffArea                            1.234800 LAYER metal1 ;
  END S

END HA2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:08 CST 2007
#
#**********************************************************************




MACRO HA2P
  PIN A
   AntennaPartialMetalArea                    0.444800 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.258068 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    1.708800 LAYER metal1 ;
   AntennaGateArea                            2.167200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.065657 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    1.904800 LAYER metal1 ;
   AntennaDiffArea                            3.101000 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.760400 LAYER metal1 ;
   AntennaDiffArea                            1.228800 LAYER metal1 ;
  END S

END HA2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:10 CST 2007
#
#**********************************************************************




MACRO HA2T
  PIN A
   AntennaPartialMetalArea                    0.633600 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.208780 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    2.273600 LAYER metal1 ;
   AntennaGateArea                            3.043200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.065662 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    2.835200 LAYER metal1 ;
   AntennaDiffArea                            4.515400 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    1.398800 LAYER metal1 ;
   AntennaDiffArea                            2.463600 LAYER metal1 ;
  END S

END HA2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:13 CST 2007
#
#**********************************************************************




MACRO HA3
  PIN A
   AntennaPartialMetalArea                    1.324800 LAYER metal1 ;
   AntennaGateArea                            0.804600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.306448 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    1.780800 LAYER metal1 ;
   AntennaGateArea                            0.906000 LAYER metal1 ;
   AntennaMaxAreaCAR                          9.580837 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    1.048800 LAYER metal1 ;
   AntennaDiffArea                            2.166150 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.732400 LAYER metal1 ;
   AntennaDiffArea                            1.241800 LAYER metal1 ;
  END S

END HA3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:16 CST 2007
#
#**********************************************************************




MACRO HA3P
  PIN A
   AntennaPartialMetalArea                    1.288800 LAYER metal1 ;
   AntennaGateArea                            1.384200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.327011 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    2.221200 LAYER metal1 ;
   AntennaGateArea                            1.479600 LAYER metal1 ;
   AntennaMaxAreaCAR                          9.422983 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    1.302400 LAYER metal1 ;
   AntennaDiffArea                            2.732400 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.749200 LAYER metal1 ;
   AntennaDiffArea                            1.249800 LAYER metal1 ;
  END S

END HA3P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:19 CST 2007
#
#**********************************************************************




MACRO HA3T
  PIN A
   AntennaPartialMetalArea                    1.264800 LAYER metal1 ;
   AntennaGateArea                            1.949400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.327005 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    2.409200 LAYER metal1 ;
   AntennaGateArea                            2.044800 LAYER metal1 ;
   AntennaMaxAreaCAR                          9.422992 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    2.181600 LAYER metal1 ;
   AntennaDiffArea                            4.358000 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    1.801600 LAYER metal1 ;
   AntennaDiffArea                            2.448600 LAYER metal1 ;
  END S

END HA3T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:21 CST 2007
#
#**********************************************************************




MACRO INV1
  PIN I
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.518600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.671814 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.101400 LAYER metal1 ;
  END O

END INV1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:26 CST 2007
#
#**********************************************************************




MACRO INV12
  PIN I
   AntennaPartialMetalArea                    0.550400 LAYER metal1 ;
   AntennaGateArea                            5.630400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.908105 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                   11.726200 LAYER metal1 ;
   AntennaDiffArea                            7.146900 LAYER metal1 ;
  END O

END INV12


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:28 CST 2007
#
#**********************************************************************




MACRO INV12CK
  PIN I
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            5.362200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.234273 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                   17.873200 LAYER metal1 ;
   AntennaDiffArea                            8.268500 LAYER metal1 ;
  END O

END INV12CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:31 CST 2007
#
#**********************************************************************




MACRO INV1CK
  PIN I
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.369000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.293763 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.035000 LAYER metal1 ;
   AntennaDiffArea                            1.004500 LAYER metal1 ;
  END O

END INV1CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:34 CST 2007
#
#**********************************************************************




MACRO INV1S
  PIN I
   AntennaPartialMetalArea                    0.224400 LAYER metal1 ;
   AntennaGateArea                            0.314400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.657130 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.716800 LAYER metal1 ;
   AntennaDiffArea                            0.656800 LAYER metal1 ;
  END O

END INV1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:36 CST 2007
#
#**********************************************************************




MACRO INV2
  PIN I
   AntennaPartialMetalArea                    0.186200 LAYER metal1 ;
   AntennaGateArea                            0.876000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.185503 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.593600 LAYER metal1 ;
   AntennaDiffArea                            1.072200 LAYER metal1 ;
  END O

END INV2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:39 CST 2007
#
#**********************************************************************




MACRO INV2CK
  PIN I
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.826200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.328489 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.181000 LAYER metal1 ;
   AntennaDiffArea                            1.288800 LAYER metal1 ;
  END O

END INV2CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:42 CST 2007
#
#**********************************************************************




MACRO INV3
  PIN I
   AntennaPartialMetalArea                    0.182800 LAYER metal1 ;
   AntennaGateArea                            1.423200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.986507 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.751500 LAYER metal1 ;
   AntennaDiffArea                            2.165750 LAYER metal1 ;
  END O

END INV3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:44 CST 2007
#
#**********************************************************************




MACRO INV3CK
  PIN I
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            1.279800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.286612 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    3.510400 LAYER metal1 ;
   AntennaDiffArea                            2.392700 LAYER metal1 ;
  END O

END INV3CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:47 CST 2007
#
#**********************************************************************




MACRO INV4
  PIN I
   AntennaPartialMetalArea                    0.303200 LAYER metal1 ;
   AntennaGateArea                            1.941600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.957970 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    2.958000 LAYER metal1 ;
   AntennaDiffArea                            2.326300 LAYER metal1 ;
  END O

END INV4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:49 CST 2007
#
#**********************************************************************




MACRO INV4CK
  PIN I
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            1.729800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.269277 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    3.262800 LAYER metal1 ;
   AntennaDiffArea                            2.647200 LAYER metal1 ;
  END O

END INV4CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:52 CST 2007
#
#**********************************************************************




MACRO INV6
  PIN I
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            2.926800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.621563 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    6.801200 LAYER metal1 ;
   AntennaDiffArea                            3.665200 LAYER metal1 ;
  END O

END INV6


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:54 CST 2007
#
#**********************************************************************




MACRO INV6CK
  PIN I
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            2.640600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.258952 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    6.209000 LAYER metal1 ;
   AntennaDiffArea                            4.185400 LAYER metal1 ;
  END O

END INV6CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:56 CST 2007
#
#**********************************************************************




MACRO INV8
  PIN I
   AntennaPartialMetalArea                    0.526400 LAYER metal1 ;
   AntennaGateArea                            3.855600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.310871 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    8.194400 LAYER metal1 ;
   AntennaDiffArea                            4.864900 LAYER metal1 ;
  END O

END INV8


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:42:59 CST 2007
#
#**********************************************************************




MACRO INV8CK
  PIN I
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            3.547800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.246517 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    8.842800 LAYER metal1 ;
   AntennaDiffArea                            5.546200 LAYER metal1 ;
  END O

END INV8CK


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:02 CST 2007
#
#**********************************************************************




MACRO INVT1
  PIN E
   AntennaPartialMetalArea                    0.864800 LAYER metal1 ;
   AntennaGateArea                            0.428400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.303416 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.586800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.734828 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.931200 LAYER metal1 ;
   AntennaDiffArea                            1.380050 LAYER metal1 ;
  END O

END INVT1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:04 CST 2007
#
#**********************************************************************




MACRO INVT2
  PIN E
   AntennaPartialMetalArea                    0.906400 LAYER metal1 ;
   AntennaGateArea                            0.707400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.652688 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    1.849200 LAYER metal1 ;
   AntennaGateArea                            1.122000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.765962 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.156400 LAYER metal1 ;
   AntennaDiffArea                            1.233250 LAYER metal1 ;
  END O

END INVT2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:09 CST 2007
#
#**********************************************************************




MACRO INVT4
  PIN E
   AntennaPartialMetalArea                    1.221600 LAYER metal1 ;
   AntennaGateArea                            0.615600 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.170945 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.190400 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.255346 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.640700 LAYER metal1 ;
   AntennaDiffArea                            3.143450 LAYER metal1 ;
  END O

END INVT4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:11 CST 2007
#
#**********************************************************************




MACRO JKFN
  PIN CK
   AntennaPartialMetalArea                    0.249600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.335862 LAYER metal1 ; 
  END CK

  PIN J
   AntennaPartialMetalArea                    0.426400 LAYER metal1 ;
   AntennaGateArea                            0.234000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.749568 LAYER metal1 ; 
  END J

  PIN K
   AntennaPartialMetalArea                    0.447200 LAYER metal1 ;
   AntennaGateArea                            0.252000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.642067 LAYER metal1 ; 
  END K

  PIN Q
   AntennaPartialMetalArea                    0.890400 LAYER metal1 ;
   AntennaDiffArea                            1.061200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.505600 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

END JKFN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:14 CST 2007
#
#**********************************************************************




MACRO JKFRBN
  PIN CK
   AntennaPartialMetalArea                    0.618800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.093434 LAYER metal1 ; 
  END CK

  PIN J
   AntennaPartialMetalArea                    0.296000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.022723 LAYER metal1 ; 
  END J

  PIN K
   AntennaPartialMetalArea                    0.400000 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.089898 LAYER metal1 ; 
  END K

  PIN Q
   AntennaPartialMetalArea                    0.713200 LAYER metal1 ;
   AntennaDiffArea                            1.495900 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.528000 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.223200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.062505 LAYER metal1 ; 
  END RB

END JKFRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:18 CST 2007
#
#**********************************************************************




MACRO JKFRBP
  PIN CK
   AntennaPartialMetalArea                    0.618800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.093434 LAYER metal1 ; 
  END CK

  PIN J
   AntennaPartialMetalArea                    0.296000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.022723 LAYER metal1 ; 
  END J

  PIN K
   AntennaPartialMetalArea                    0.400000 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.089898 LAYER metal1 ; 
  END K

  PIN Q
   AntennaPartialMetalArea                    0.825600 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    1.002400 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.223200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.062505 LAYER metal1 ; 
  END RB

END JKFRBP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:21 CST 2007
#
#**********************************************************************




MACRO JKZN
  PIN CK
   AntennaPartialMetalArea                    0.255600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.603534 LAYER metal1 ; 
  END CK

  PIN J
   AntennaPartialMetalArea                    0.426400 LAYER metal1 ;
   AntennaGateArea                            0.234000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.757268 LAYER metal1 ; 
  END J

  PIN K
   AntennaPartialMetalArea                    0.435200 LAYER metal1 ;
   AntennaGateArea                            0.252000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.649206 LAYER metal1 ; 
  END K

  PIN Q
   AntennaPartialMetalArea                    0.893200 LAYER metal1 ;
   AntennaDiffArea                            1.063300 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.505600 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.311900 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227898 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.246400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.222224 LAYER metal1 ; 
  END TD

END JKZN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:25 CST 2007
#
#**********************************************************************




MACRO JKZRBN
  PIN CK
   AntennaPartialMetalArea                    0.643200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.142674 LAYER metal1 ; 
  END CK

  PIN J
   AntennaPartialMetalArea                    0.234400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.488632 LAYER metal1 ; 
  END J

  PIN K
   AntennaPartialMetalArea                    0.345600 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.041415 LAYER metal1 ; 
  END K

  PIN Q
   AntennaPartialMetalArea                    0.857200 LAYER metal1 ;
   AntennaDiffArea                            1.370300 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.760400 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.348000 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.785639 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.395200 LAYER metal1 ;
   AntennaGateArea                            0.439200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.256372 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.336000 LAYER metal1 ;
   AntennaGateArea                            0.280800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.358259 LAYER metal1 ; 
  END TD

END JKZRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:27 CST 2007
#
#**********************************************************************




MACRO JKZRBP
  PIN CK
   AntennaPartialMetalArea                    0.643200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.142674 LAYER metal1 ; 
  END CK

  PIN J
   AntennaPartialMetalArea                    0.234400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.488632 LAYER metal1 ; 
  END J

  PIN K
   AntennaPartialMetalArea                    0.345600 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.041415 LAYER metal1 ; 
  END K

  PIN Q
   AntennaPartialMetalArea                    0.653200 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.938000 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.348000 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.785639 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.395200 LAYER metal1 ;
   AntennaGateArea                            0.439200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.256372 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.336000 LAYER metal1 ;
   AntennaGateArea                            0.280800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.358259 LAYER metal1 ; 
  END TD

END JKZRBP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:30 CST 2007
#
#**********************************************************************




MACRO MAO222
  PIN A1
   AntennaPartialMetalArea                    0.180400 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.617042 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.516400 LAYER metal1 ;
   AntennaGateArea                            0.540000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.617034 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    1.300800 LAYER metal1 ;
   AntennaGateArea                            0.543600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.869154 LAYER metal1 ; 
  END C1

  PIN O
   AntennaPartialMetalArea                    0.682000 LAYER metal1 ;
   AntennaDiffArea                            1.630550 LAYER metal1 ;
  END O

END MAO222


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:34 CST 2007
#
#**********************************************************************




MACRO MAO222P
  PIN A1
   AntennaPartialMetalArea                    0.212000 LAYER metal1 ;
   AntennaGateArea                            0.410400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.989281 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.522000 LAYER metal1 ;
   AntennaGateArea                            0.820800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.989275 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    1.220000 LAYER metal1 ;
   AntennaGateArea                            0.824400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.989276 LAYER metal1 ; 
  END C1

  PIN O
   AntennaPartialMetalArea                    0.965600 LAYER metal1 ;
   AntennaDiffArea                            1.452900 LAYER metal1 ;
  END O

END MAO222P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:36 CST 2007
#
#**********************************************************************




MACRO MAO222S
  PIN A1
   AntennaPartialMetalArea                    0.207200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.556819 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.630400 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.414141 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    1.165600 LAYER metal1 ;
   AntennaGateArea                            0.320400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.761727 LAYER metal1 ; 
  END C1

  PIN O
   AntennaPartialMetalArea                    0.570000 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END MAO222S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:39 CST 2007
#
#**********************************************************************




MACRO MAO222T
  PIN A1
   AntennaPartialMetalArea                    0.212000 LAYER metal1 ;
   AntennaGateArea                            0.410400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.989281 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.522000 LAYER metal1 ;
   AntennaGateArea                            0.910800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.989277 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    1.208800 LAYER metal1 ;
   AntennaGateArea                            0.914400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.980680 LAYER metal1 ; 
  END C1

  PIN O
   AntennaPartialMetalArea                    1.210400 LAYER metal1 ;
   AntennaDiffArea                            2.691000 LAYER metal1 ;
  END O

END MAO222T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:42 CST 2007
#
#**********************************************************************




MACRO MAOI1
  PIN A1
   AntennaPartialMetalArea                    0.353500 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.808406 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.210700 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.687476 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.345400 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.073793 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.193600 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.526537 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.219600 LAYER metal1 ;
   AntennaDiffArea                            1.876700 LAYER metal1 ;
  END O

END MAOI1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:45 CST 2007
#
#**********************************************************************




MACRO MAOI1H
  PIN A1
   AntennaPartialMetalArea                    0.234800 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.282800 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.001064 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.306800 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.796233 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.314000 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.683939 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.470000 LAYER metal1 ;
   AntennaDiffArea                            2.842200 LAYER metal1 ;
  END O

END MAOI1H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:47 CST 2007
#
#**********************************************************************




MACRO MAOI1HP
  PIN A1
   AntennaPartialMetalArea                    0.229600 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            2.194200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.907845 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            1.018800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.692580 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            1.018800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753042 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    2.709200 LAYER metal1 ;
   AntennaDiffArea                            5.126400 LAYER metal1 ;
  END O

END MAOI1HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:50 CST 2007
#
#**********************************************************************




MACRO MAOI1HT
  PIN A1
   AntennaPartialMetalArea                    0.229600 LAYER metal1 ;
   AntennaGateArea                            3.317400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.781335 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            3.321000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.859982 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            1.528200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.770318 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            1.528200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.770318 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    3.724400 LAYER metal1 ;
   AntennaDiffArea                            7.265400 LAYER metal1 ;
  END O

END MAOI1HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:53 CST 2007
#
#**********************************************************************




MACRO MAOI1S
  PIN A1
   AntennaPartialMetalArea                    0.188800 LAYER metal1 ;
   AntennaGateArea                            0.230400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.412326 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.210700 LAYER metal1 ;
   AntennaGateArea                            0.230400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.144963 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.188600 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.241038 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.193600 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.649646 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.533200 LAYER metal1 ;
   AntennaDiffArea                            0.862400 LAYER metal1 ;
  END O

END MAOI1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:55 CST 2007
#
#**********************************************************************




MACRO MOAI1
  PIN A1
   AntennaPartialMetalArea                    0.220000 LAYER metal1 ;
   AntennaGateArea                            0.581400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.722053 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.186800 LAYER metal1 ;
   AntennaGateArea                            0.568300 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.786560 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.220500 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.223234 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.193600 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.015152 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.825600 LAYER metal1 ;
   AntennaDiffArea                            1.707150 LAYER metal1 ;
  END O

END MOAI1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:43:58 CST 2007
#
#**********************************************************************




MACRO MOAI1H
  PIN A1
   AntennaPartialMetalArea                    0.190000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.630103 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.322800 LAYER metal1 ;
   AntennaGateArea                            0.468000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.744446 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.294800 LAYER metal1 ;
   AntennaGateArea                            0.468000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.744445 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.855600 LAYER metal1 ;
   AntennaDiffArea                            3.380400 LAYER metal1 ;
  END O

END MOAI1H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:01 CST 2007
#
#**********************************************************************




MACRO MOAI1HP
  PIN A1
   AntennaPartialMetalArea                    0.190000 LAYER metal1 ;
   AntennaGateArea                            2.194200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.751435 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.680866 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    3.094000 LAYER metal1 ;
   AntennaDiffArea                            6.717900 LAYER metal1 ;
  END O

END MOAI1HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:04 CST 2007
#
#**********************************************************************




MACRO MOAI1HT
  PIN A1
   AntennaPartialMetalArea                    0.190000 LAYER metal1 ;
   AntennaGateArea                            3.267000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.793389 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            3.267000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.793388 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            1.690200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.696486 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            1.576800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.746575 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    4.265200 LAYER metal1 ;
   AntennaDiffArea                            9.990000 LAYER metal1 ;
  END O

END MOAI1HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:07 CST 2007
#
#**********************************************************************




MACRO MOAI1S
  PIN A1
   AntennaPartialMetalArea                    0.220800 LAYER metal1 ;
   AntennaGateArea                            0.205200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.818717 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.683200 LAYER metal1 ;
   AntennaGateArea                            0.203400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.054371 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.236000 LAYER metal1 ;
   AntennaGateArea                            0.160200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.320851 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.220800 LAYER metal1 ;
   AntennaGateArea                            0.160200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.590513 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.295800 LAYER metal1 ;
   AntennaDiffArea                            1.525500 LAYER metal1 ;
  END O

END MOAI1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:10 CST 2007
#
#**********************************************************************




MACRO MULBE
  PIN M
   AntennaPartialMetalArea                    0.816800 LAYER metal1 ;
   AntennaDiffArea                            1.096900 LAYER metal1 ;
  END M

  PIN M0
   AntennaPartialMetalArea                    0.554400 LAYER metal1 ;
   AntennaGateArea                            0.551400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.861809 LAYER metal1 ; 
  END M0

  PIN M1
   AntennaPartialMetalArea                    1.090400 LAYER metal1 ;
   AntennaGateArea                            0.551400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.550888 LAYER metal1 ; 
  END M1

  PIN M2
   AntennaPartialMetalArea                    0.560800 LAYER metal1 ;
   AntennaGateArea                            0.586200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.676770 LAYER metal1 ; 
  END M2

  PIN S
   AntennaPartialMetalArea                    0.816800 LAYER metal1 ;
   AntennaDiffArea                            1.096900 LAYER metal1 ;
  END S

  PIN Z
   AntennaPartialMetalArea                    0.912000 LAYER metal1 ;
   AntennaDiffArea                            1.096900 LAYER metal1 ;
  END Z

END MULBE


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:13 CST 2007
#
#**********************************************************************




MACRO MULBEP
  PIN M
   AntennaPartialMetalArea                    1.554000 LAYER metal1 ;
   AntennaDiffArea                            2.369800 LAYER metal1 ;
  END M

  PIN M0
   AntennaPartialMetalArea                    0.608000 LAYER metal1 ;
   AntennaGateArea                            0.551400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.861812 LAYER metal1 ; 
  END M0

  PIN M1
   AntennaPartialMetalArea                    1.076000 LAYER metal1 ;
   AntennaGateArea                            0.551400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.315594 LAYER metal1 ; 
  END M1

  PIN M2
   AntennaPartialMetalArea                    1.345400 LAYER metal1 ;
   AntennaGateArea                            1.218000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.823232 LAYER metal1 ; 
  END M2

  PIN S
   AntennaPartialMetalArea                    1.554000 LAYER metal1 ;
   AntennaDiffArea                            2.361800 LAYER metal1 ;
  END S

  PIN Z
   AntennaPartialMetalArea                    1.768800 LAYER metal1 ;
   AntennaDiffArea                            2.581800 LAYER metal1 ;
  END Z

END MULBEP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:16 CST 2007
#
#**********************************************************************




MACRO MULBET
  PIN M
   AntennaPartialMetalArea                    1.850400 LAYER metal1 ;
   AntennaDiffArea                            4.342000 LAYER metal1 ;
  END M

  PIN M0
   AntennaPartialMetalArea                    0.608000 LAYER metal1 ;
   AntennaGateArea                            0.551400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.861812 LAYER metal1 ; 
  END M0

  PIN M1
   AntennaPartialMetalArea                    1.076000 LAYER metal1 ;
   AntennaGateArea                            0.551400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.315594 LAYER metal1 ; 
  END M1

  PIN M2
   AntennaPartialMetalArea                    0.392800 LAYER metal1 ;
   AntennaGateArea                            2.335200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.067062 LAYER metal1 ; 
  END M2

  PIN S
   AntennaPartialMetalArea                    1.836000 LAYER metal1 ;
   AntennaDiffArea                            4.239600 LAYER metal1 ;
  END S

  PIN Z
   AntennaPartialMetalArea                    1.886800 LAYER metal1 ;
   AntennaDiffArea                            4.287600 LAYER metal1 ;
  END Z

END MULBET


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:19 CST 2007
#
#**********************************************************************




MACRO MULPA
  PIN M
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.141972 LAYER metal1 ; 
  END M

  PIN M0
   AntennaPartialMetalArea                    0.354400 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.219982 LAYER metal1 ; 
  END M0

  PIN M1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.775534 LAYER metal1 ; 
  END M1

  PIN P
   AntennaPartialMetalArea                    0.620400 LAYER metal1 ;
   AntennaDiffArea                            1.489100 LAYER metal1 ;
  END P

  PIN S
   AntennaPartialMetalArea                    0.470400 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.957355 LAYER metal1 ; 
  END S

  PIN Z
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277777 LAYER metal1 ; 
  END Z

END MULPA


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:22 CST 2007
#
#**********************************************************************




MACRO MULPAP
  PIN M
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.141972 LAYER metal1 ; 
  END M

  PIN M0
   AntennaPartialMetalArea                    0.354400 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.219982 LAYER metal1 ; 
  END M0

  PIN M1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.775534 LAYER metal1 ; 
  END M1

  PIN P
   AntennaPartialMetalArea                    0.660400 LAYER metal1 ;
   AntennaDiffArea                            1.533400 LAYER metal1 ;
  END P

  PIN S
   AntennaPartialMetalArea                    0.482400 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.942195 LAYER metal1 ; 
  END S

  PIN Z
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277777 LAYER metal1 ; 
  END Z

END MULPAP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:25 CST 2007
#
#**********************************************************************




MACRO MULPAT
  PIN M
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.141972 LAYER metal1 ; 
  END M

  PIN M0
   AntennaPartialMetalArea                    0.354400 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.219982 LAYER metal1 ; 
  END M0

  PIN M1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.775534 LAYER metal1 ; 
  END M1

  PIN P
   AntennaPartialMetalArea                    1.584800 LAYER metal1 ;
   AntennaDiffArea                            3.012800 LAYER metal1 ;
  END P

  PIN S
   AntennaPartialMetalArea                    0.538400 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.942198 LAYER metal1 ; 
  END S

  PIN Z
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277777 LAYER metal1 ; 
  END Z

END MULPAT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:28 CST 2007
#
#**********************************************************************




MACRO MUX2
  PIN A
   AntennaPartialMetalArea                    0.526400 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.232324 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.324000 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.959596 LAYER metal1 ; 
  END B

  PIN O
   AntennaPartialMetalArea                    0.604100 LAYER metal1 ;
   AntennaDiffArea                            1.356500 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.428000 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681190 LAYER metal1 ; 
  END S

END MUX2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:30 CST 2007
#
#**********************************************************************




MACRO MUX2F
  PIN A
   AntennaPartialMetalArea                    0.509200 LAYER metal1 ;
   AntennaGateArea                            0.419400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.886505 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.419400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.944686 LAYER metal1 ; 
  END B

  PIN O
   AntennaPartialMetalArea                    1.436000 LAYER metal1 ;
   AntennaDiffArea                            2.804800 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.427600 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.700811 LAYER metal1 ; 
  END S

END MUX2F


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:33 CST 2007
#
#**********************************************************************




MACRO MUX2P
  PIN A
   AntennaPartialMetalArea                    0.789600 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.867386 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.324000 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.817207 LAYER metal1 ; 
  END B

  PIN O
   AntennaPartialMetalArea                    1.010800 LAYER metal1 ;
   AntennaDiffArea                            1.375000 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.317800 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.244210 LAYER metal1 ; 
  END S

END MUX2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:36 CST 2007
#
#**********************************************************************




MACRO MUX2S
  PIN A
   AntennaPartialMetalArea                    0.238000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.643935 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.790399 LAYER metal1 ; 
  END B

  PIN O
   AntennaPartialMetalArea                    0.878000 LAYER metal1 ;
   AntennaDiffArea                            0.602700 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.716800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.150254 LAYER metal1 ; 
  END S

END MUX2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:39 CST 2007
#
#**********************************************************************




MACRO MUX2T
  PIN A
   AntennaPartialMetalArea                    0.489200 LAYER metal1 ;
   AntennaGateArea                            0.414000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.898067 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.419400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.944686 LAYER metal1 ; 
  END B

  PIN O
   AntennaPartialMetalArea                    1.336000 LAYER metal1 ;
   AntennaDiffArea                            2.600150 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.430400 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.700810 LAYER metal1 ; 
  END S

END MUX2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:42 CST 2007
#
#**********************************************************************




MACRO MUX3
  PIN A
   AntennaPartialMetalArea                    0.340400 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.451903 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.237200 LAYER metal1 ;
   AntennaGateArea                            0.247800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.565776 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.296800 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.050510 LAYER metal1 ; 
  END C

  PIN O
   AntennaPartialMetalArea                    0.670000 LAYER metal1 ;
   AntennaDiffArea                            1.338600 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.545800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.653406 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.375600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.241794 LAYER metal1 ; 
  END S1

END MUX3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:46 CST 2007
#
#**********************************************************************




MACRO MUX3P
  PIN A
   AntennaPartialMetalArea                    0.340400 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.451903 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.242800 LAYER metal1 ;
   AntennaGateArea                            0.247800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.565778 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.361200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.050508 LAYER metal1 ; 
  END C

  PIN O
   AntennaPartialMetalArea                    1.008000 LAYER metal1 ;
   AntennaDiffArea                            1.431900 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.551500 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.653404 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.375600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.109214 LAYER metal1 ; 
  END S1

END MUX3P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:50 CST 2007
#
#**********************************************************************




MACRO MUX3S
  PIN A
   AntennaPartialMetalArea                    0.270100 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.702988 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.119662 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.207200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.699499 LAYER metal1 ; 
  END C

  PIN O
   AntennaPartialMetalArea                    1.130000 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.457600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.542296 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.270800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.327812 LAYER metal1 ; 
  END S1

END MUX3S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:53 CST 2007
#
#**********************************************************************




MACRO MUX3T
  PIN A
   AntennaPartialMetalArea                    0.352400 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.451912 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.247800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.565778 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.337200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.050510 LAYER metal1 ; 
  END C

  PIN O
   AntennaPartialMetalArea                    1.272000 LAYER metal1 ;
   AntennaDiffArea                            2.755350 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.492400 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.653407 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.375600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.055394 LAYER metal1 ; 
  END S1

END MUX3T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:44:57 CST 2007
#
#**********************************************************************




MACRO MUX4
  PIN A
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.141972 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277777 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.214400 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.164202 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.153084 LAYER metal1 ; 
  END D

  PIN O
   AntennaPartialMetalArea                    0.620400 LAYER metal1 ;
   AntennaDiffArea                            1.489100 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.525600 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.731356 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.916944 LAYER metal1 ; 
  END S1

END MUX4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:01 CST 2007
#
#**********************************************************************




MACRO MUX4P
  PIN A
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.259200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.344138 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.259200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.513886 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.235200 LAYER metal1 ;
   AntennaGateArea                            0.259200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.344133 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.259200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.479942 LAYER metal1 ; 
  END D

  PIN O
   AntennaPartialMetalArea                    0.697600 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.554400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.563488 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.129064 LAYER metal1 ; 
  END S1

END MUX4P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:05 CST 2007
#
#**********************************************************************




MACRO MUX4S
  PIN A
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.754480 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.951609 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.770611 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.754483 LAYER metal1 ; 
  END D

  PIN O
   AntennaPartialMetalArea                    0.620400 LAYER metal1 ;
   AntennaDiffArea                            0.672000 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.514800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.725714 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.856344 LAYER metal1 ; 
  END S1

END MUX4S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:09 CST 2007
#
#**********************************************************************




MACRO MUX4T
  PIN A
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.259200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.344138 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.259200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.513886 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.235200 LAYER metal1 ;
   AntennaGateArea                            0.259200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.344133 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.259200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.479942 LAYER metal1 ; 
  END D

  PIN O
   AntennaPartialMetalArea                    1.218400 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.554400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.563488 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.231200 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.028061 LAYER metal1 ; 
  END S1

END MUX4T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:13 CST 2007
#
#**********************************************************************




MACRO MUXB2
  PIN A
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.986867 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.986869 LAYER metal1 ; 
  END B

  PIN EB
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.471600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.792193 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    0.815600 LAYER metal1 ;
   AntennaDiffArea                            1.323800 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.815658 LAYER metal1 ; 
  END S

END MUXB2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:16 CST 2007
#
#**********************************************************************




MACRO MUXB2P
  PIN A
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.986867 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.986868 LAYER metal1 ; 
  END B

  PIN EB
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.946800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.794677 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    1.478800 LAYER metal1 ;
   AntennaDiffArea                            2.439000 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.815658 LAYER metal1 ; 
  END S

END MUXB2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:19 CST 2007
#
#**********************************************************************




MACRO MUXB2S
  PIN A
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.325054 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.325058 LAYER metal1 ; 
  END B

  PIN EB
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.150292 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    0.818400 LAYER metal1 ;
   AntennaDiffArea                            0.961000 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.815658 LAYER metal1 ; 
  END S

END MUXB2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:23 CST 2007
#
#**********************************************************************




MACRO MUXB2T
  PIN A
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.986867 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.986868 LAYER metal1 ; 
  END B

  PIN EB
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            1.420200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.828897 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    1.702000 LAYER metal1 ;
   AntennaDiffArea                            3.180900 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.815658 LAYER metal1 ; 
  END S

END MUXB2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:26 CST 2007
#
#**********************************************************************




MACRO MUXB4
  PIN A
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.560930 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.758069 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.239200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.560935 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.718643 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.473400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.857622 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    0.972400 LAYER metal1 ;
   AntennaDiffArea                            1.392700 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.496800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.041871 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.327600 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.700851 LAYER metal1 ; 
  END S1

END MUXB4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:30 CST 2007
#
#**********************************************************************




MACRO MUXB4P
  PIN A
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.560930 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.758069 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.239200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.560935 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.718643 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.946800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.759189 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    1.511600 LAYER metal1 ;
   AntennaDiffArea                            2.657400 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.496800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.041871 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.263200 LAYER metal1 ;
   AntennaGateArea                            0.327600 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.492061 LAYER metal1 ; 
  END S1

END MUXB4P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:34 CST 2007
#
#**********************************************************************




MACRO MUXB4S
  PIN A
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.560930 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.758069 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.239200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.560935 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.718643 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.187133 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    0.916400 LAYER metal1 ;
   AntennaDiffArea                            1.009000 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.496800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.041871 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.327600 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.700851 LAYER metal1 ; 
  END S1

END MUXB4S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:38 CST 2007
#
#**********************************************************************




MACRO MUXB4T
  PIN A
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.560930 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.758069 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.239200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.560935 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.223200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.718643 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.420200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.835094 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    1.660400 LAYER metal1 ;
   AntennaDiffArea                            3.180900 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.496800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.041871 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.263200 LAYER metal1 ;
   AntennaGateArea                            0.327600 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.492061 LAYER metal1 ; 
  END S1

END MUXB4T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:41 CST 2007
#
#**********************************************************************




MACRO MXL2H
  PIN A
   AntennaPartialMetalArea                    0.275200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.735535 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.275200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.735535 LAYER metal1 ; 
  END B

  PIN OB
   AntennaPartialMetalArea                    2.145600 LAYER metal1 ;
   AntennaDiffArea                            4.221900 LAYER metal1 ;
  END OB

  PIN S
   AntennaPartialMetalArea                    0.193600 LAYER metal1 ;
   AntennaGateArea                            1.602000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.030461 LAYER metal1 ; 
  END S

END MXL2H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:44 CST 2007
#
#**********************************************************************




MACRO MXL2HF
  PIN A
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            4.507200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.816294 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            4.507200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784345 LAYER metal1 ; 
  END B

  PIN OB
   AntennaPartialMetalArea                    6.144000 LAYER metal1 ;
   AntennaDiffArea                           14.182700 LAYER metal1 ;
  END OB

  PIN S
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            6.400800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.927040 LAYER metal1 ; 
  END S

END MXL2HF


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:47 CST 2007
#
#**********************************************************************




MACRO MXL2HP
  PIN A
   AntennaPartialMetalArea                    0.232800 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END B

  PIN OB
   AntennaPartialMetalArea                    3.370800 LAYER metal1 ;
   AntennaDiffArea                            7.541200 LAYER metal1 ;
  END OB

  PIN S
   AntennaPartialMetalArea                    0.275200 LAYER metal1 ;
   AntennaGateArea                            3.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.939447 LAYER metal1 ; 
  END S

END MXL2HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:50 CST 2007
#
#**********************************************************************




MACRO MXL2HS
  PIN A
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.673056 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.673056 LAYER metal1 ; 
  END B

  PIN OB
   AntennaPartialMetalArea                    0.890400 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END OB

  PIN S
   AntennaPartialMetalArea                    0.185600 LAYER metal1 ;
   AntennaGateArea                            0.846000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.128845 LAYER metal1 ; 
  END S

END MXL2HS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:54 CST 2007
#
#**********************************************************************




MACRO MXL2HT
  PIN A
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.821086 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.193200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END B

  PIN OB
   AntennaPartialMetalArea                    4.818000 LAYER metal1 ;
   AntennaDiffArea                           11.061700 LAYER metal1 ;
  END OB

  PIN S
   AntennaPartialMetalArea                    0.275200 LAYER metal1 ;
   AntennaGateArea                            4.806000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.953638 LAYER metal1 ; 
  END S

END MXL2HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:45:58 CST 2007
#
#**********************************************************************




MACRO MXL3
  PIN A
   AntennaPartialMetalArea                    0.269600 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.523234 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.004043 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.866157 LAYER metal1 ; 
  END C

  PIN OB
   AntennaPartialMetalArea                    0.609200 LAYER metal1 ;
   AntennaDiffArea                            1.278600 LAYER metal1 ;
  END OB

  PIN S0
   AntennaPartialMetalArea                    0.504800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.493056 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.282000 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.712278 LAYER metal1 ; 
  END S1

END MXL3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:01 CST 2007
#
#**********************************************************************




MACRO MXL3P
  PIN A
   AntennaPartialMetalArea                    0.275200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.523231 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.004043 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.782827 LAYER metal1 ; 
  END C

  PIN OB
   AntennaPartialMetalArea                    0.580000 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END OB

  PIN S0
   AntennaPartialMetalArea                    0.507600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.493057 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.254000 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.731222 LAYER metal1 ; 
  END S1

END MXL3P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:05 CST 2007
#
#**********************************************************************




MACRO MXL3S
  PIN A
   AntennaPartialMetalArea                    0.269600 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.523234 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.004043 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.866157 LAYER metal1 ; 
  END C

  PIN OB
   AntennaPartialMetalArea                    0.956400 LAYER metal1 ;
   AntennaDiffArea                            0.769300 LAYER metal1 ;
  END OB

  PIN S0
   AntennaPartialMetalArea                    0.504800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.493056 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.254000 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.731222 LAYER metal1 ; 
  END S1

END MXL3S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:08 CST 2007
#
#**********************************************************************




MACRO MXL3T
  PIN A
   AntennaPartialMetalArea                    0.286400 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.523235 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.004043 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.782827 LAYER metal1 ; 
  END C

  PIN OB
   AntennaPartialMetalArea                    1.180000 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END OB

  PIN S0
   AntennaPartialMetalArea                    0.504800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.493056 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.254000 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.731222 LAYER metal1 ; 
  END S1

END MXL3T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:12 CST 2007
#
#**********************************************************************




MACRO ND2
  PIN I1
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.418800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.000000 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.418800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.000004 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.747600 LAYER metal1 ;
   AntennaDiffArea                            1.079900 LAYER metal1 ;
  END O

END ND2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:16 CST 2007
#
#**********************************************************************




MACRO ND2F
  PIN I1
   AntennaPartialMetalArea                    0.963200 LAYER metal1 ;
   AntennaGateArea                            2.274000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.969449 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.162800 LAYER metal1 ;
   AntennaGateArea                            2.150400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.943493 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    3.362000 LAYER metal1 ;
   AntennaDiffArea                            5.207550 LAYER metal1 ;
  END O

END ND2F


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:19 CST 2007
#
#**********************************************************************




MACRO ND2P
  PIN I1
   AntennaPartialMetalArea                    0.220400 LAYER metal1 ;
   AntennaGateArea                            1.068000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.765730 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.204400 LAYER metal1 ;
   AntennaGateArea                            1.062600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.771316 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.337200 LAYER metal1 ;
   AntennaDiffArea                            2.587350 LAYER metal1 ;
  END O

END ND2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:22 CST 2007
#
#**********************************************************************




MACRO ND2S
  PIN I1
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.343200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.267485 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.343200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.267485 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.742000 LAYER metal1 ;
   AntennaDiffArea                            0.896300 LAYER metal1 ;
  END O

END ND2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:26 CST 2007
#
#**********************************************************************




MACRO ND2T
  PIN I1
   AntennaPartialMetalArea                    0.939200 LAYER metal1 ;
   AntennaGateArea                            1.717800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.039684 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.822200 LAYER metal1 ;
   AntennaGateArea                            1.656000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.553178 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    2.681000 LAYER metal1 ;
   AntennaDiffArea                            3.849150 LAYER metal1 ;
  END O

END ND2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:29 CST 2007
#
#**********************************************************************




MACRO ND3
  PIN I1
   AntennaPartialMetalArea                    0.200000 LAYER metal1 ;
   AntennaGateArea                            0.471000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.001272 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.212000 LAYER metal1 ;
   AntennaGateArea                            0.472200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.772558 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.184000 LAYER metal1 ;
   AntennaGateArea                            0.484200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.728622 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.105600 LAYER metal1 ;
   AntennaDiffArea                            1.668350 LAYER metal1 ;
  END O

END ND3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:32 CST 2007
#
#**********************************************************************




MACRO ND3HT
  PIN I1
   AntennaPartialMetalArea                    0.261800 LAYER metal1 ;
   AntennaGateArea                            1.501200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784172 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.223600 LAYER metal1 ;
   AntennaGateArea                            1.501200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784172 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.252000 LAYER metal1 ;
   AntennaGateArea                            1.443600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.888616 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    2.457600 LAYER metal1 ;
   AntennaDiffArea                            5.261000 LAYER metal1 ;
  END O

END ND3HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:35 CST 2007
#
#**********************************************************************




MACRO ND3P
  PIN I1
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.977400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.965827 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.068000 LAYER metal1 ;
   AntennaGateArea                            1.011000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.897760 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    1.268700 LAYER metal1 ;
   AntennaGateArea                            0.988800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.887140 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    2.234000 LAYER metal1 ;
   AntennaDiffArea                            2.826000 LAYER metal1 ;
  END O

END ND3P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:38 CST 2007
#
#**********************************************************************




MACRO ND3S
  PIN I1
   AntennaPartialMetalArea                    0.188000 LAYER metal1 ;
   AntennaGateArea                            0.302400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.785057 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.244000 LAYER metal1 ;
   AntennaGateArea                            0.302400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.479502 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.208000 LAYER metal1 ;
   AntennaGateArea                            0.302400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.523149 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.165400 LAYER metal1 ;
   AntennaDiffArea                            1.183250 LAYER metal1 ;
  END O

END ND3S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:42 CST 2007
#
#**********************************************************************




MACRO ND4
  PIN I1
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.607322 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.243200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.857326 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.199200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.176764 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.361107 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.774400 LAYER metal1 ;
   AntennaDiffArea                            1.460400 LAYER metal1 ;
  END O

END ND4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:46 CST 2007
#
#**********************************************************************




MACRO ND4P
  PIN I1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.584263 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.243200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.329634 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.746296 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.716670 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    1.080500 LAYER metal1 ;
   AntennaDiffArea                            1.440800 LAYER metal1 ;
  END O

END ND4P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:49 CST 2007
#
#**********************************************************************




MACRO ND4S
  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.392677 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.215200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.256314 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.199200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.438134 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.574497 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.858400 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END ND4S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:53 CST 2007
#
#**********************************************************************




MACRO ND4T
  PIN I1
   AntennaPartialMetalArea                    0.232400 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.182774 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.205200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.345560 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.206400 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.742777 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.729448 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    1.335600 LAYER metal1 ;
   AntennaDiffArea                            2.677200 LAYER metal1 ;
  END O

END ND4T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:46:57 CST 2007
#
#**********************************************************************




MACRO NR2
  PIN I1
   AntennaPartialMetalArea                    0.196800 LAYER metal1 ;
   AntennaGateArea                            0.439800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.877674 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.205200 LAYER metal1 ;
   AntennaGateArea                            0.439800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.033194 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.716800 LAYER metal1 ;
   AntennaDiffArea                            1.211050 LAYER metal1 ;
  END O

END NR2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:01 CST 2007
#
#**********************************************************************




MACRO NR2F
  PIN I1
   AntennaPartialMetalArea                    1.644800 LAYER metal1 ;
   AntennaGateArea                            2.463600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.859399 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.639900 LAYER metal1 ;
   AntennaGateArea                            2.458800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.015829 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    4.631800 LAYER metal1 ;
   AntennaDiffArea                            5.111300 LAYER metal1 ;
  END O

END NR2F


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:04 CST 2007
#
#**********************************************************************




MACRO NR2P
  PIN I1
   AntennaPartialMetalArea                    0.300000 LAYER metal1 ;
   AntennaGateArea                            0.905400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.011045 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.214000 LAYER metal1 ;
   AntennaGateArea                            0.907200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.234647 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    2.848600 LAYER metal1 ;
   AntennaDiffArea                            2.781900 LAYER metal1 ;
  END O

END NR2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:07 CST 2007
#
#**********************************************************************




MACRO NR2T
  PIN I1
   AntennaPartialMetalArea                    0.923900 LAYER metal1 ;
   AntennaGateArea                            1.342800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.857370 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.921600 LAYER metal1 ;
   AntennaGateArea                            1.342800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.047013 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    2.725200 LAYER metal1 ;
   AntennaDiffArea                            3.159000 LAYER metal1 ;
  END O

END NR2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:10 CST 2007
#
#**********************************************************************




MACRO NR3
  PIN I1
   AntennaPartialMetalArea                    0.312000 LAYER metal1 ;
   AntennaGateArea                            0.408600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.183067 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.209200 LAYER metal1 ;
   AntennaGateArea                            0.408600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.091038 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.408600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.165443 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.203200 LAYER metal1 ;
   AntennaDiffArea                            2.413700 LAYER metal1 ;
  END O

END NR3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:14 CST 2007
#
#**********************************************************************




MACRO NR3H
  PIN I1
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.768600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.791565 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.278800 LAYER metal1 ;
   AntennaGateArea                            0.831600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731603 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.334800 LAYER metal1 ;
   AntennaGateArea                            0.831600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731603 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.615200 LAYER metal1 ;
   AntennaDiffArea                            2.399400 LAYER metal1 ;
  END O

END NR3H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:17 CST 2007
#
#**********************************************************************




MACRO NR3HP
  PIN I1
   AntennaPartialMetalArea                    0.198800 LAYER metal1 ;
   AntennaGateArea                            1.184400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.984801 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            1.184400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.984800 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.370800 LAYER metal1 ;
   AntennaGateArea                            1.247400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.865802 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    2.174400 LAYER metal1 ;
   AntennaDiffArea                            3.051300 LAYER metal1 ;
  END O

END NR3HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:21 CST 2007
#
#**********************************************************************




MACRO NR3HT
  PIN I1
   AntennaPartialMetalArea                    0.198800 LAYER metal1 ;
   AntennaGateArea                            2.431800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.985940 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            2.431800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.985932 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.370800 LAYER metal1 ;
   AntennaGateArea                            2.431800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.985940 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    4.173600 LAYER metal1 ;
   AntennaDiffArea                            5.255400 LAYER metal1 ;
  END O

END NR3HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:24 CST 2007
#
#**********************************************************************




MACRO NR4
  PIN I1
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.950245 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.314000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.071306 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.178600 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.715586 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.253800 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.690711 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END O

END NR4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:28 CST 2007
#
#**********************************************************************




MACRO NR4P
  PIN I1
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.940295 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.356000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.019066 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.843287 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.263200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.110279 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.593600 LAYER metal1 ;
   AntennaDiffArea                            1.456600 LAYER metal1 ;
  END O

END NR4P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:32 CST 2007
#
#**********************************************************************




MACRO NR4S
  PIN I1
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.108621 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.190000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.154232 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.251200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.166671 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.436977 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END NR4S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:35 CST 2007
#
#**********************************************************************




MACRO NR4T
  PIN I1
   AntennaPartialMetalArea                    0.254800 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.940295 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.356000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.019066 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.843287 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.263200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.110279 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    1.092400 LAYER metal1 ;
   AntennaDiffArea                            2.690400 LAYER metal1 ;
  END O

END NR4T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:38 CST 2007
#
#**********************************************************************




MACRO OA112
  PIN A1
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.237600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.966329 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.359200 LAYER metal1 ;
   AntennaGateArea                            0.237600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.125425 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.359200 LAYER metal1 ;
   AntennaGateArea                            0.336600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.715388 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.299600 LAYER metal1 ;
   AntennaGateArea                            0.336600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.190133 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.971200 LAYER metal1 ;
   AntennaDiffArea                            1.593250 LAYER metal1 ;
  END O

END OA112


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:42 CST 2007
#
#**********************************************************************




MACRO OA112P
  PIN A1
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.279000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.668097 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.348000 LAYER metal1 ;
   AntennaGateArea                            0.279000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.810038 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.348000 LAYER metal1 ;
   AntennaGateArea                            0.414000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.368600 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.305200 LAYER metal1 ;
   AntennaGateArea                            0.414000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.967632 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.806800 LAYER metal1 ;
   AntennaDiffArea                            1.928100 LAYER metal1 ;
  END O

END OA112P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:45 CST 2007
#
#**********************************************************************




MACRO OA112S
  PIN A1
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.279038 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.359200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.517673 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.359200 LAYER metal1 ;
   AntennaGateArea                            0.205200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.147173 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.205200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.285570 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.817200 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END OA112S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:49 CST 2007
#
#**********************************************************************




MACRO OA112T
  PIN A1
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.306000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.520918 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.334000 LAYER metal1 ;
   AntennaGateArea                            0.306000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.650327 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.334000 LAYER metal1 ;
   AntennaGateArea                            0.486000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.132507 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.305200 LAYER metal1 ;
   AntennaGateArea                            0.486000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.824276 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.356000 LAYER metal1 ;
   AntennaDiffArea                            3.278800 LAYER metal1 ;
  END O

END OA112T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:53 CST 2007
#
#**********************************************************************




MACRO OA12
  PIN A1
   AntennaPartialMetalArea                    0.286800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.630339 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.238800 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.096190 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.428800 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.041462 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.657600 LAYER metal1 ;
   AntennaDiffArea                            1.321700 LAYER metal1 ;
  END O

END OA12


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:56 CST 2007
#
#**********************************************************************




MACRO OA12P
  PIN A1
   AntennaPartialMetalArea                    0.295200 LAYER metal1 ;
   AntennaGateArea                            0.379800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.922069 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.216000 LAYER metal1 ;
   AntennaGateArea                            0.491400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.764750 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.491400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.934879 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.839600 LAYER metal1 ;
   AntennaDiffArea                            1.554600 LAYER metal1 ;
  END O

END OA12P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:47:59 CST 2007
#
#**********************************************************************




MACRO OA12S
  PIN A1
   AntennaPartialMetalArea                    0.282800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.097226 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.322800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.691241 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.275200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.620725 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.931200 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END OA12S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:02 CST 2007
#
#**********************************************************************




MACRO OA12T
  PIN A1
   AntennaPartialMetalArea                    0.295200 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.926458 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.216000 LAYER metal1 ;
   AntennaGateArea                            0.486000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.765846 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.486000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.937864 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.192000 LAYER metal1 ;
   AntennaDiffArea                            2.659200 LAYER metal1 ;
  END O

END OA12T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:06 CST 2007
#
#**********************************************************************




MACRO OA13
  PIN A1
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            0.217800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.723598 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.197200 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.039687 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.239400 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.997887 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.234000 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.202642 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.774400 LAYER metal1 ;
   AntennaDiffArea                            1.165100 LAYER metal1 ;
  END O

END OA13


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:10 CST 2007
#
#**********************************************************************




MACRO OA13P
  PIN A1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.262800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.431128 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.197200 LAYER metal1 ;
   AntennaGateArea                            0.460800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.814669 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.239400 LAYER metal1 ;
   AntennaGateArea                            0.460800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.814669 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.234000 LAYER metal1 ;
   AntennaGateArea                            0.460800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.986547 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.540000 LAYER metal1 ;
   AntennaDiffArea                            1.488100 LAYER metal1 ;
  END O

END OA13P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:14 CST 2007
#
#**********************************************************************




MACRO OA13S
  PIN A1
   AntennaPartialMetalArea                    0.364800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.861112 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.225200 LAYER metal1 ;
   AntennaGateArea                            0.313200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.112391 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.368000 LAYER metal1 ;
   AntennaGateArea                            0.313200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.112392 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.427800 LAYER metal1 ;
   AntennaGateArea                            0.313200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.154530 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.778400 LAYER metal1 ;
   AntennaDiffArea                            0.597800 LAYER metal1 ;
  END O

END OA13S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:18 CST 2007
#
#**********************************************************************




MACRO OA13T
  PIN A1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.262800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.431128 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.197200 LAYER metal1 ;
   AntennaGateArea                            0.460800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.814669 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.239400 LAYER metal1 ;
   AntennaGateArea                            0.460800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.814669 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.234000 LAYER metal1 ;
   AntennaGateArea                            0.460800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.986547 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    1.108000 LAYER metal1 ;
   AntennaDiffArea                            2.706750 LAYER metal1 ;
  END O

END OA13T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:22 CST 2007
#
#**********************************************************************




MACRO OA22
  PIN A1
   AntennaPartialMetalArea                    0.301600 LAYER metal1 ;
   AntennaGateArea                            0.250200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.333334 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.340000 LAYER metal1 ;
   AntennaGateArea                            0.250200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609117 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.185600 LAYER metal1 ;
   AntennaGateArea                            0.250200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.193843 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.202400 LAYER metal1 ;
   AntennaGateArea                            0.250200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.111907 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.971200 LAYER metal1 ;
   AntennaDiffArea                            1.253400 LAYER metal1 ;
  END O

END OA22


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:26 CST 2007
#
#**********************************************************************




MACRO OA222
  PIN A1
   AntennaPartialMetalArea                    0.360000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.612773 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.296000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.223053 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.239400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.462819 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.300000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.626039 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.116090 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.296000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.108623 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.931200 LAYER metal1 ;
   AntennaDiffArea                            1.335400 LAYER metal1 ;
  END O

END OA222


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:30 CST 2007
#
#**********************************************************************




MACRO OA222P
  PIN A1
   AntennaPartialMetalArea                    0.324000 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.086420 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.324000 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.167900 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.322200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.936688 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.080862 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.325800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.295887 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.325800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.390422 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.911200 LAYER metal1 ;
   AntennaDiffArea                            1.456700 LAYER metal1 ;
  END O

END OA222P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:34 CST 2007
#
#**********************************************************************




MACRO OA222S
  PIN A1
   AntennaPartialMetalArea                    0.360000 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.366453 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.296000 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.036323 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.185400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.471412 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.300000 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.393166 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.316000 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.688036 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.292000 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.678421 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.931200 LAYER metal1 ;
   AntennaDiffArea                            0.592900 LAYER metal1 ;
  END O

END OA222S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:37 CST 2007
#
#**********************************************************************




MACRO OA222T
  PIN A1
   AntennaPartialMetalArea                    0.324000 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.926457 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.324000 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.843917 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.641269 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.921689 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.401400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.957651 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.348000 LAYER metal1 ;
   AntennaGateArea                            0.363600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.173264 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.224000 LAYER metal1 ;
   AntennaDiffArea                            2.638350 LAYER metal1 ;
  END O

END OA222T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:40 CST 2007
#
#**********************************************************************




MACRO OA22P
  PIN A1
   AntennaPartialMetalArea                    0.352800 LAYER metal1 ;
   AntennaGateArea                            0.491400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.878711 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.353600 LAYER metal1 ;
   AntennaGateArea                            0.491400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.793243 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.412000 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837329 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.316000 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.741005 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.850400 LAYER metal1 ;
   AntennaDiffArea                            1.680100 LAYER metal1 ;
  END O

END OA22P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:44 CST 2007
#
#**********************************************************************




MACRO OA22S
  PIN A1
   AntennaPartialMetalArea                    0.296000 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.695513 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.340000 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.264961 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.185600 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.111107 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.192400 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.063032 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.774400 LAYER metal1 ;
   AntennaDiffArea                            0.583100 LAYER metal1 ;
  END O

END OA22S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:47 CST 2007
#
#**********************************************************************




MACRO OA22T
  PIN A1
   AntennaPartialMetalArea                    0.352800 LAYER metal1 ;
   AntennaGateArea                            0.491400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.878711 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.353600 LAYER metal1 ;
   AntennaGateArea                            0.491400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.793243 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.412000 LAYER metal1 ;
   AntennaGateArea                            0.496800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.850642 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.316000 LAYER metal1 ;
   AntennaGateArea                            0.496800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.757449 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.175600 LAYER metal1 ;
   AntennaDiffArea                            2.739500 LAYER metal1 ;
  END O

END OA22T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:51 CST 2007
#
#**********************************************************************




MACRO OAI112H
  PIN A1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.190000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.556400 LAYER metal1 ;
   AntennaDiffArea                            3.666600 LAYER metal1 ;
  END O

END OAI112H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:54 CST 2007
#
#**********************************************************************




MACRO OAI112HP
  PIN A1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.190000 LAYER metal1 ;
   AntennaGateArea                            2.194200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.751435 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            2.224800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.741101 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    2.847600 LAYER metal1 ;
   AntennaDiffArea                            7.293600 LAYER metal1 ;
  END O

END OAI112HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:48:57 CST 2007
#
#**********************************************************************




MACRO OAI112HS
  PIN A1
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.798012 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.821441 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.821441 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.798013 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.275200 LAYER metal1 ;
   AntennaDiffArea                            2.402200 LAYER metal1 ;
  END O

END OAI112HS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:01 CST 2007
#
#**********************************************************************




MACRO OAI112HT
  PIN A1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.190000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    4.335600 LAYER metal1 ;
   AntennaDiffArea                           10.999800 LAYER metal1 ;
  END O

END OAI112HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:04 CST 2007
#
#**********************************************************************




MACRO OAI12H
  PIN A1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.704296 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.863200 LAYER metal1 ;
   AntennaDiffArea                            3.250400 LAYER metal1 ;
  END O

END OAI12H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:07 CST 2007
#
#**********************************************************************




MACRO OAI12HP
  PIN A1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    2.902400 LAYER metal1 ;
   AntennaDiffArea                            5.928800 LAYER metal1 ;
  END O

END OAI12HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:10 CST 2007
#
#**********************************************************************




MACRO OAI12HS
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.665247 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.534600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.799849 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.774583 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.062400 LAYER metal1 ;
   AntennaDiffArea                            2.646100 LAYER metal1 ;
  END O

END OAI12HS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:12 CST 2007
#
#**********************************************************************




MACRO OAI12HT
  PIN A1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    3.970400 LAYER metal1 ;
   AntennaDiffArea                            8.750200 LAYER metal1 ;
  END O

END OAI12HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:15 CST 2007
#
#**********************************************************************




MACRO OAI13H
  PIN A1
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.797400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.773517 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.456200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.652383 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            1.456200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.959759 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.245200 LAYER metal1 ;
   AntennaGateArea                            1.330200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.995037 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    2.599200 LAYER metal1 ;
   AntennaDiffArea                            3.483600 LAYER metal1 ;
  END O

END OAI13H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:18 CST 2007
#
#**********************************************************************




MACRO OAI13HP
  PIN A1
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            1.594800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.806621 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            2.912400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.787529 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            2.912400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837453 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.298400 LAYER metal1 ;
   AntennaGateArea                            2.849400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.900676 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    4.431200 LAYER metal1 ;
   AntennaDiffArea                            5.356800 LAYER metal1 ;
  END O

END OAI13HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:22 CST 2007
#
#**********************************************************************




MACRO OAI13HS
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.453600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.865078 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.892800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.681451 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.892800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.681451 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.892800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.681452 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    2.037600 LAYER metal1 ;
   AntennaDiffArea                            2.223000 LAYER metal1 ;
  END O

END OAI13HS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:25 CST 2007
#
#**********************************************************************




MACRO OAI13HT
  PIN A1
   AntennaPartialMetalArea                    0.258400 LAYER metal1 ;
   AntennaGateArea                            2.392200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.757294 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            4.305600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.845365 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            4.305600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.925168 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.298400 LAYER metal1 ;
   AntennaGateArea                            4.242600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.979636 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    6.610400 LAYER metal1 ;
   AntennaDiffArea                            8.749400 LAYER metal1 ;
  END O

END OAI13HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:28 CST 2007
#
#**********************************************************************




MACRO OAI222H
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.235200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    2.456800 LAYER metal1 ;
   AntennaDiffArea                            4.368600 LAYER metal1 ;
  END O

END OAI222H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:31 CST 2007
#
#**********************************************************************




MACRO OAI222HP
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            2.158200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.763970 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    4.470400 LAYER metal1 ;
   AntennaDiffArea                            8.673600 LAYER metal1 ;
  END O

END OAI222HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:34 CST 2007
#
#**********************************************************************




MACRO OAI222HT
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.285000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.789041 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    6.570400 LAYER metal1 ;
   AntennaDiffArea                           13.042200 LAYER metal1 ;
  END O

END OAI222HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:37 CST 2007
#
#**********************************************************************




MACRO OAI222S
  PIN A1
   AntennaPartialMetalArea                    0.334000 LAYER metal1 ;
   AntennaGateArea                            0.584400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.599244 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.334000 LAYER metal1 ;
   AntennaGateArea                            0.584400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.754794 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.362000 LAYER metal1 ;
   AntennaGateArea                            0.585600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.620561 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.295500 LAYER metal1 ;
   AntennaGateArea                            0.579600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.710486 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.325600 LAYER metal1 ;
   AntennaGateArea                            0.601800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.807576 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.310000 LAYER metal1 ;
   AntennaGateArea                            0.604200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.632575 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.482400 LAYER metal1 ;
   AntennaDiffArea                            2.698150 LAYER metal1 ;
  END O

END OAI222S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:41 CST 2007
#
#**********************************************************************




MACRO OAI22H
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            1.067400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.661046 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.206000 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.626198 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.656400 LAYER metal1 ;
   AntennaDiffArea                            3.340800 LAYER metal1 ;
  END O

END OAI22H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:44 CST 2007
#
#**********************************************************************




MACRO OAI22HP
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.122200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.776929 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731629 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    3.043600 LAYER metal1 ;
   AntennaDiffArea                            6.673200 LAYER metal1 ;
  END O

END OAI22HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:47 CST 2007
#
#**********************************************************************




MACRO OAI22HT
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766774 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.249000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.797784 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    4.430800 LAYER metal1 ;
   AntennaDiffArea                           10.053600 LAYER metal1 ;
  END O

END OAI22HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:50 CST 2007
#
#**********************************************************************




MACRO OAI22S
  PIN A1
   AntennaPartialMetalArea                    0.312000 LAYER metal1 ;
   AntennaGateArea                            0.543600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.793229 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.339600 LAYER metal1 ;
   AntennaGateArea                            0.543600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.741356 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.315600 LAYER metal1 ;
   AntennaGateArea                            0.555600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.633545 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.210900 LAYER metal1 ;
   AntennaGateArea                            0.560400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.694152 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.120000 LAYER metal1 ;
   AntennaDiffArea                            1.780250 LAYER metal1 ;
  END O

END OAI22S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:52 CST 2007
#
#**********************************************************************




MACRO OR2
  PIN I1
   AntennaPartialMetalArea                    0.228000 LAYER metal1 ;
   AntennaGateArea                            0.291600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.367627 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.198509 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.068000 LAYER metal1 ;
   AntennaDiffArea                            1.124200 LAYER metal1 ;
  END O

END OR2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:55 CST 2007
#
#**********************************************************************




MACRO OR2B1
  PIN B1
   AntennaPartialMetalArea                    0.210800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.064392 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570464 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.548800 LAYER metal1 ;
   AntennaDiffArea                            1.448100 LAYER metal1 ;
  END O

END OR2B1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:49:58 CST 2007
#
#**********************************************************************




MACRO OR2B1P
  PIN B1
   AntennaPartialMetalArea                    0.252800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.678030 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.441000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.006351 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.998800 LAYER metal1 ;
   AntennaDiffArea                            1.396700 LAYER metal1 ;
  END O

END OR2B1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:01 CST 2007
#
#**********************************************************************




MACRO OR2B1S
  PIN B1
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.252000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.682536 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.292000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.952016 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.838000 LAYER metal1 ;
   AntennaDiffArea                            0.721000 LAYER metal1 ;
  END O

END OR2B1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:03 CST 2007
#
#**********************************************************************




MACRO OR2B1T
  PIN B1
   AntennaPartialMetalArea                    0.275900 LAYER metal1 ;
   AntennaGateArea                            0.176400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.651931 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.885600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.252711 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.372800 LAYER metal1 ;
   AntennaDiffArea                            2.724250 LAYER metal1 ;
  END O

END OR2B1T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:07 CST 2007
#
#**********************************************************************




MACRO OR2P
  PIN I1
   AntennaPartialMetalArea                    0.252800 LAYER metal1 ;
   AntennaGateArea                            0.453600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.938711 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.453600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.046295 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.814400 LAYER metal1 ;
   AntennaDiffArea                            1.462600 LAYER metal1 ;
  END O

END OR2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:09 CST 2007
#
#**********************************************************************




MACRO OR2S
  PIN I1
   AntennaPartialMetalArea                    0.359600 LAYER metal1 ;
   AntennaGateArea                            0.214200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.929035 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.286400 LAYER metal1 ;
   AntennaGateArea                            0.214200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.055092 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.642800 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END OR2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:12 CST 2007
#
#**********************************************************************




MACRO OR2T
  PIN I1
   AntennaPartialMetalArea                    0.224000 LAYER metal1 ;
   AntennaGateArea                            0.874800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.102881 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.224000 LAYER metal1 ;
   AntennaGateArea                            0.900000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.177331 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.596000 LAYER metal1 ;
   AntennaDiffArea                            2.780050 LAYER metal1 ;
  END O

END OR2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:15 CST 2007
#
#**********************************************************************




MACRO OR3
  PIN I1
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.415200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.034196 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.304000 LAYER metal1 ;
   AntennaGateArea                            0.415200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.973503 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.328000 LAYER metal1 ;
   AntennaGateArea                            0.415200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.973509 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.080100 LAYER metal1 ;
  END O

END OR3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:17 CST 2007
#
#**********************************************************************




MACRO OR3B1
  PIN B1
   AntennaPartialMetalArea                    0.292000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.021466 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.370000 LAYER metal1 ;
   AntennaGateArea                            0.367200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.100765 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.367200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.037033 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.563100 LAYER metal1 ;
  END O

END OR3B1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:20 CST 2007
#
#**********************************************************************




MACRO OR3B1P
  PIN B1
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.146469 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.370000 LAYER metal1 ;
   AntennaGateArea                            0.414000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.114490 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.414000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.976331 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.774400 LAYER metal1 ;
   AntennaDiffArea                            1.315000 LAYER metal1 ;
  END O

END OR3B1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:23 CST 2007
#
#**********************************************************************




MACRO OR3B1S
  PIN B1
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.952019 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.284000 LAYER metal1 ;
   AntennaGateArea                            0.259200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.559411 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.284000 LAYER metal1 ;
   AntennaGateArea                            0.259200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.559411 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.931200 LAYER metal1 ;
   AntennaDiffArea                            0.666400 LAYER metal1 ;
  END O

END OR3B1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:26 CST 2007
#
#**********************************************************************




MACRO OR3B1T
  PIN B1
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.146469 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.370000 LAYER metal1 ;
   AntennaGateArea                            0.432000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.068059 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.432000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.935652 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.122400 LAYER metal1 ;
   AntennaDiffArea                            2.643500 LAYER metal1 ;
  END O

END OR3B1T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:31 CST 2007
#
#**********************************************************************




MACRO OR3B2
  PIN B1
   AntennaPartialMetalArea                    0.188000 LAYER metal1 ;
   AntennaGateArea                            0.534600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.786385 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaGateArea                            0.534600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.850732 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.341800 LAYER metal1 ;
   AntennaGateArea                            0.190800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.553455 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.629200 LAYER metal1 ;
   AntennaDiffArea                            2.232900 LAYER metal1 ;
  END O

END OR3B2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:34 CST 2007
#
#**********************************************************************




MACRO OR3B2P
  PIN B1
   AntennaPartialMetalArea                    0.448800 LAYER metal1 ;
   AntennaGateArea                            0.190800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.392039 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.224000 LAYER metal1 ;
   AntennaGateArea                            0.190800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.483226 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.224800 LAYER metal1 ;
   AntennaGateArea                            0.438600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.987230 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.964000 LAYER metal1 ;
   AntennaDiffArea                            1.419500 LAYER metal1 ;
  END O

END OR3B2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:36 CST 2007
#
#**********************************************************************




MACRO OR3B2S
  PIN B1
   AntennaPartialMetalArea                    0.412000 LAYER metal1 ;
   AntennaGateArea                            0.261000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.638316 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.193800 LAYER metal1 ;
   AntennaGateArea                            0.261000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.888121 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.200000 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.280191 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.366400 LAYER metal1 ;
   AntennaDiffArea                            1.116500 LAYER metal1 ;
  END O

END OR3B2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:39 CST 2007
#
#**********************************************************************




MACRO OR3B2T
  PIN B1
   AntennaPartialMetalArea                    0.349600 LAYER metal1 ;
   AntennaGateArea                            0.190800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.392035 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.244000 LAYER metal1 ;
   AntennaGateArea                            0.190800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.367924 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.236000 LAYER metal1 ;
   AntennaGateArea                            0.432000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.043754 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.328000 LAYER metal1 ;
   AntennaDiffArea                            2.673000 LAYER metal1 ;
  END O

END OR3B2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:42 CST 2007
#
#**********************************************************************




MACRO OR3P
  PIN I1
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.415200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.022636 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.304000 LAYER metal1 ;
   AntennaGateArea                            0.415200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.973503 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.328000 LAYER metal1 ;
   AntennaGateArea                            0.415200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.973509 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.750400 LAYER metal1 ;
   AntennaDiffArea                            1.511200 LAYER metal1 ;
  END O

END OR3P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:45 CST 2007
#
#**********************************************************************




MACRO OR3S
  PIN I1
   AntennaPartialMetalArea                    0.232400 LAYER metal1 ;
   AntennaGateArea                            0.313200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.355682 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.304000 LAYER metal1 ;
   AntennaGateArea                            0.313200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.290544 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.328000 LAYER metal1 ;
   AntennaGateArea                            0.313200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.290546 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.665200 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END OR3S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:48 CST 2007
#
#**********************************************************************




MACRO OR3T
  PIN I1
   AntennaPartialMetalArea                    0.280000 LAYER metal1 ;
   AntennaGateArea                            0.444000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.946849 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.316000 LAYER metal1 ;
   AntennaGateArea                            0.444000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.910358 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.340000 LAYER metal1 ;
   AntennaGateArea                            0.444000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.910364 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.132800 LAYER metal1 ;
   AntennaDiffArea                            2.610900 LAYER metal1 ;
  END O

END OR3T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:50 CST 2007
#
#**********************************************************************




MACRO PDI
  PIN EB
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.622477 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    0.471200 LAYER metal1 ;
   AntennaDiffArea                            0.663000 LAYER metal1 ;
  END O

END PDI


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:53 CST 2007
#
#**********************************************************************




MACRO PDIX
  PIN EB
   AntennaPartialMetalArea                    0.194000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.699493 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    0.346000 LAYER metal1 ;
   AntennaDiffArea                            0.239200 LAYER metal1 ;
  END O

END PDIX


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:56 CST 2007
#
#**********************************************************************




MACRO PUI
  PIN E
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.804297 LAYER metal1 ; 
  END E

  PIN O
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaDiffArea                            0.801450 LAYER metal1 ;
  END O

END PUI


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:50:59 CST 2007
#
#**********************************************************************




MACRO QDBHN
  PIN CKB
   AntennaPartialMetalArea                    0.353200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.580812 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.288400 LAYER metal1 ;
   AntennaGateArea                            0.253800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.443652 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.600800 LAYER metal1 ;
   AntennaDiffArea                            1.406300 LAYER metal1 ;
  END Q

END QDBHN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:01 CST 2007
#
#**********************************************************************




MACRO QDBHS
  PIN CKB
   AntennaPartialMetalArea                    0.353200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.648992 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.288400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.396463 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.640000 LAYER metal1 ;
   AntennaDiffArea                            0.784000 LAYER metal1 ;
  END Q

END QDBHS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:04 CST 2007
#
#**********************************************************************




MACRO QDFFN
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.517678 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.285600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.890850 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.893200 LAYER metal1 ;
   AntennaDiffArea                            1.063300 LAYER metal1 ;
  END Q

END QDFFN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:07 CST 2007
#
#**********************************************************************




MACRO QDFFP
  PIN CK
   AntennaPartialMetalArea                    0.297600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.704542 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.959957 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.878400 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END Q

END QDFFP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:10 CST 2007
#
#**********************************************************************




MACRO QDFFRBN
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.977273 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.778958 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.628000 LAYER metal1 ;
   AntennaDiffArea                            1.218700 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.193997 LAYER metal1 ; 
  END RB

END QDFFRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:13 CST 2007
#
#**********************************************************************




MACRO QDFFRBP
  PIN CK
   AntennaPartialMetalArea                    0.297600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.579542 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.233600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839421 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.666400 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.289600 LAYER metal1 ;
   AntennaGateArea                            0.898200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.763977 LAYER metal1 ; 
  END RB

END QDFFRBP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:16 CST 2007
#
#**********************************************************************




MACRO QDFFRBS
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.977273 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.778958 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.810000 LAYER metal1 ;
   AntennaDiffArea                            0.769300 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.233600 LAYER metal1 ;
   AntennaGateArea                            0.608400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.357332 LAYER metal1 ; 
  END RB

END QDFFRBS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:18 CST 2007
#
#**********************************************************************




MACRO QDFFRBT
  PIN CK
   AntennaPartialMetalArea                    0.249600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.472222 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    1.616000 LAYER metal1 ;
   AntennaDiffArea                            2.917300 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.898200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.791361 LAYER metal1 ; 
  END RB

END QDFFRBT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:21 CST 2007
#
#**********************************************************************




MACRO QDFFRSBN
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.392673 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.612000 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.459600 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.212610 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    1.568400 LAYER metal1 ;
   AntennaGateArea                            0.493200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.503791 LAYER metal1 ; 
  END SB

END QDFFRSBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:24 CST 2007
#
#**********************************************************************




MACRO QDFFS
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.517678 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.285600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.890850 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.893200 LAYER metal1 ;
   AntennaDiffArea                            0.626500 LAYER metal1 ;
  END Q

END QDFFS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:26 CST 2007
#
#**********************************************************************




MACRO QDFZN
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.494948 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.893200 LAYER metal1 ;
   AntennaDiffArea                            1.063300 LAYER metal1 ;
  END Q

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277069 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END QDFZN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:29 CST 2007
#
#**********************************************************************




MACRO QDFZP
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.494948 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.844800 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END Q

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277069 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END QDFZP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:32 CST 2007
#
#**********************************************************************




MACRO QDFZRBN
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.506313 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.779200 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.193997 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227899 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END QDFZRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:35 CST 2007
#
#**********************************************************************




MACRO QDFZRBP
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.494953 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.896000 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.898200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.787128 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227899 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END QDFZRBP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:38 CST 2007
#
#**********************************************************************




MACRO QDFZRBS
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.506313 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.841600 LAYER metal1 ;
   AntennaDiffArea                            0.769300 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.608400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.378043 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227899 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END QDFZRBS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:40 CST 2007
#
#**********************************************************************




MACRO QDFZRBT
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.494953 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    1.590400 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.898200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.787128 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227899 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END QDFZRBT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:43 CST 2007
#
#**********************************************************************




MACRO QDFZRSBN
  PIN CK
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.506313 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.612000 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.455600 LAYER metal1 ;
   AntennaGateArea                            0.666000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.212616 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    1.566000 LAYER metal1 ;
   AntennaGateArea                            0.493200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.486108 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.227899 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END QDFZRSBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:47 CST 2007
#
#**********************************************************************




MACRO QDFZS
  PIN CK
   AntennaPartialMetalArea                    0.225600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.494948 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.273600 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.753048 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.893200 LAYER metal1 ;
   AntennaDiffArea                            0.626500 LAYER metal1 ;
  END Q

  PIN SEL
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.423000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277069 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.869950 LAYER metal1 ; 
  END TD

END QDFZS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:49 CST 2007
#
#**********************************************************************




MACRO QDLHN
  PIN CK
   AntennaPartialMetalArea                    0.353200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.717172 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.288400 LAYER metal1 ;
   AntennaGateArea                            0.253800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.443652 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.600800 LAYER metal1 ;
   AntennaDiffArea                            1.406300 LAYER metal1 ;
  END Q

END QDLHN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:52 CST 2007
#
#**********************************************************************




MACRO QDLHP
  PIN CK
   AntennaPartialMetalArea                    0.353200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.717172 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.480400 LAYER metal1 ;
   AntennaGateArea                            0.271800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.348054 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.580000 LAYER metal1 ;
   AntennaDiffArea                            1.641600 LAYER metal1 ;
  END Q

END QDLHP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:55 CST 2007
#
#**********************************************************************




MACRO QDLHRBN
  PIN CK
   AntennaPartialMetalArea                    0.494200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.790401 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.306800 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.525924 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.709600 LAYER metal1 ;
   AntennaDiffArea                            1.411200 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.323200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.230859 LAYER metal1 ; 
  END RB

END QDLHRBN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:51:58 CST 2007
#
#**********************************************************************




MACRO QDLHRBP
  PIN CK
   AntennaPartialMetalArea                    0.494200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.790401 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.306800 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.204674 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.647400 LAYER metal1 ;
   AntennaDiffArea                            1.647000 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.323200 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.166081 LAYER metal1 ; 
  END RB

END QDLHRBP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:00 CST 2007
#
#**********************************************************************




MACRO QDLHRBS
  PIN CK
   AntennaPartialMetalArea                    0.494200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.790401 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.306800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.601011 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.709600 LAYER metal1 ;
   AntennaDiffArea                            0.793800 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.323200 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.350949 LAYER metal1 ; 
  END RB

END QDLHRBS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:03 CST 2007
#
#**********************************************************************




MACRO QDLHS
  PIN CK
   AntennaPartialMetalArea                    0.353200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.785352 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.288400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.396463 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.640000 LAYER metal1 ;
   AntennaDiffArea                            0.784000 LAYER metal1 ;
  END Q

END QDLHS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:06 CST 2007
#
#**********************************************************************




MACRO QDLHSN
  PIN CK
   AntennaPartialMetalArea                    0.487600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.251267 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.282800 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.556389 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.435700 LAYER metal1 ;
  END Q

  PIN S
   AntennaPartialMetalArea                    0.304800 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.953568 LAYER metal1 ; 
  END S

END QDLHSN


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:09 CST 2007
#
#**********************************************************************




MACRO RAM2
  PIN D
   AntennaPartialMetalArea                    0.204000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.529041 LAYER metal1 ; 
  END D

  PIN QB
   AntennaPartialMetalArea                    0.826000 LAYER metal1 ;
   AntennaDiffArea                            1.156400 LAYER metal1 ;
  END QB

  PIN QBZ
   AntennaPartialMetalArea                    1.981200 LAYER metal1 ;
   AntennaDiffArea                            2.288650 LAYER metal1 ;
  END QBZ

  PIN RD
   AntennaPartialMetalArea                    0.233600 LAYER metal1 ;
   AntennaGateArea                            0.651600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.321978 LAYER metal1 ; 
  END RD

  PIN W
   AntennaPartialMetalArea                    1.350400 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.580804 LAYER metal1 ; 
  END W

END RAM2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:14 CST 2007
#
#**********************************************************************




MACRO RAM2S
  PIN D
   AntennaPartialMetalArea                    0.221200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.237375 LAYER metal1 ; 
  END D

  PIN QB
   AntennaPartialMetalArea                    0.564400 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END QB

  PIN QBZ
   AntennaPartialMetalArea                    1.013600 LAYER metal1 ;
   AntennaDiffArea                            1.504300 LAYER metal1 ;
  END QBZ

  PIN RD
   AntennaPartialMetalArea                    0.348000 LAYER metal1 ;
   AntennaGateArea                            0.392400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.654940 LAYER metal1 ; 
  END RD

  PIN W
   AntennaPartialMetalArea                    1.328400 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.785358 LAYER metal1 ; 
  END W

END RAM2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:17 CST 2007
#
#**********************************************************************




MACRO RAM3
  PIN D
   AntennaPartialMetalArea                    0.198400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.324495 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.651600 LAYER metal1 ;
   AntennaDiffArea                            1.251250 LAYER metal1 ;
  END Q

  PIN QZ
   AntennaPartialMetalArea                    1.804400 LAYER metal1 ;
   AntennaDiffArea                            2.486650 LAYER metal1 ;
  END QZ

  PIN RD
   AntennaPartialMetalArea                    0.213600 LAYER metal1 ;
   AntennaGateArea                            0.651600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.396562 LAYER metal1 ; 
  END RD

  PIN W
   AntennaPartialMetalArea                    1.318800 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.050521 LAYER metal1 ; 
  END W

END RAM3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:20 CST 2007
#
#**********************************************************************




MACRO RAM3S
  PIN D
   AntennaPartialMetalArea                    0.192800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.324498 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.657600 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END Q

  PIN QZ
   AntennaPartialMetalArea                    0.971600 LAYER metal1 ;
   AntennaDiffArea                            1.504300 LAYER metal1 ;
  END QZ

  PIN RD
   AntennaPartialMetalArea                    0.348000 LAYER metal1 ;
   AntennaGateArea                            0.392400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.807340 LAYER metal1 ; 
  END RD

  PIN W
   AntennaPartialMetalArea                    1.335600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.050491 LAYER metal1 ; 
  END W

END RAM3S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:23 CST 2007
#
#**********************************************************************




MACRO RAM5
  PIN D
   AntennaPartialMetalArea                    0.257200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.324493 LAYER metal1 ; 
  END D

  PIN QZ0
   AntennaPartialMetalArea                    1.501600 LAYER metal1 ;
   AntennaDiffArea                            2.494600 LAYER metal1 ;
  END QZ0

  PIN QZ1
   AntennaPartialMetalArea                    1.769600 LAYER metal1 ;
   AntennaDiffArea                            2.353800 LAYER metal1 ;
  END QZ1

  PIN RD0
   AntennaPartialMetalArea                    0.229600 LAYER metal1 ;
   AntennaGateArea                            0.634800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.433521 LAYER metal1 ; 
  END RD0

  PIN RD1
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.634800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.450535 LAYER metal1 ; 
  END RD1

  PIN W
   AntennaPartialMetalArea                    1.239600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.050521 LAYER metal1 ; 
  END W

END RAM5


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:26 CST 2007
#
#**********************************************************************




MACRO RAM5S
  PIN D
   AntennaPartialMetalArea                    0.257200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.324493 LAYER metal1 ; 
  END D

  PIN QZ0
   AntennaPartialMetalArea                    0.597600 LAYER metal1 ;
   AntennaDiffArea                            1.312400 LAYER metal1 ;
  END QZ0

  PIN QZ1
   AntennaPartialMetalArea                    0.883600 LAYER metal1 ;
   AntennaDiffArea                            1.260600 LAYER metal1 ;
  END QZ1

  PIN RD0
   AntennaPartialMetalArea                    0.241600 LAYER metal1 ;
   AntennaGateArea                            0.392400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.103462 LAYER metal1 ; 
  END RD0

  PIN RD1
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.392400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.103464 LAYER metal1 ; 
  END RD1

  PIN W
   AntennaPartialMetalArea                    1.225600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.050513 LAYER metal1 ; 
  END W

END RAM5S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:28 CST 2007
#
#**********************************************************************




MACRO TIE0
  PIN O
   AntennaPartialMetalArea                    0.314400 LAYER metal1 ;
   AntennaDiffArea                            0.493000 LAYER metal1 ;
  END O

END TIE0


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:31 CST 2007
#
#**********************************************************************




MACRO TIE1
  PIN O
   AntennaPartialMetalArea                    0.314400 LAYER metal1 ;
   AntennaDiffArea                            0.586000 LAYER metal1 ;
  END O

END TIE1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:34 CST 2007
#
#**********************************************************************




MACRO XNR2H
  PIN I1
   AntennaPartialMetalArea                    0.275200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.789849 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.347200 LAYER metal1 ;
   AntennaGateArea                            1.602000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.083641 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.881600 LAYER metal1 ;
   AntennaDiffArea                            4.322200 LAYER metal1 ;
  END O

END XNR2H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:36 CST 2007
#
#**********************************************************************




MACRO XNR2HP
  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785943 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.006740 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    3.263200 LAYER metal1 ;
   AntennaDiffArea                            7.983200 LAYER metal1 ;
  END O

END XNR2HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:39 CST 2007
#
#**********************************************************************




MACRO XNR2HS
  PIN I1
   AntennaPartialMetalArea                    0.235200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.631165 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.303600 LAYER metal1 ;
   AntennaGateArea                            0.838800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.243204 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.916000 LAYER metal1 ;
   AntennaDiffArea                            1.706400 LAYER metal1 ;
  END O

END XNR2HS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:42 CST 2007
#
#**********************************************************************




MACRO XNR2HT
  PIN I1
   AntennaPartialMetalArea                    0.232400 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.813632 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.480400 LAYER metal1 ;
   AntennaGateArea                            4.806000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.936242 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    4.636000 LAYER metal1 ;
   AntennaDiffArea                           11.210500 LAYER metal1 ;
  END O

END XNR2HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:44 CST 2007
#
#**********************************************************************




MACRO XNR3
  PIN I1
   AntennaPartialMetalArea                    0.287600 LAYER metal1 ;
   AntennaGateArea                            0.463800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.079775 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.248000 LAYER metal1 ;
   AntennaGateArea                            0.484200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.269515 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.614198 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.498600 LAYER metal1 ;
  END O

END XNR3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:47 CST 2007
#
#**********************************************************************




MACRO XNR3P
  PIN I1
   AntennaPartialMetalArea                    0.287600 LAYER metal1 ;
   AntennaGateArea                            0.463800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.079775 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.248000 LAYER metal1 ;
   AntennaGateArea                            0.484200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.269515 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.229600 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.503088 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.697600 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END O

END XNR3P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:50 CST 2007
#
#**********************************************************************




MACRO XNR3S
  PIN I1
   AntennaPartialMetalArea                    0.243600 LAYER metal1 ;
   AntennaGateArea                            0.192600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.934582 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.248000 LAYER metal1 ;
   AntennaGateArea                            0.484200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.310825 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.391978 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.914400 LAYER metal1 ;
   AntennaDiffArea                            0.666400 LAYER metal1 ;
  END O

END XNR3S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:52 CST 2007
#
#**********************************************************************




MACRO XNR3T
  PIN I1
   AntennaPartialMetalArea                    0.287600 LAYER metal1 ;
   AntennaGateArea                            0.463800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.079775 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.248000 LAYER metal1 ;
   AntennaGateArea                            0.484200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.269515 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.261600 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.425313 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.428800 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END O

END XNR3T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:55 CST 2007
#
#**********************************************************************




MACRO XNR4
  PIN I1
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.422400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287880 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.806000 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.266660 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.859851 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    1.271600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                         10.669811 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.750400 LAYER metal1 ;
   AntennaDiffArea                            1.340400 LAYER metal1 ;
  END O

END XNR4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:52:58 CST 2007
#
#**********************************************************************




MACRO XNR4P
  PIN I1
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.422400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287880 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.873200 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.906108 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.439391 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    1.293400 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                         10.669798 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.878400 LAYER metal1 ;
   AntennaDiffArea                            1.464900 LAYER metal1 ;
  END O

END XNR4P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:01 CST 2007
#
#**********************************************************************




MACRO XNR4S
  PIN I1
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.422400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287880 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.786800 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.160632 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.439391 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    1.293400 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                         10.669798 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.750400 LAYER metal1 ;
   AntennaDiffArea                            0.769300 LAYER metal1 ;
  END O

END XNR4S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:05 CST 2007
#
#**********************************************************************




MACRO XNR4T
  PIN I1
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.422400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287880 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.782000 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.160600 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.439391 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    1.293400 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                         10.669798 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    1.221600 LAYER metal1 ;
   AntennaDiffArea                            2.683200 LAYER metal1 ;
  END O

END XNR4T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:08 CST 2007
#
#**********************************************************************




MACRO XOR2H
  PIN I1
   AntennaPartialMetalArea                    0.275200 LAYER metal1 ;
   AntennaGateArea                            1.126800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.735535 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.347200 LAYER metal1 ;
   AntennaGateArea                            1.602000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.056181 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.922400 LAYER metal1 ;
   AntennaDiffArea                            4.364100 LAYER metal1 ;
  END O

END XOR2H


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:11 CST 2007
#
#**********************************************************************




MACRO XOR2HP
  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            2.253600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.731630 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            3.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.006740 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    3.263200 LAYER metal1 ;
   AntennaDiffArea                            8.051400 LAYER metal1 ;
  END O

END XOR2HP


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:14 CST 2007
#
#**********************************************************************




MACRO XOR2HS
  PIN I1
   AntennaPartialMetalArea                    0.235200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.631165 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.239200 LAYER metal1 ;
   AntennaGateArea                            0.833400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.257743 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.902400 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END O

END XOR2HS


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:16 CST 2007
#
#**********************************************************************




MACRO XOR2HT
  PIN I1
   AntennaPartialMetalArea                    0.246400 LAYER metal1 ;
   AntennaGateArea                            3.380400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.766773 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.494400 LAYER metal1 ;
   AntennaGateArea                            4.806000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932589 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    4.636000 LAYER metal1 ;
   AntennaDiffArea                           11.030500 LAYER metal1 ;
  END O

END XOR2HT


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:19 CST 2007
#
#**********************************************************************




MACRO XOR3
  PIN I1
   AntennaPartialMetalArea                    0.255600 LAYER metal1 ;
   AntennaGateArea                            0.443400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.017595 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.248000 LAYER metal1 ;
   AntennaGateArea                            0.484200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.336435 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.794758 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.577800 LAYER metal1 ;
  END O

END XOR3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:22 CST 2007
#
#**********************************************************************




MACRO XOR3P
  PIN I1
   AntennaPartialMetalArea                    0.255600 LAYER metal1 ;
   AntennaGateArea                            0.443400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.017595 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.248000 LAYER metal1 ;
   AntennaGateArea                            0.484200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.336435 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.741358 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.697600 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END O

END XOR3P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:25 CST 2007
#
#**********************************************************************




MACRO XOR3S
  PIN I1
   AntennaPartialMetalArea                    0.255600 LAYER metal1 ;
   AntennaGateArea                            0.194400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.737655 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.248000 LAYER metal1 ;
   AntennaGateArea                            0.484200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.336435 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.201600 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.683638 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.749200 LAYER metal1 ;
   AntennaDiffArea                            0.666400 LAYER metal1 ;
  END O

END XOR3S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:30 CST 2007
#
#**********************************************************************




MACRO XOR3T
  PIN I1
   AntennaPartialMetalArea                    0.247600 LAYER metal1 ;
   AntennaGateArea                            0.443400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.017588 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.248000 LAYER metal1 ;
   AntennaGateArea                            0.484200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.328995 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.229600 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.669758 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.428800 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END O

END XOR3T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:32 CST 2007
#
#**********************************************************************




MACRO XOR4
  PIN I1
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.422400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287880 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.786800 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.215132 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.439391 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    1.305100 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                         10.669866 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.766400 LAYER metal1 ;
   AntennaDiffArea                            1.340400 LAYER metal1 ;
  END O

END XOR4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:35 CST 2007
#
#**********************************************************************




MACRO XOR4P
  PIN I1
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.422400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287880 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.839600 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.942384 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.439391 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    1.305100 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                         10.669866 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.858400 LAYER metal1 ;
   AntennaDiffArea                            1.502700 LAYER metal1 ;
  END O

END XOR4P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:39 CST 2007
#
#**********************************************************************




MACRO XOR4S
  PIN I1
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.422400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287880 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.760400 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.215106 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.439391 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    1.305100 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                         10.669866 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.766400 LAYER metal1 ;
   AntennaDiffArea                            0.769300 LAYER metal1 ;
  END O

END XOR4S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:53:44 CST 2007
#
#**********************************************************************




MACRO XOR4T
  PIN I1
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.422400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287880 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    1.782000 LAYER metal1 ;
   AntennaGateArea                            0.356400 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.215200 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.268000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.439391 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    1.321600 LAYER metal1 ;
   AntennaGateArea                            0.316800 LAYER metal1 ;
   AntennaMaxAreaCAR                         10.669783 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    1.204400 LAYER metal1 ;
   AntennaDiffArea                            2.695500 LAYER metal1 ;
  END O

END XOR4T



END LIBRARY
