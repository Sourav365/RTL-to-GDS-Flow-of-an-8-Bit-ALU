//////////////////////////////////////////////////////////////////////
// (C) Copyright 1993-2003 Faraday Technology Corp. All Rights Reserved.
// 
// FTC Verilog Simulation Library
//   Cell Library            : fsa0m_a
//   Library Release Version : 2009Q2v2.0
//   Date                    : Tue May  5 13:35:36 CST 2009 
//////////////////////////////////////////////////////////////////////
//
//   Note : This library uses delayed signals to support negative
//          timing checks.
//          Please add command-line options
//             "+neg_tchk" and "+nowarnNTCDSN" when runnning simulation with Verilog-XL
//             "+neg_tchk" when runnning simulation with NC-verilog
//          to support negative timing checks.
//
//////////////////////////////////////////////////////////////////////

`timescale 10ps / 1ps

//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN2(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
ic5NCSQ:5DT^<iYa3NmfM9nR^_K;n5EEi]G>SK:R<_J`PIDCoAL?n_LLgQAa8[U9
1Ep;alJJa3I^nOD0JXY\MegVf>WRTR;>bG4DYDoTFN7JIV@\H@>J?Mi^o@APIFVn
m`Yqnkkf5eBhJa\CN3K^igkBHkP=D:ViRG4l7A`L3@6BM8E_fe6b\hlCgV9q:j0R
\Mq7c_l2iUYN38k5GHj2i7:nQS@U4>ccbmqUlL\CHjpbN@9=@qIZd\PSdUYA1XC7
cBPNkdM79lVQjU97<SVhCc`>T[:oUNicNdd6X0X8Di6\0@B\\>Ie^M[8h:FU^Y:]
KPmmXqmN1>3ESl^b7o0nR87hiEl_[?c=YKICCCcMSj]1^4^7?HQ2Im`\iHq6BN<=
OO>C=b73`cj;lmPWI@e?RjC7hHKZ4aYjGQL:2m5<W[kC7X]<3WIH27]TKIA6O]^1
gd0Hj[7e3FfiPFpXeKLDhD$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN2B1(O, I1, B1);
   output O;
   input I1, B1;

//Function Block
`protected
Xj954SQV5DT^<IUKhBcB:KJ?TA\oKa<me\8Sf`I;nn6AkWDaV9CmdJ@?HQAU8[[9
IEpF0ClGX^b1H^m9M1U;d^^ilj^M15O4WjQ0;]932oMbSjKeWANOafp`O3f?Vo]7
jk[gF9QOGJk9<mc[DepUj@VFbq077\PL^c[5<mhkkYUkYOb:nlM?>qN8IbkJ@dPa
<`=8GT4YPS522JIDXD>m?qdfBana@qS76^O1poDo?6L[HVDE_H8fTdncNLD=`Yem
@\6W0<RheWSDH:3]j=4J2Zck3\cR23\f\CYdgo8iO\VAonIX;V761Tilq2EJaAnk
ce0f>XRRU=g`j][i552^]gfDZb4;co8>SYQl1E_oaHc7696igKSG^PbOa2n3gj\G
bK0NdgJXHh1fq\P@KYU6$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN2B1P(O, I1, B1);
   output O;
   input I1, B1;

//Function Block
`protected
gnO39SQH5DT^<::hU^aj<EgdSWjIH5HC^Mo^7:3Qa6iTR]_>OoIDH>>3RbMB70Fa
pBKDeO<AMHJ>4RDFQEbX`S_emTcUmY1=nSh43h9:6[Q7MQNqYS>_ml\Z5kKMBVkh
:C[^=>YMJRI?EJOLB3j@TQ5N5PX[f@jqMXLI>bp4FQDOm@FW45^cC\]?h=k2<6[g
@;pd8GCGN4ZFh2jW3edZBHG`o^>QjIa@moq6jnCEcEqk@`Na1pON73J:SV>N;GGR
MT[X9D?@ojbAEO_I9E2:I\fK>aRD:`6Qc43lT?6EIlBER`J:B3O4bnk]7JSY<a6K
C];=2p`nRXC8ZRZDR]aK28Tl3OjC3e@E_M@fiQFT]OUPcIHdB@maRdHQm\hhj__k
fVFk=lPL`jlXIQUP\2:\ll`:lm5FM9bCKpbE6i`H079BR?Y`la5XREP[k2>N[mdB
?9]m63g@Y5hC1@=HIXoo[LI<pco_QCc@$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN2B1S(O, I1, B1);
   output O;
   input I1, B1;

//Function Block
`protected
Nfi@;SQd5DT^<?e1fjoX8nIEdh>=F?m9[ROJWNc:LVNmdhC29ja_NZXmRbMB7P[G
pZ2VSH@fJK?OQR048BMg1QbPiUN7cig?<0X5fQFWoo6]5?1Y^@PLE4?b<N@pHJUl
>V<727Y9F3np?LA\ngqQIe?fboE1ZF>NIiD72@7?JgQoTGq4WGeFkJUlJ8Y1aLDj
M_9AS@B`\IJ1VCpg];DKG@p_<l@EXpT?ZZUfGYDDSUJoeMQ;hF17EH5U7AZNU:9X
E=g<C86nCRY>H8ZST\cjEZ?m=>CaQ<TP3iFVBYUa\28k\60h4q;0\amF0lEZATdi
MO9j:UeUcMD4^0Tc\55NhhMnZ11bmNRT4AU5Mcnn><[YUXkh_j;d[>EKo9Pb02>h
FefERpV0IbRST$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN2B1T(O, I1, B1);
   output O;
   input I1, B1;

//Function Block
`protected
PBG4gSQd5DT^<kahdA^[4S<k14j[fQFcV<OkPVB[ceP2W1I0H`UibG4HX<coMKPq
8KSYV7?dJQo?IaMVEi6o\bZ`A=l0OblH9h;WnNOCCQ:[8;Zc;]g=_c>1_OlR01Nk
=nCf5WpiGMI?i39gW\Q]]J\PL2Qn:o<M`_BW`4<93_5I6HK=mOFN3Vq5i1jBGqI>
c5ajPm[Ek3bV7k[S?eQ3M[bQ[pfE?nK^ee]5FI1VkdJe_Do4?ZLj?<Xf0qT_XWiV
:p2RFR=g2E>bWK2n>Xk1QnS<VU4dbUDGXaT0`>@KYqRQN]77pBWF^j0Z0G@lCKfA
Z2GG:h0o`?WBVKAgBX:QGZ1g[WXXUWD2H`2BGK[G=i8k;Mf3YB8jnVBhWCKlZ7FS
7bS3piTDl?NhAi`]\:@AXbDZc\VL?V;7lb:d;]k9:i9WW89K^lniYFjMbXJ<6S\b
7:SF]1RN]^A3\Pc`DT8i=cXd7RZ4q:b]?^B2$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN2P(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
>\3HlSQd5DT^<<mhMnX<TfKoeS\1Ic?QeL3aW>;N4X>WkYE`9Kd7mG4kX<co7EPq
\1Fg?5TJ?g8FZV[Y=0=NP_2;07a79;37\\S>eJD29BU4]e@>7b\ARU7IqmMU`ooI
:3IZ]>T4g4VTc4cGV=NXGFcFHq9[9E``p3SO>=3W<1UL2gWEJgIb4^:o0cW>\\A2
pc9<VTc3qJ2jDF<jdPBk`:1V9XgII<Mh<=DU]@8hSOnGdCBmDRafN@T]5fXKOmM>
0AA]<8?`Yq>@WHQmq?1c<]6_4B1cFLEBmM\A>LAK4SB2nNoYMO_YADOo;eciX_8K
H?0W?C>T1^TgLO;_O?mV]H[OB5@aDU?IXXL^qdKA<o0bPEblA_F<[f@3j:_P[kfE
RI1;Bj`<8AJHm@7aUb=`]mQDbYWjGC>IcZonAd?WMJa@4<Qe7D=g]PeRqJRkfPO9
$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN2S(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
?:;YHSQH5DT^<C_:X;me0AnCmX2?0gIUI11E0k:lAOI0HEh?RQJUMjo4GBG>kop:
@\H:2[^i2M5;]oOhJ[b7?djZQW[p<n1fUP=Ke?lPl8j^E=JSCY[17ZmFOFX0RNl^
H4bmhNDKmAmpWQLM``pR]EP]97M;e0TYLLN3kY4>YZV?O_K^6kqNF<LjLKpD9UG]
OqbZ;8LCMd5H:lSH]Dh_96F4Ka\cGBT^[^^i5]=MVj57VIU?k]ZM?EE_YORBOcBf
:jb1X<ld3LenmG>bG4b:3pF][QaDkQW=:i2P6nXgMghX=<B9^=IAUj;e1bh;_]ZA
Ah5\GK0Cg6\75McfY=0CO:FIcF2JCllJD<<TTi60aq@8HFCSC]:][j^80X[cl7d9
?@^<2[WJ7Xcegp`o8OoZ:$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN2T(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
Xb_DmSQ:5DT^<n@Y?<fFW:5;PLbgio02]o=jUQK`]knL>CLIMWBG0f?M_o7_q5FK
TCM0Um<1f<JpUgCEDX_Ok]@C21<>3@^nm5a7jWnf?m=ofGL<RcM]fRJW]1\l<3NP
<bk7`f3pK<9i3`q98ijYGhR\V\ge8Q2FA>c5gI_cOQUgH3pc\_=MEBqWHl:T0AE4
I3ZiHbp2ll0?Oq77PW9Ib_<JK9o7kV]EP]5GWL]lm^jL]OOlhonFlW]TA`b>0hQP
ZB@<hmPXj[Cn727_=onHY=D:6fgeML24]pX4COJgW>eMVc5=gfeY9CnUND[LRLi0
FKkjVMjM9JK;HZW:cG2mT:HS356Lk;??_9XJedlY:\YXB7`IAk:4iqeJkFERQ$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
U?_^`SQ:5DT^<nY:[@DRglV4m8ImCb`7N?B2ehImo2NUHV9LF6M]0f?M_f7nq[@I
[K5^V6HT`ED0Plf1[_7Dm\oQP4S`TLb_WLU8CGOS@5[hG[ClQ`2p3S^fKXEgl6f>
RL>3HPDhZVk@SL7H\mRScHSpDiC4Fbq;V_>bD50HZNiEE64KooIO3=Ah^Q=df\:b
]J>q@`7H`_eqNa7\[Gq\]?cH7J_C;2WD1C]C5jEmd1CFj<I@4<53Fb90mUY[RD@]
=05:NZn]nTm2HLZ4VQM\[U^LVe1o[\X?bhNaMjpElo0LMIOb\2An:`g3J`LP3UGl
8LIBK<llLR6hcF7ZUJD]<n@an]Hl<A@m7XK5j4HEKcoY5c>a``_AGSi5^=p0?OR5
OF4BjeAdULfMU>8jnaR;G>W\[hQXC@_GAeXK_DBn;W?;Z[CNifIEYP[m@590d=:_
S];UbkD:98=\VEqiYl;BnA$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3B1(O, I1, I2, B1);
   output O;
   input I1, I2, B1;

//Function Block
`protected
o?l=?SQV5DT^<K4iE>i3]LMnC@_9hod@n=ec6a0\JZC4W]@6=BfoCZJ9Gkmp85A_
REVT9dW\Kkq0JTZMfahH>6c<S[7bJ@YB046P<W5TLT;[7GKNl7KG3UAT?KV>LjqX
85XXjpg<;\B;<62GIhBcRVXjj=[J1K8=HqBC=ncDTGO`OkS2KOCmdJgbj2nWQ3>5
NkB[FbqGfd7W]YpSReD?OpgF@WIVam=CGN;BHbF9DakGP:>b_V90=S`mTWY^W38;
Z\8GT<N6<XiccioHmmN;Dig8AUldMA6`RnQ4TJS;hqGUUimhXR3h:a0E5l<B?<>T
KhFoYF2N`lPdM5=QS3F@E@caoM9:ne]@XJFPF>kFm4GM0k@bBnN\HOUQH02BWpb\
_<gciP8dHZFLB:CML:S=o11[omNd04]?XRNTmOLg>1F>8VjGDE3nZIiD0NS3]?pg
ibPkW?B1S3aDGOE[lFEnVA@c@B[liPUWQ\I:fMWO6^daV<mBgT[3UJoTaBP7k\m:
ATiOhWbCn4;_CNmAh;Jl;nq8cA4V`:$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3B1P(O, I1, I2, B1);
   output O;
   input I1, I2, B1;

//Function Block
`protected
<1K3ZSQV5DT^<cjaCH`>nBXLi14j4BdaE@P1f[HD=\FK5RY1:@fZCZJ96^=pl[f2
B6MJKg<\ORfVmXXRAdMq]2B1G`I:Xo?>jB_lpFNUR7?qC^VDaGXdX?0Yl<V\5^_7
9X;c8UhqJC[:jO<[QoNO_>H0_<CK0ISaN7b2MPc2b<23q2L33E:3pOO0b\Mq8H=e
3d0`[DLdQ_RX7GYV=KGE9`Uo@h;HX3[1RR_`7Cq\YT<iRDg1A2\ZkDYSYM[fb8Lg
ZO?SLaO;2PkZNn]e=:Ri7RSBTMadi?D35OOE?0<NPPUcgGU[@n5V@9hPY`^dZ@>G
m[pg6?o86A9DQ:PW=Goe08HGKZ<9`@A`7J9aYdMbDHCHQIccF1GGdC:5=[<2UVIG
AEN[`6>ihIG9?FBjDAWO5CMX39DT;>p_5lF[E9P^`YZWWi[6fKIjTBL[6XI7V_Nm
899YOML6Mh2EHIS]geXbgm:n]klmHmjY_`nAXmQ@S`e2@[\5f]mKi4FBYdph8fGj
H1$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3B1S(O, I1, I2, B1);
   output O;
   input I1, I2, B1;

//Function Block
`protected
RK3FXSQ:5DT^<OobHG\jSnFSOj>`Y8G>K5Ua?LZ1b0UC0FPbUlQNjj9EAYqFEWhi
>olmPYiE>l4m:Dfbho>BUDF:V78_FY3fCXg]bq7e\jSN4WYSZilGb5CZL2gk7]@c
FGi8iMRRml81`41m\MDd995C?RPU\GMDI_9;CVVeS;p56eb^Xp5S_QJW1[Hd3[X4
H<i`UPkVS`:Ddq]fPX1=GYYEdV_^QUOeGkK]79k;6VC;R5l4`Mpl:h?hZ6q5DgS\
lqPJ=>2?4NXZZECQE<aAl0E]T`;EQlW6jNo6SI2R3Y@D3[nA39oWcW>;5I^ASiBE
5cPPBfhNo2fg_]0b1JV`^pbPoaRKj`@j`I_Y5CZcJXL@73L:17]Sf7cSS>`@DaKY
a2:Dhh6G0`Q9lT?X<ClLEPb9]C@`3:e046\l=ih?>q[47:Mo>Q1UB5Cga4m>k@9G
Y`Kf6H_Z3>2oZd^jeSV4Ih34JUMf1gfJXZL6FFj\;S[?eUNOO6FKX8TigZF`1q0i
UUQEm$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3B1T(O, I1, I2, B1);
   output O;
   input I1, I2, B1;

//Function Block
`protected
BkE>@SQV5DT^<O]i01fT9K8J1fJhPRSR77E_I_ZNeI_VSJJ5GlQkjj3;9YpA]E74
nG`Jf_DYV=BMga0c?>?iAWo:D@6LGoE;]VmYP;V99LMGeDJpO4751]@Jk4aY2hgK
9;2A\d=832VoSWUV1BCm:JBRW:GNPb<A38p[@n73`q\cKK_Cemacn>WfYJFg^`fg
hXm_@qO>G4o2]gkac^:0;K6f8HX=G0c]acf0lOE:UkpEiRXG6\p]DP8:?qBLD;AC
kH66:G=b:E4FJY[QoOmDAOY^:S4Td3hhcD@g?hl]kA;fm@GH5UmE>oNhXFC^X06<
QCq^;dhNe\3dJm>1=6nKjUNHh4Y9TT?\?cYA9:W7hZ]3IWJSFC<]LASO6bTL;GNY
1<<Bi4Be0;TSPM4Ic1bbW;TT;1:9YXqJWJ]iCNR9l<UQgnSEj4ickk`?>CO5:d?l
dTRmTMLmY`gk[R6BTEoi84LQ7OA`1ie`BKRW0KSFTRd><2U2\b=FTgmPK5p_ZGPR
;Rh\XN:CRBHhC4W6QOJF[6>n6F9YPG:XB9oHIFH7WmYkKXUlZM;lR]S?mWobR[aL
U@M_a\@1X@aS]F_W9@6DXBp0Y7nD6Q$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3B2(O, I1, B1, B2);
   output O;
   input I1, B1, B2;

//Function Block
`protected
WY5a[SQd5DT^<EFRHCF>P93G8NU]363Na4B9jai1VI9>Q:a9We<f4RFIq7NJQeL;
^D0@hjJGl0miLkO6O4h?IVaO>;KnZh:`T6Zm5X>VS<5peX=9heYFW>Ml6S@WWQ0Q
8V3BI[e:pflT\bDpB>]Og^eoF4kW4MGCb@VM1VDWH]:pMaDDZNZh<gWm8e`GWnU_
mNB7O?B^5X]mXnX8q>LF9oZN]@;OiLCBX1XN>86WY@BYpZdDK4\<qRUAW64q9jOa
:4hf00V?HlFY<W04ToXKXFRX5@>=U:SL=FITL3[\hFE:oE7NC3hBVK35kmD1915[
jNJ0cQO<Y7S@F:<pb;>^g_T4NICe>J3=?G]GTi<`Y?=oagke];j6_nak[Q>i`JnL
Eja7Ud8O[2mR<PT`RI:gZ]4RMOVZ<9ITN@B6QaTpEa0Fhi>>mZQnS6f0dT?iGb3i
B@EXB7cWlX8f@oHi2kbnon8lLg1JE=QV@?GUd8Yo8^_^?W__UI:SNMhe<\H7VEmq
^9U6QVWN5B>93E_63PG8e`1a8BJlPhqVj6ZXg<$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3B2P(O, I1, B1, B2);
   output O;
   input I1, B1, B2;

//Function Block
`protected
gjhUcSQV5DT^<HVYV[g8WXSgVW>nXQ:KW>W8G3>7>Aj`HlUUWe<f4iFZqd@GnDUn
[2Kd`kBXgqS<_PLP<UhT^UaF2a3PIT];;NY:\RJK^ZX;4N^h]=T@P;UI5@Doa5bQ
V;YX4q9;HFUjqlHK5e\29NocYEYZoKVoCaifC;<aqDdUCGk3a0oBW<dS=SU_G5[B
b=4G4cNhhFPW[qWb`TNmedP<Fi\dd72;C9?G[D_7hqHA<llHjqZ874=@qCZO;9eX
dV@^T1Bea]L;??lCVWhHAeiF9d[?Gm_SE\V_=2Wh`WJ3A@6_==lLaGX\6:^AHqnB
I0P4fOGDUj6NQ63ZoObIUIj;EX>NJoL@C@7??8\l4GWB^QmRnKM@XYKI:EZV8DI8
2Em5]8iRTCT6YDM_n_4@Eof`epgiX\ULf_<N;Zk1RdWOU269P`:h:LS<bCKi8@1P
mJdm98<1So\RNREm]61B`Yc2kAAD@eglLH8FeTY4ok==bm^B5A\NGpQ@5BNGKEVk
fFZh@XF\CQa=o6GDaVEY0fZIC<:]_fJakDD\A:DTgeL=PLhh0k3eTO3XNJAG`0S0
1Gd]@8o\@O]b^?_AmqV<je<36$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3B2S(O, I1, B1, B2);
   output O;
   input I1, B1, B2;

//Function Block
`protected
2o]edSQV5DT^<1ah^UTod=o[PBjKjS;VfFbbl`E;:;C\Bmi56=dg:W4phjR8X?BZ
4S3ZMH9d:b1=F`TokV;>gUf0GIMU>C3of_gK]AdgP0eTgUY[0g@P:;fp3[JO8G_\
jL36;B[7H0V:4GFH0nEfnWJ;5GKi>;VAJiI;J=KkV6ZE@WRoNc[3FP:ETnp2D69S
lpnXbATYdZl]]RFF3ZR5Bbc@0=HB=pC@5_`cjDbfc@W@Cej;H1@LAc\WbbVgi;PZ
[Xp?E7ZT?M`=?c;[R?l?aOe@0B?>0Fq^E6e>lXqNGZPACVZhjeQ2?<6YCaME1`Mo
hB[LYn`aS_Gm0L=Q>RFn_K_f4<UFDk77SeZcd3ZUK_Mcongp]OBc\lpCYRF=`^GL
0GQKd@<?3<B5X>]IR?dBVMgZJacVNlaOMkmahCb0U[X6Gg]S=>ME=D^CUcFgV8b;
bAYldG@M=cq0eU9Y]RaG34cMH0`;eOWaX`=`jOCB\2ko>0>f]6MJojXF1QdK<mOo
PDVNYTchb?G0anTB3o`jfFcKj<ZIhcpn;Z9nU>hTeJdcJSiISSW:aecm;gIhD[<C
CD6<;Z;TGN99Xn>1I1dbmMl\1X6SU:lnbD?3QJh7c2IRiZ4:FEqJDg`0?R$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3B2T(O, I1, B1, B2);
   output O;
   input I1, B1, B2;

//Function Block
`protected
3k8dISQV5DT^<i5aaCLC\U91ee?:VAC7MkY9AY:eJ1noj8i46=dgfiPp?4f2kbZ;
8l2o<J2g6T\XEPA15__5iFWCS]0=;>dK;7Vc;M;oS6U25_d]?[V5hcQhG8p^fUk1
FWW5fA5;`pK<9i3`pm;K2ZFg:4INe=WaBlS5feX3_PYlq[dmNCWfEFDD=\B>VZRM
IH?3KF_4RN]PVPa8hpn29Q;d::TfOVggRL6fG3i3Yhd_Yq;k]H?>fpWATlg<q4[B
GO]7LNceJ72XV=kgUb31BWF\l9SOH4PO8U<]oKW0UFagYH=V>]DjWSDj95c3WNh6
IV46P`N?<Da6go\82fAC>;d`p0[0O<\cXAo3k9A5:7ISD?=@0Mm[EBShH5a_fhol
=LXTo:iKg]fb^8==CfV]=kSeD2c3U7oJ?GI4[`9G`;US5C\c\e]CpDBO\AiP2Bc\
AeFh<:E;NH08PgG`_H06YMaOi[LNRjfGfVk9TF`KSPFScbm\bR5i3lY`c90I9D@i
b\;;G]5MCkbVUm3Pq]D\L@3BeCoQmO2Af=;N:i4jO`jL1ZGAWNo>h9hE3FXSLhk:
Q[TpI`Oh<UE$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3P(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
eOFE2SQ:5DT^<OjK@DDXa5IEc:KibCRAbinB^NcRTGnOjK8oo;C[J6p0Vm8iBk7k
_]=3jjV5ilA[BC3`6jf][Lo@45XGfh5Y5G2ZAn4<S^8g`A<J@@3b^5qCJETLm^1U
63XBbZeM?`WCM3>4`LPY8cqHO]UFbq>??ml1m1;d`]<^K7IU:aFE:\GTn]jnBeb9
AoplOimIB8qi\nH8Gp7PTX^Lj:R74EZ>0Pk58W<NJPlBQ6G3d2>cZI1@E2m:V58`
IXQEkTPBCCj93MVMo2l_IbMF^_HjSAILcB=gEEd2;R12@pS[`LdBQKM;gY`EDS10
l140kcV2gg=eD69MNJE2BIk7OC]1bZG<8nqmFeF6\jggAbb58;7?3oF3i6f9@`_^
7KVA7W`Tcaa@Ym0R3M3k;a8F2_0^VFLfPXHWX4gAYBbkNXi6@BU[P_T3dBncQXqh
3kQKSBg;<5N@7KXj9G]:<SN]@o]gK3?UUI`4]9PjR`3T;ZAn5Il8XFk07C2h5C^Q
c\O1W2@jn^TTal24:2R=B7VX8=pX9O9Hi?$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3S(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
<i[eVSQ:5DT^<k2DYgXHQEDeXDXOEV\OiVR:@MaX0a`VMYc?m5F=p?Nm:<hiBV:\
jIV28>h?F3IdDg8YWM6kQI3pA3m]\:aBJ3^k^L1Njho]MZe\[DAVOLYK[:n3XM`0
UPLEM\b>q^l`JD=pglLNO2Z:`fM6e=<5Q@kJON=02IB:Ed5hG8BYqeF>>^UipmnE
m>7pXT^:_@BeI]DgchRI6HI=RKgknZJSho]f[k6lGk5@H5a4HYga?BeV[2abDPCd
BS^3Xg\<N@1i6fDMN[JV^;OpoeMgNoSn;?7QVG?>I8^`75gfS=AlgnbLH28aD9hB
_^9FeObn9BkjCQe5Z9hMF5S6oGDYDn3\c^R896>T3\oqocU47_kjk9:4i8GbhGGE
5J<JmKnNO^JTC=]QBf6g2CHal5T?<oPQYmUQK5]FQIn:oCI1mMnGbKdB?E<c:naq
0LDlKe9$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN3T(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
H2kJlSQd5DT^<JK]WWJmORU?^d19;\_YPDGT_4[6THT3MYc?mVFipOEb7^MTP<Pd
EL7lc>:8AROe?7RV=hNXN@?PAd7qgj3@`jE<5I^8^5DAInbCI@2Pfg_56]`Wcd>9
A=6VFEMST1qSboZD=po_?AmHb:LBnIjRIY\N6YafIRYUihQd8>j>`Yq<U`jAEHqT
?LH?>pQG05jfI5^I>?Y\<9\;mWHI3YPZYX6WY5aTfZWaSMA845>OF0<h@:_NO]lj
0eIcd[^hn3ga^:^FTkF?CB0=2_i@7pF8hA0<SPbO1GPD_bUWLD8J845f3PY[<XC7
`cokME8JlJ]gjM<7MUTdf5Xb`jk`^;n4SVNZQEP6U0R^=NfjCPiIAG1f;qO8_6Nh
ZFMW\OoS2T[bZ5V4OXBbkbFBL?5@YoVgoJZ;:3WDRN[41_=3i81@JbN:>]NThU4O
_[Bd>2OU7P7gXfDlYck`_qaGfaL5N$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN4(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
YJeKRSQ:5DT^<KFlR@?D74]ZSPemH[YT_^E1]PAeZJBZ>YV;EXiqn@lZe\cY7Fg7
E5]dE9cFICYLi@4<qHPD?g[i^3Gb<0VH3TYYQmgLC8o;RaZe_DcCY<MW3[Z<8DWf
1mOK`190i<?i4?5@e9;dS?Anp4:@:Fbpba>Z?3XK3f5[S@V8AaN]YBb]fYLdm7cL
j@AJMl?7AWqf_PUHKcp7aP_>7p_R2VXJD@H\SPDQm]l=J]ThO3hAdk8_l8ZaigBV
m462VG_U9_TdXkZ>Im9kf7[8hd_3EgWcmPMbMH7h1?HbOpKb2_L1Ee2T?g8G6Kh[
o4^jq1ND;[QB6e5PUJGeOk`[Y_8b2TG;3`YF?ha^4^<mNjQ6TIilJ`gNR4^5^g;C
[`W;61:FGkMGfbJ2emaMfO8VpOa3GK57ZS\SoKjA1<7VV;1V^VU16GHXa0kbK^dW
TbB]=i7?eX\GbI:cQU9c]FY7gOd66Bi8Y_@ORVAWN;0fq^gAeKCSg@:NY@X3eEf^
;I<:C^S8alilb`DUVGbQ\d<Cki8RLN\\PWXMX:XFLZ8MC^L=biVI06YW;<NL2``g
pY;S7kC9$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN4B1(O, I1, I2, I3, B1);
   output O;
   input I1, I2, I3, B1;

//Function Block
`protected
>gGDkSQd5DT^<oi`BiGDA@5<::nK1AONPh]hMa4f_6BS>YV;:k6qV5m@[_e2Z`3<
jNg[D27>@N6W:\0_lZhXpQ8@H6KNIf\l3;g`a7D1]m]>LW:BkGLR>JSl1h\mQH5_
9A_T]o_hk6Bp;4Q64Oq3649U2cfJT7Y<be^6OD78SRHdWlQJ;`d5c8fiPnHM0pPC
IV8MINZ01XS?1Yc56kXOd\>dlp[XQ_ZEWRMk13]DWb7WQGGOEEWB5I@Q@h=M9[UY
qFDWT=U3pN:YDY?q^_QU2=O4<J5C\M@AQBgJNd6\Wa^CGKCJLlCg5h0?=2N4^1l?
T:^jO45W2Ig]W]kj^dBMT?I>I;D:KbO0_^op75RaF\KgZ><cgb:?FKCA93?ULZPm
eKdEZ<aCbLcgCWYQ8HI\FNVOC0@CWmXOegX87<Z3\4c6:D7YK2BKKkipC]0bCKE`
CCE:JUBk_[OdNaKQY4oj6\L8;FKmJ0NQI?D>HdZj9GGkdIA<76GW`KMkC[mcM@Lh
WdmR072iPBZqn=:jPPaNACN1W14Q1dGlYT18CeBFKZ>5gnjD=@TQWGj`1Ah;;SV5
Q:W5ncT5]Y]Gng57o<3lgBUETO?>nSEpIXZd`Yb$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN4B1P(O, I1, I2, I3, B1);
   output O;
   input I1, I2, I3, B1;

//Function Block
`protected
C7c5TSQd5DT^<ZEljCf1_[iDiG8PjUlkMCQ6>LP737SM<l?Mf6pk5o_QZD_[6hAD
;MNcMqZlV>]79N0i5[M9JU6eg>06aEe3aSW^AdTN]fWLXZV;I4ClQ=XgLm5:Tm5d
E0JBOp9=LnC1qnWZA9gkgI3f8LD=RR0i0:gVfAOUHLYXfSm9\:QcCO=q3kW93WA<
[Z?GKZ[;PXd2dm8ejD3qXTX?U[SL^<>cTnUn0mPRB6W`:?Tp:7FYS@lpeEK4;Bpd
omeoBNJ[7[n=mFP0A:J`ANYUUgOGUnUgDN?Nj1hi<nJ6?8hbHj`A;<nCZQ@@D[ld
hf3W:aX7;[gCS`]EPoq_nDIj6_c[OXdSLQq\ldYm7DDF;U73\5VFfO63lcM^aJjG
H4M;9399O9PfQ0clk=T2<khG]\LP1O5VVnY2>RAX9iff1B\GaS4CR;9;=Ap><W3n
dADZLd]8oE_[kgUI228bi<OgQJh;[HINn0QeBANmXZ3[6b;c391EKG1@ZdWF`O9J
l8enPV4m8MdY5dH5R>pMIZ[EA@PP@PP58CLZgncV8>K9oM5<kS>NMO[JCZ5S:M3f
E76^W1U@@<?@NYY3:bPMN^B6i0iO@05VdOE;Y?p?7\DAng$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN4B1S(O, I1, I2, I3, B1);
   output O;
   input I1, I2, I3, B1;

//Function Block
`protected
@c@NUSQ:5DT^<am:1T7;I\c_Xh:fXXjS?J]S6Fkei7S\<l5MI6qjLOk1=MS=IK_o
]?Q]W@S^0P\NVX@U\XpmaD<AMnVooY9H59\:MMKlK>9DIF9ZNQMe3_QhHh7]9>>6
]TC`OB6Bd_WY5eUp6WBONcqjARWdSbj_E5b__D1T5cL<`EHeP>`\cT\lAYZ>XhNS
@pmQjULRlB0FhGE3f4?HlKcC\?XVCqKok\TMBqBg?FZmpao7E[I_g5cWSAB\9mh:
bg8W_QFk5K68c]2X^m^qAg^ACUlik3ETH;M`RSn;29K>Il0[0640FoBoGRdjRFhN
QW9\1=lnFgXGM>15kaJTAP]1ejCG2jEUlWnkRofp@l0\99hjenF`EU5K1\@PjIG@
Nc\IL7]a[bd@Rj24Mg_gW0`VbLd0VQXCYDC63HYP@eI?AEP@j4a6dCk6;EIpl6Vi
D;NkaO7GNOWX59?<iMBU]XnH_P^hkXR2aWkD@m7begM^[5L8>Sl6\TOZD?[@lI96
92<?b3SdT2Yo^4Pq6faGXXZL;Af:Vn?pFn\[dHQ8U]0=;YX3[iAjChI3^ib0J:1j
RKPalTFk3mS<Kdb1_M=_aV;7h6ObeoIiF7iUW[M\:Q4A?TT1<?mqd9jm:YB$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN4B1T(O, I1, I2, I3, B1);
   output O;
   input I1, I2, I3, B1;

//Function Block
`protected
[P[\LSQH5DT^<0b`icU4GCNKe_?M>WM8_iS]9[?]X\i??m46pS1W78hlb=W]R[0^
CVF4cqo9j9_RP>5M8GGemNIRfY1KOgUjAgFDLbJ8XfX<iE66l2X]BJmVW;R68X<?
Bq[b05o2p4DJM`DBYH5HoZ8YY:?iT^O2fDb8df9J1Wl;eGlUjUQp=coR\c:ANTXW
?90bSha@LbQiSGPq>=FQV9gpUV8HYmqTA\=FUb3UAkhDZVEL>l]igbQoLUHnDWH2
JTObOQ;7nhT_HOkS9Qn8Gh=\mE9VI=g?LA0<QYcc\^d3omBC6676`<qe=]Mc3He2
Dj:4LbnY`;gY;]OXFhZ6VL_?STJgTn:U>OY^V_:X4c9pGh6Hj6c[Ui@2m=LN[:jD
2h?hOGDKaWP=`aZR9\:0D]`J_2W8<>\[ane?Mj`H1OlLSZ77V]gYX@6@dChSBD1l
@jmq>9>AB9i>[h:=W\8?>i=]Rof>_5McR[k;X[`del35MRAm0:b:gQ2J^VNdH9Xl
UCL_;g=ncA0NmKlThEhnd]FFfkXpOK:OFBQFU0jOE?]a?24:K3HXYTQ<4BE>l1i6
n2mF=QVDlDcL]R7:>jIIgMB]YdaIOgo764l1V0YOUTOdeU6pZ^;Z>\U:IVUDlU^p
W3I?=Oi$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN4P(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
KFC[HSQV5DT^<NiD:TjX9l=H``oFM74eC:4h0\73X\i??IMWp_>RHCSPk_nR1bT3
B:8@7YB6`Fm?JM5E?A0aJQ=EpZfPY8kT495V^6f;j`XJ98gdNbmUR^_4]K;?K:jo
EJlDfCVG4GJ__k04Z<8[AeV^Lg\<ApJSo_Fbp:hO=DT36PW:Od>02?=gR46`>YPM
QBEQn_Y6god^K_WpC@77d\hq<i4PO1pGVRCah\?FKW6;@mLC:M\OmK7K5g_m::Ci
mW:MfbA]=55bQgH7NHK\Zj;7K=PE?GJ\E0@MG9k1<X:oBH:eSF;ShVqlY2joCA_Q
mG2[RhkVVZ8cUM02eUA8bclT9YRcId[T<4im2oO`PF09:130iC<URJ7VNA\AUB:V
QBD=GAAQVIBG99pFmlZbQ^k@j76iG:HG;^3NIn5R<ISX9;;IRo@NQRQ`U^oMPdUl
QGTbQDkF3lYc?;iF3n`5;amj^1V6CW2jKMqK2WiHIHIlFi3E9ZTd@WLlQFgQ1\ke
lA7Po=O>?^aRg27imlHYjE8HB]DQfN>AKh@K65TdG=@Pm5>G5kBKVhpXfAjnLB$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN4S(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
LIYB@SQd5DT^<o6aTdSSW>mdMFmJGkaGmNTSE1mG\M`d1[Xq_`T5X>XX39?Q1HC3
^8[ldMiY8N2q?NDP`0;jfag14FQY5_hec338?73fcRI0oKGN^`5aLbJ\d=A=5oTF
JI\<DJg<A48BG>9MNm7pJBgJbDpBI0_NgD4]^lP?]VmUO6bfJ6SFlFWVcF2Y7=g_
1[?HdpBLn<_^cp80g?CHpn0LdZO[oSZT6AW]`3JR@kdDoei[0``4\L`K>AU0GhhX
eZ@R4>FP0IZ[IN5Aah=d\n<VA^C\HRN_Eo@5GDkCp8>ThLbA4Dl0\3=A<>g`j\NX
DLhVDB1Sh;_\7J;Llj>HaIYZIcWW?8m\dM^oh29aW8eeJX39IdX:;cROLZTUp6>e
bWQ5`mfmMN_K1E3FUTeg]VPYmJ\S^:XY`[fMEoQSNNN1eCj6]PBNoDF?B996T64U
dD]INXGhaPe[`J3IqjJX0a>j2G]B?c[?Cn8hmK@KloNo2R<o<T8Z0Do03m_4[:8=
kg^=eoGAEFof5gYk;OeqC=Qhb_mOllVBZK<Bcn<2J]0@KDcB<M>\8c=cG8jP@d`<
`MHB2\CDYhQ4Winc?_agCJg9Lo?UD:VU8aBk@MPp0Gm^@>4$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AN4T(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
;2X0ASQV5DT^<g9XD8KJR@Jg`A]SfG8S3chC3RmQ\M`dnTEpdiQSddH5<Z>XhdOY
^EjP]0q;VS<\XFT8UjC]J2H8[=k2Sp]X\];=qghgi2LbnTg0`o:UnaO45aUhXCVe
ZeY0FEO6@6Ac<81q01X`IX?pdloiD=p?k=bCaS9;:3Z\HiVBK^C8<\36_eK36LPB
flABYO2i4IIoN[?WKfBgL]lU?kcS8m]XEWgXT<[o<HV_>_JhC1clGcqML1`1CX]5
<AS<kFf05;g=^9i3F5HAN29O5T<>5<EnTl]?O9SL5U8_6HfeOVE`jS4m[^NmQ?^R
MS5YSINAmQ8iR`pOQEl65e`Mm0MLfVP4C\j6Me:aJNVho4jP95VTYld_ndiFR81[
fID2FoF`W`fFHmb07FI?OC8ofZ6;AI_6I[c7bQqA:LadHVHTcLOn\H@7J7DidCEB
eSb_8=H>9U[jE5Df<_TmAaOKeSjbf@V^<`B?bYZa@C1=<lP551c2W;8X_@_9^QpW
W>jf\[_bOSg^nl;\2ggo1QlJZ1WA_P:_npENNm>GX$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ANTENNA(A);
  input A;

//Function Block

//Specify Block

endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO112(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
WZYLYSQ:5DT^<4^bCT4cg8ABZU9><HPaXCYgDC\^TS;TJIp2LF6KHR>F<O[fbR42
[T:IRU?_Sb?92p=AOUM<MWDkRcJjR@f><\G=58FBXK?gJlDfXA9``5;j?jQea0n7
hpZhA6Xjq4Sf[^\Rg`\H787[Wk5TLWPjUR\;Gjdd8_?pS]Xd;hE?Cc7Em;GM<?mf
cb8d=G6;J4<e@GRl6iD0pUWeO1n>W32ZXfL0;J5:SGa8jdlpPGc6klQUZfTS>M;i
g]g>3T:U18NIPN7`T\0CF8S@^>:UNLQg^Nb6>b>ajNVmM6BD:>fqXSE;ia9pdhgZ
bVpHDd1e;eAMDib4^n_Unb9CT`2e76LADXW7Pn0:]SLC>:XW]L]RB0B9`6I6j\<2
:oaG[ffZ`?7W9`>i?A@b0P9_[T>AUFRhI=I=18Q5]Q8Zl_?bigM`bl4?>Xc@5q>F
1M=acicVdJ[jA_GhKbO3TR>0H@o_k<i2eb_3dFZ^]kbN2R<aPIX2ZeYK`9EY86A?
bX[_L@<S94830d6FfGKDLNg6S56hg5kN2Fe3MDfZI2icO:ifanmWl5Y\p]8239i[
IIST2Jfk2?HUDmViCH:nU>8EB42?48>Fh:a9P5UT_:EaOLM4<iRYL\\ZG]n[3bn?
DmF0UnEX6HaMcdD7mRca0U3I6B2546f\Ihl3YNZHZoF;3i7q9W74aDeNL1eT^=PK
S_cA3L:ammQc_2C]HT4cjQmljCg\A2;IKG>K@60CKeM8Gd1V9okoP0fS^G3^<KX<
Z<V?SWp6Dj_koYVcSEZDA2Ng=Y^oVk60J^0S8OgkRPRIJc2KA9TjI5Cdj93_6EK1
]dG>fG:65T5`YoWG:PLQUXV_Oc=dMOl7;d7QF56URnlO?gXZNTC;FO2hl@YoHqU6
Hn0VVO@nEVP@jpj4J[6TB<jcCFAb0loQkk:60gXjML>`^hhThm;Dfa18Ji5iO\MB
X]gYZ^>_G2:mKEjELYO3<A[BJO>0l5fI1We:FX0\5E^Om?gTliaHRon4eSa;[IAE
O;BZqhn9?\6_6Uo:K8Ef:[U33hZLReVK5R@L8S1B^UfTLC^0`O1I6<lZUCO@b1_S
L288?hY6NX@QDn`K6OoQdhV=LJkFCVJXH[0?Sj16Y5S^45B_bH8;S_k0JKeqnFX3
6LlFC35VBbn;4]4KVC4YFQ4IoAeTle`\9?2DADko5VFf;nQ\07ilX58`^Y_\n:N;
A1`0\7DlbQJn8KS=IDq[bf3]Cp=Q2\i@a^_]GWR0PeXmjH2I8ea]T1`>YR9[aYTX
hb3GB]6]d0UUN1@a@DlPfI<oZI5QVF;Fn@VLf8:6JIUE]Z^j8pHGUbchW2k>;jT:
99f^=]lJ1bNOof^>jIEQdDe>G:j0dL>jm4biNX7PaV?A46IKNUa_I`0bam?h3kcP
_:60LBJ5Yq;:ok4\\$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO112P(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
^P^STSQH5DT^<S@aj5[^S]1:56\5JOiiePXWYj<2Q?Nlqk:WCH]e?^]Ugc?E>o?0
N6;m@;fW:M2fk0AdqT]\Q9glbj[dV=KiqaeCF6kplamRk4h?HeeHJ[?l2MhlWVS:
CVZLJU0<:Mq^D6Y2Ho64jX]1fF_bbTkJdK]?<oBe<d\@ER5ENAhqOO4ePP7hg<fS
OoZg1Rh7@kjLABpJm;Rb^cq^GQQgHpT5FKh<m:_md?IZ4n:n87d7A;7X74UElfdI
;9G_NRLPi\Bl5GF_BMcfd`F@o^Y0jDV0]hF4VW>=:6EH=RgQ^0S?FaKg]_`Gl@O6
6Q]_FU;ZgGa^>5IoUhbAeDPDp3Mc2nHPPGZRI4d3jHdEU7C2KkSh2=4d8MKP4N5>
EPb3nQP4e804>ZfkZT^B\[D?eRo3Boaj5`h1k_CY\0n783@EB6L[F^f7`3N66`5>
BMNaWk7Bee5[IQSJ>N2q4?iJ8K2]bYWPL6[^?FS0A9bC4YBVWBZ;^h\S2>hc[TfV
gTaiV<7kjG9A8h:CISpXe>34e89lhGo6M6YM:91mefk^Z1Af=gfg>HWOT;2eEjCS
ce6JA[H:7^77<DfA0d[WhX0If12LO;aT9PZP]4`JaRbU4a`XGW2^B@N0TEW`gZcR
oN4aK;ggnkb\Iq[>T?RB7NoBCj?XiOBVaSRoiYb?U9Y3kQ;[FMIEoCV3_cHZRRUE
`WFdW090cPR5ocWGGQh<]lG^TS5PadHh5W?[a>3Wpd^99YD9SQ<^8E]lgbfAK<QM
7:RH?:LY4EjXBe<[dIhfLgJoZCO4DaG_[cSooXF]4dG[39A\h[QQ5Lc;O<R]V2i?
GCjFef9Un[jOl<[Dd7J<GNk[B74=Wdap49eR@8QKP9[Eii?@1KQ\mj;]aRZO_7@2
CZQaQEfG2h\O08Y\gjH9?U^gPEKWYGS38Dk=o4Pof\VbX@Z[=[?c<R6K39iS[OX8
bMKc5E_B0Q<gTS6N97A[mh22OSpfLMEPU57h3?o;Man9L7b5jIH2Ph?`lLfdmSSF
hC0g3m6:2>2Agk[e?A3GbLIg7g5YN;Sn^nW??n`4kg0HlD=QWaDBOK^acAMXh>fS
h65:1M]FmfYK7m?`d_RM=qXbGUM30OiRe\A1D?=X]^CcA=>Ja5NVjZmOQCHZ3Cdo
lZ7:S@hlJg\FojS6a?3^WX:O8Q]GKVgiY<LNXEa:^OP<NcVaq`k`@io5:5ETTHdl
IbC0iLWSJCWGinb=dd>kpb?j]=9q`kT0J4T>ik56]Zi\PNMn9doFhU4Ead\_<\6Z
J>olZ[MSL\;eG0GI9FEW9hRT?Y5K\mV_0_<]\\<KMCjSOWEf<KZpABC@jKZPhRGk
e_@?7C]DSN6j45jeS9hFhkFe_gQGg_YX63FEX;e0F:A<WQ1Ok0o\9ECUE^F0G;Cj
HVMD6@^PbSApYo=i^=R=:GoNPYeEM;C66fTQj4N9Nm;mbNg1Ge_APoHb1KI@lE7S
0^fRTG\`c[cFO8[qQcLBVKe$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO112S(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
\^ICUSQV5DT^<M_1eVVBb6NRQ2NVM=V^e6FQYj<2QjO`q0:0b@TGC`o5WgFCPF7W
Ncm\N6`;KKW25C;jobUPd`gmJpCJU<D4`0V<=be8NH<G<@bIpWLfikRp:EmjO86C
gQJ;]41VL[dC>oYEk5@n;S_G67pVe:Z`C<]^f8_P8\VQfXi>^;UPa4hXAI`cN57E
]IQq;AFiScZBG[SlCZ@2mS_YW\Tj@=p02j^26Rp34faF^F1<0FJR6Nl`<;J1C;kA
le1X0JdU_8UjGVdnS>pHdID^Wpdaa9V6[FPFf@:\i8[]U6KmbYFf;A_CJMPcnIBa
jW9BdDgU:K^?T3FMW45b56kT>Yi<6OnWKGjUBfjkh\=SRj7D]AQ2962PY^7BVHUa
CW5[:N67i8jS4RXC@FOBp`9G3>>][?QbXm^R@:dHe2Ve3o]Q`_[dI@ZoS4T;:eg0
3flA5C`027B7eKRce^WGcjmn;UdSNM\j^iL3Xh9]KO4`?0I4n9gKdNVmN1T2A]f`
091oh;VJP21S<@YqKGeMUkZ3L2mVZ];WLP3HD6niaN=:=PWPVeGN>]^=fZdIU3[6
R5Z7L682b0dVjhfjKaUMMkmm[6hj;8>_5gbAd?i`l?c]B]Vj`e1PEm]lD8?Ygc6M
8@;FN9p>SJN9`[jlA8X0geK=9<L?3XM^OSljINdQ:9oBD]Ukd9@Tgo8GXb3deR[E
jJ<QXR7>^jjUdiDSeTU\D>G:NAA1Ip>XKAa>@C3^0PjhM`Dab2aFj<m_kGl7cHR1
`lGEX3P88`;de_50nOY5?]LKk5Dk5;>8YFH9c[W0aWaf4Ud[CP:Ra;d>QASb2c^1
QH1`98l@D:Lj;Em]KAI1p^>SIbeIDZmQ>MNO^YYWDMReHqh;PeBGBL0Xi1Y9ZX1V
TZc;F8m1jJk>E[WCN3A:1ZTM6oo]1gnN4Vj:I6]G09UT:?hLjZm2Y_N:cf52jnlk
cTYP1_n95KY2BTTCKVIg\@M_^n`8YE:k0c06qEhcfMn;eSPM]D99C7Y7bZKC:I[H
JAP8S7E?5PEL[g<[RUcCO8nP;56N?^e3MUR:MEH3TbmJFXNWU\WGSmL@onB\>2^Y
XTM]9eE6F;I6EZ@l^MXo2AG1lf;qbdA_DlgaENVa@f0QCZfMO15B7E[QTU>EnV[\
M4_48`m27_Fnl`RknKg=47oAhkkkb[nZ?dde0=^QVBdB`o@NeIp[`@DncqM7[X@^
74fnXS`DeW:mh>>ZCg_Q=E`_57jec?b:_\LSX=5fG`5Z:kP3dPjH<C>6V=<g=kZg
BROXcUB]F5S9I7QRBp27U@<VdPPGmlXe=i]S?B8g6J8`80?ZBn0P\5od`Aj;]\of
^O9VfWJ9NfUBYC33HRTT6R:VU73?kSlX1cD\k1BA^pRbPiV26$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO112T(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
YnLF8SQd5DT^<HIXBCl1d1^CXOPY2ljH4YJcIdP5Jfop^fHASdecFS8LiK0I2Mnb
cVgCb=h;fo_1N]V6meKiUVqU;aL=>3Xi:W83kE?Ya7_`Be7JZ?\iF9lE9Vc<7hIn
74B651=qKMf5?6qmOI]hi`EoFAndb2\iBZLej_5[@YN>BPIQ^p>]dV07?mfknn^g
QH]^XCAQdZK70NNgkd]lB>ShA`p7g8F8m1\[VTk67dDlYRKARaF1A;CZ2HcPCl6h
WU7`lR0ScEiBf;N=<i]LEDqnh]26TK\Z13G=N?PT[R2n=4bU1pVV4eZZGpA>?h\l
p^<8g3l_TjF^YVO^n542hFGM4JEDA06Fj@@iAeI:6DBLPMVc?`3S9TSD@SibmS6I
O6H>H`ni^7_I^07m^;4j4k>1kHdLiS?H@coW]8I>;c:ED3MYdhF`MPJ\kA:pf@ji
1H_U`;bg@e`L]e@T[NldGBH4@OlPVfP;7P2K:T=ZoBmXXHoo3SX3FnU3Z@0icU?<
LmZ1^A7?I2PM5JHJ5`<5_9WA2\CWc;iA5P2bMJcM`VN6:?A^F3V1M6pU:V@Xi9OE
IdBikY2W@OoZ`b8<CS]nRcO_PEj<XAFAFC;>OF>jT<jfY9JTYm5DN5D=Q[ZV^E77
OWGWm_b<V<6JiJ2>P?llLWblJOW=XCnXHhn8ZRUg<Oj?jKlSVqXImU@:\RUfm6AP
XaPW^j:]l@Flqn`1ZjTjBH[QgRD:`PYcn>Z39IlcY2i@E;U`MPM1a`9<`i4H1HFP
dmXV<CgnWfQLg]3I0JjY8H]LPghOQeiW;3a`C8Ip5X?Y7DIXAE8?_^Glj76Uf3iR
B_Z_6jXSB2WP<j5?YLfP7HiA:ZRJW6faIZ?G:Ee@@gU9\ARH5Oih\1DjK[j2kh0K
25Q5GhieQ:3dEj\gOC8CeFN7EUE0lLWe^GqlDa9\gW\NcDe`::C<O_PO;J3eVL[l
99mOh\Id=l^?H]WC0?DVN_<NV=a]3TK]1jDJf4^b<VK1hDJNW[QZeAelRmke:U?[
Alg`?8TX=hKd9B9>RB0l:;gS:`mCYqW5_E2=[BJXJHO]D0g[m]6K8K5^j@bLM8gA
f8<l999XNAW;^dC8mP349<CN^6Z@IcCTi>M[[M_M]OY]m8AU3\?c>hR7h=SBl[2H
2m2lbXIBSN8_8`a7ccZ\N6AKq_a3C36fCT7\Kj[MSNTI5g;^RO76mDR8ecWbC>1N
VfgJ\T<RYObEU?8e<UT>[k_Ale[VeH7jMR1?lag@CGHmO1MOQ8UqKj6mA:GCBLDK
VX2N]CAQN\6WEZ:mMJ:WK6g8N0W2GOIH3G:gg2>n4[CR3f@NKISb6^q\_KIb9pUd
>Q:?7ZmVNV2<9lhcMH71E>b0l]9Z_e<KS6U4mhJ9lMkYD6[6>l9=`BSl[8Fhhdf7
8IaoAQcYLF6?dM=__dda=pFiX>lN:;`Pfg6WRE5V9\23=l]4lW_Rblg9]a]JCZXH
9>:0J@;?JHEaYd3cS_]9:chgPdSkfTZVP=>P_e_V2J;53A7Qnqj35EKcf$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO12(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
gj9P0SQd5DT^<NfD\6f90oZDlP@A`D48]\J[IdP5cH^p3OQ::F5=Ac^DhZmA3>:E
k:T\2jdGYB?7<lBLpUA;2IDndkR:mi_WBZg=Zk]\8?cW@eAXNh9mJqcWYaNcp0=O
TQPBclSeOiA`mTNnehF4]87H64NPXClq:A55mM5ohDm[eXmDA;U\d`7JLZdmB<dE
9<pF1TF=7D\o9A0Q389l<__CL\48Wq5Un3VA3qIX2=CSp]B<\8g;Pn88`UP0;FH@
l1de<?dQ6gOTVhaYDBUOS4mV`PYI4Fk^oNli<U?ZjoEjO]=FAmm8=Vo7D:fVT^k>
[;NF[h`nm1dH3@a?D\:mDl=UI;TijKCGL^Qq6ShGW2[7Fk\1EE5LF[`L@H]CSbF@
Po2fLQEC4KoXE7^hXh1:Kl_^^a1gjc7R]Q`]okOXl1R7P8@Ldm:=oRn9?@8IjjhX
nThnm@D6SKo7O4`13MWeHKbDii305aq0i5[nX=\8e]^4aDcQ3CFc;F4hh>@UhA=M
APKgkMgSN<0TP?mg[HOIGLLP2F[h<mq]o;2S0F2[oV62\YeCf`cQ\>]6iV_Q6HBT
GVVV0hC@iJB6T8A:`9Veg=3A9]mlZ6?dS:DE]o@5@og858Yom<N^fnln6YL^dn5B
=Tao0`VWQb^Fn2l8?nlVXZZd0q03e^BkOD`0[;SH]C]ZT9V05SF5TH0aC_FYSF=:
o1H>;H<9b4bihlTn:cBFOEn8T\kGk0F<^mOQZWUK5]jPJ4TL:AmlpFK8V:?p;;80
MagdRki5;m0_L2<^cVD<hLP7_o\SfOWnHj>ic?YD4\m4lQAL9;\IOd``eFe@;@DO
K5=[QWQDYjZ2=M:qU=B3EmAko\;91\c43kSQ?XKQT]ng6[]b;39k`WGYBZc@jXFD
1bI;\[9_AoD9Wld3U]f3Lm_X^>Q:nWEYE[[qCo5]ZD2$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO12P(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
Eem[BSQ:5DT^<AWH_;^[E;iLASOYJ5\Anm]FVIhD_cq1D8MZnX=>oa2XZ^gk@iO7
4mHYQXqo9lX4=2SkNDYbHT9GgRfbfRjjR_NhYIOUieI:?2C4TA`@AbQE=_>:jE>8
hIcGZkg?=oq6Ln2d6p>k98=Rj>jL]Ch7L[3RElW_Kb_R>Y@LiPlQpGagL8>i9VA6
[FDN7LP_[nQmk>66DmgKi6XqmI6Z55i=<\C^[U;VD9d`Z=^g_dqNZOoR6PpFT]L2
?pm1f@>WGLCPD<WD=7Eg]8SSVY\K[?7l7fi<Le5eN:<=A6ZcPU]R137I1eo^cRln
c[m^CRi6;3O8WXPJPdkW4Y^l^Z>0A7]MT:d<LjQgG9Y5^3QjY`H3<d7lpT?;^Hmn
7BI@f^b6:3Y[\iQV_YhlYV\onPQ=P2_a:KC8RZk7F?J9n^]G`c:PG1Ih^I5m3MYB
>oAe9a3jY5696ag:k1K3dZAJ=RTWYm_dc5<cB34GDf::5n`o]ZmpkFJj=IiX]j4O
DJNI=lTJDcnSKkRIe?Nc5o_cPYT^kY8QQ4Ea`Eod\=[0c:]_S\g?V[bJ^bgG<31D
YdkC_@K;]VnidYVWF5OSk\hS3YT4@Fc=Ugn_L7k?fX_H\YqWjGJDf6<@_PAdFbJT
J\d<^6qm>>Y<i]UMlLadifZ\I4DLf7LFkE==[lFd]TF5Ga4T\j0I\0fa_2oDJLFI
XOA9R7UdH\5UCRGBoB5]oH27GX4EX=^ZVqfOJ@DjpGD2nS4BjN5_5RVf1JCf2:DE
8CXZ4DonE2[1gj`RK4NkAZjHBi4Bd[C7gBM_Z05Zi8J\OQWDiiGNOSW?kcPU>h48
pmO8_ULPE>a4E2K1X?1V`Q^IRf\972V=YWeD?;=>][UaV1d0GhZYcQZMZ[Ui[a@=
oHf>ojDP>7=6UXmIjnCXX>NNqLie^i5m$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO12S(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
kb_T2SQH5DT^<Pj]Oa`l:A735ZF;THN13m]GVI^FOcp>?G5oF7IG;`<2K>SH6<J2
Qq;C0o;AkGWOJfZfm35IAi?5k1OM4E[KjV=Ce]1CJEEVYmE`cqS2>=n4p?9fM_BO
Gf_7gV<JkJH`TkP@=joK>i@MlVlpkgl8j]S7j2<GHBM=::;FHCSn8h>GGI=<`0pY
O]HkPcaO@e6kBf9_cZghmo2C`pO93[`3PqWF^iNoLdYDU:Nh>:=B1QRmp]2]1ASq
`T]\gZ1T]lg;_8T\[d;?<Z9XN4PNAlmGT<QFRFZk]E>SUm^;1lHWBleAD_f:]YMH
`AjfYbk5:2Pof1;1fgKbU96oaAk8OA@X5<^@P:LTI:KQa9F2=Z9CP6qGGJJ2Gg=a
KC1[8F>BHBe=MoFK]N\<GKH2[I4`d@b0\_fP2QnER_m_Y\2S\aMfkSn>2<e>OKJ]
H:c;M^k:KVY1]IR3EKGIZjiKlFghdmb__K6KWg[PUVgXB94:cp>`lgT@Mnl[7j2I
dB<CID:4;SVeGGYio7dHiY7IJ_A`;e@T2dj:9eModN_5VKVLT>>Tb\aTTYhEcVmJ
>U0B2G3o?en\9TMPP_nHiYO2<cT[cFkINiKFi:O^p:ogVa^XIc]ooh1Ta4o<Mmdj
U4<4Q=V;_2R]V4X_]nFE]cXJ5HmY2_TXn3_E6_jLE:8N2TSZ9fbnO;OV0D0Ve42q
LAEKDoqND556Gj`U_\>K_nXElE<LLRgjk;>FWiVT[KIRmc\IG23=X^;j^bkQ2QHe
_i[k5GANQk@fNKN:HEdg`TK@BhpF8>e7?FV1jQiYJ]`L[UL[37V504k<B0TAd7Jg
FDkW:_gIF<^=WHITk`[5GLD>`i2FhkfE61O7NZm:A1c1=BpkC[lPb>$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO12T(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
_:SVHSQH5DT^<JM12agm::Kdf6M;W=8nmOHnf80OpRm2O4;IFG4X28[H[=c=K>IH
Vd_k]4Sp8C8<dj0KWcAeI_>^:H=kR;KBQ[^T6n=QK;]a\hG?0_OQPdVjfXTpU^ai
iSpOfA78BOYM;Z`8QcbKXN>h`DZd1`QlJXNYlp]3NFbHLbm<6_;AmG2330maOA2j
YkJ8NL54p><?Bg[PhB0Qi]DojjFVgh9S29FgI\no4DWP1[BlLHWiM[1]:nC]8p21
ZCJLeW63OEXJ`Km78d8N4oQop?iAEZLOq42`_]dqg8Xm1S4BBn[\GX;ab;f5heWI
ZYBdG=E4^LRi2mBWZknZ=VMRAmU^F?;K`I3MT?8VgkU;g7gf6gHOem@7T:``oXQB
\0\C:WlK4L=he`SD0[LEOLiX@biXgWqVDb\\eJY1I:aWe_5hTCSN\4I]^jaZi?SF
7AJ4=`GFQR[b_ANJ9cF?K^kKjI=6hoD>M>q3BbXWgP>1Uoij=>ldb5?9N]l@VD_B
JJAV>a]CE2k]o^E=[DmgcIl\gfJ?IfYkF[dJON4GX=\_KBE;nA?ncPV?RD8Y_d<h
B3R_e5=aEUkAk;EXYn5N8jmEDSFhNp;h3P?n>;]T4e;e8TKIIhohF\fY0bknJC18
9a4Zm7lQ^So>LoS9DFR_YO6122MdO>\BU_cODQakDcN\a\aoVV7l`BF9kioh>BN4
;`QZm713;G:8C^KkR5j7<gbEpKIT1ln?[=T\hl>g>iQ\nXfaL5FE@Rc5BEL2AOKn
=0VQUdX]8gXAA35R2nA?VQeilZ`R3HUl4MLm1I7>119iE=2K5M@q4C>chJq@Lkk3
b8[>^XQ_5G`pgINBD@eDV25iDO0>>e;Za>8;8LJTi380:gVGk9<HciC^iWGoicB0
58gS9Mi`@;<[g=V[B2>^Y^<iS3`aFJ>pImNJ]RjHDQMkW3?RYKHC=iD3i4CdNEE2
ECo9N6_V?^ICKfEAEJV\T49MUoWbNfWY=eD_oZ:oKGeJ]9jjFU5cTISqnY\NL\_p
IgnjSD@GHPl05@o^<B;PjbM`>ef[PV@lE?=b6UX7PK9L9Y19Vf=_00_BQ<==U7m@
$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO13(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
A2OPCSQ:5DT^<S4h[4abd>bJWMC;NJI;mOHnfbQAqiA\e3a6NM7jEJnG=Bk:M]72
cA[Gfn^iXhMh<A4aqcnB@ARSb>YjR_X?I6DE2_TnhOYS5\jgd]RgFKGcA5464Jg_
1<iHhTbo:j8_dYCVOE`qU4\0HmqHO8PgOGDf6iijG0eX2_221n2l0F:5mMiIa`J8
a`7pfP_0k1Gn^mQ[QiJnJ@EkOeSnRfmemBeE;lp_K51d:gA1=l99N<kD?l?cA`Dc
dDR0:B2MlL_]aeK[CX]h:i2>S3qkEHXMIPdG8nPLe0Gc_JoVF3e:DqKAc_Li<q@A
:@c8q5d1^Y[hjD\f=Bi:^SCJG1j@21RDgO`f?Y53R1d^ZOGC4@9EVeil9i76\8Mn
>BG>h5E7X5OIaBH4ZFBh26ZZGT^QYMM3A[DTlF5mg8>\_A41Xa1S?`>C[^nZ7PUU
SPSFj<UBoX?qelEi<no2mhNU9ZTBDnZBha8BSm2[GC>cS``k4c@70DTf=UBJJJm?
Ecm6?Cja7R0ke<mNO=<m=Gjgd4AM22=>NMWjA@96Vk:lc`loMVZo4Z;G2FG?ng=X
]XH0aTEWm^oDo2K9L\p:ZLRbN6R]dbdgC`=nEiTd;EZ1]3K;KJJValoJPZJ8M;[m
1kaT1OhkiIa3\^1d;5I:JGK?e[2PoS^B<H0m\E8]nXkiULdRIZEEaO6S[4K5BbGG
Y;YaPMgkMJYVP3K5diJR\e>m8pJRO\=4fbd>EFXhc66K]R]n971jNnK[3Pi1T7DF
_64FjJpbeSkkVJ9FbTK\>`;hGeS5[V`>XYWEboaC8Ph:IZ\\^:6RQ:m@jVO;?3M<
7g7Rk[@blW`3MYMN:IO?IlQS?iYAkX0I;nGnD=BK8m2F0_POX\WdkkaAc9WSj^oK
91;VmbB^4_UWWqfn<4m3\l80U7Hn=XcZ0A@5`M[^B;idkddWJHD[7oU7V26c_O6k
U0OQhmn<QKVHSffIcZ0MWNeLJbY]02[Uj3e6SeL^ZOohW?XWiG`=[G7O;\N?D\EA
bKbCP2G;iEe7R=?e1K27qa2D[X?9<DTKjnlZjjeEack:e]E\d0KACO2mUd@IH]:6
eW9c?6^e>GIFA_YmR=;3Zabc[[e7WSO[8Oo4g3:PD<GI33L2MDYXA`2:Ue<6`Q<3
id5YlR8L]o`m@URf4e1Y5`Ho8A_p:V<7jiQM3nGPE?:>dgVT=lcS[AM9FPfkC2WG
:E::1nD:P>7kQYDE]GU7AoEkJeIB:YRWAeOEHIGWXZ`hMkMI28WFiI@WiK5NH25Z
\fAZ2`;8EHVfF7RR40gZD6=98BG:>W`3U6qa`SVQFQ0;aU@dSgZ2WVW99QBmHA8]
c7YPn_dK4H95^X8[Cne\Wa6=]QJ98dkj9<IaceQOAW[5H>iX?ho_]IZ6Ipj665Ta
qeH:j=E6Rd;>FP:ocjgNKoF[MWlK_GgXe\<@GM_3R:=_o[n<AooRTRiX]UJb7=gU
6e1P?L@JA1ii>c0OW;9SqZ>485fN3i`h@6OF>Q1Q;FTHDV;@kQ1fQL;A@Q7YahQH
]PD_bJNLcO4?6jVJf3;GDN:d`<7U0J8e8iA@EiYfLR8;po`:afUe0P6C:iClXAXB
W:DqCB4h]iA=?=NiL_`Al>EOZ\NiF]1maa0cD\XB4E<WY0NMhh0kk`T\5JYENaG3
VCmI7]PBof8h]f=gBAl1He`]`BepKUoVC^P$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO13P(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
QJJEASQV5DT^<071cY=RW52Y7OEk;N2mKe:LKJVqY]1d<BBlDi5lZEPHP[]fX:9X
ICU@0m=2QM3k>D=b0LZOGVL9ZJgadm6I3X=p?\73U8T2M?L:VMWi7L[2?2o]X`3P
bj\GTaaq4doIB1q\46PR[eeRjAXE06ah1Ynh1WkN3E93IgFS1I:_RX1pY08g\cn3
BhMSEfS?7C<@QWl0<ZZ]C_E=UBpV;ZV;VLOcd6MnY_TeHO1FJ9fglqebb6T:hmMA
d@YoS`c<bkNX@AlCD8efoOZPE^D^Oh2`qnIK^>F_qLTT`ZBp1`QQl7Slmm^@W<8\
BISPDO>cLI^2VoUVb1=[76JjJGLG]RLIZV4@6nJh\U7cecc31M8XIlJLFIUbjOdF
[7cP:GEhKoJ[OJ:TM1JGQ2ggc1mC4E<AlJ0W>DXEHhWOB\1Q6Hne:Wp5A@41QA\j
oWdZ\ZY_gh6QBR5mLgonQEh05WI3QbUIl_iAKMaBNW5cN6J;oOi2Kmf5X=S1KZ8H
\=3oKKkT6HQ^NSTbcBoWHMLE5=413Rk86iDO4o:GZR::3?d5LRjoR]D1R@j^[q4>
=>645VYbPlJahSJLW4`94TiKlDZ1@2jL4=Wb0g8aKl3N6f4LhUj3JiM9ihfPh>4n
B_>l0JMmHoWhH8fBNBjDTBBBi]n\HXSLn\T6Hglf4e4KBjNUk6Q[9JY<>BX6fIKE
h=e2pC889HHV1=Q2b7NG=[0C\VeBV<c<:^]hd0QeAEHAM8AN`hmILSFLEY7m2njA
MX9omCLZHOWabh^e=0IeBIQFDB1XifR8HdgMafQedB_R;cmeDHV0=Ig;hb68a\_[
7gbF>`M?n_0q?`EDFMh8LkCd[4lV4PQ;NU9;g5Wn7mPj?3ATl>`i^JGFnRi_OGEj
h[]P6e_oog1O?c4D:D:i52WEG`VYUdlmn:_lb9AJhIfVO3Kg6?`kHnoJBZZbTL=l
A0;HC`QIN8T7=hJ6TdqWDIoo_P]_D^JlA=QCe]L6SYjmh;GNAS]FQkP>N575>@b:
E0W3X>7F@\ZP7V498biW[eFF::P50aV@^dCPSX6SW?cLJSh:6XO@Q5<\:>dbhURU
[4oc4NDl[OCI;X38[lC9h?n=UqR=g<mO<M]lLDo?^T?HZ00dGa:2d`Qfo;iQf63E
F;I2cRODSC`nTcMQ`]0`p:b=DZ6NAJe^gQ0f@E6C0eLYSVi3:h@OdhYQ]nG7aTWD
m3a=RR7HMV?Q\37KPd`IQ:0V?A:IMDP7iDCXD`8Wk>a:L]ioFa52]3YMRnI^E7VH
<QVRZ2BJeaR0dHTEkDN:[d3?0DNqK?PFcSbgYT6c_MIf8dnmi3EA1MeDe<Y2e885
EQBic?YL>T^fhbc:GodBZLI3nAJ>K`2Qi4FMSIMP?hFG1]8h`0q_SEXX5pGTGY]a
?M_7J2@UQL]LfLLU:Mhkm\5g>9E:T:\W9k07NL;`?fjP2<ViCC<Thp;O^?HcHD7^
HkZG]D]I`LaRCnh:\3]\O`Wf`GT=BN@<Qa8Af=DldVQn=H9][UFM;c;c6O<BM3W_
?hVcKHWUVqDlaIe7@dLNjaoh7o;g5bS6i]MCA;Z_l6Jgoie6n;GUR6iK_MSKlh0L
LYBAL7SIWYCYk^>OC_F3jUmRLFI<TcG?lpXK4cCJ9:XUnWOLj=ajKQ_PYPQV`5VG
;6Pk=L8]3OGihCY6jogE]BZm7:2\P_FAbNU4FaQ;DX7[hAIKB=]3MfjQfpcZCHRK
c$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO13S(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
nnIHSSQ:5DT^<KbHjFc:`[g[MBZ77W28Ke:LA92p_2a5VQmehJL@VN>7j_^j<]BC
[4g_WOVFLUUc4eCYR<5nC;JkoZYP3b@m4bY[l:ZE]c4<p?4nQo;WaVH0ddc1M`@6
EBMeC8l:UhNP=46C@0;@>4=0TpA\YG``p`oQ8nJm]>If?20X?iF>5[^=2Z59I>[b
5f\K`@:i^pmm6J;HAWC20XY93VMPmH;4N5l]V2IHW<;6qg9i4=K`_UVNUKME;F<W
ldYBA@1q@QbHhf0=d0M`57p:1dn]JYpRRH^j3p^hkBIVaj>0O0LaKlkf4eT2TZce
;AUFPZFDfJmDUoKUNCA<MQg^Q?VI^1=^DQhKNh^m5_B=Jka53lm:K9URkW6f2]M^
?D6a2:>D0Jcg8j@Fj::Dn_d_^fP]gcM6_M^m\]@So0EXpZRdHSKK3lNDEoUPqT\Y
c:`:16L;Je=GeT?JS\S]@_;=OomH`iTd0FFiXXNeei:X;Y44kcGOBQHf\5?<5TU_
>RTFO?m[Em[;3i^TbLKS7WMLa_Rgj<TLB3:IK57I@Y4EM1f7ohcdH5_>^OIoll^2
jMTp?TbkaDPXCE>KN^kQ9jG0=V8_h6l[21k<JJ6EQoY;9DQT3H?;]9I6C_:cEF99
cUN:?c?SM>3BR4jSedX<TPT>7VEJ]3AAbA;I5JLQ[\n<:fSC3A[Lkc>29;BSRgmT
PX@_5^1;c6qi0Dg2gZ0QhAWGJYf6R4\O>5bleReV[=@YB5CGGT4[Dma0o@EHD@hI
HgGQQ`oZiEaP?@fck:dn4Pa`2S]m`AS_X8Sd^lTNG52_Oc7HG2S86<8?;a7YThQ]
FiGDKj^1j?jC1W1f>[Nn=qo:on_ed8`809Tki3`Te`UPOb4Co8S4J[lJ2bhJ;`fH
RPZh@X5LCnS\PecTcR[SiPRUWLf[2K@N0OcPEL``=2DMPE<UmJI2?OgmYIXJ\KUP
FLCA;\mWEZUeNP2hM8Uf9^BJCK:iF6i7qD]1bmmW?Cd0QK>OQ3C;[Zm\W3:_<78R
]aDWNfNZb3a37GO2[HT8DmIlQ2b:;OIBcDeRV5Y[E@ZD<_;i464b6F5K[XOK`bO<
lmD?Jh?>;6IKBI6=cJQ6LI1eBiJi`7S@HWg2B^kp?jL7]>Q4EM`f8[3>i3g3TY>g
:JaR:FdB:1Gc\a6e1J^a8Oc<T[Y@PP089bP8B3f_?X[lHMX0>kSm>4dMRW5j7D7h
>97W2ER>o1LbNF4?``o0n]R>VSbT3MgCki[kdMFUG9gR8nqHDd1e;DAMHR<`[@Ok
=gUjYf_QA=EjOEWU0`RGHHkT[QbHiXX;CMef3MnmWPFGVbDH>glC<dTODlCA7\Gj
mK=11qE;Q`>4q_:3`?_FGWRh5gd_H]nImF\^h=m4[6Ie0QE\;;Xp<_LUEZiEmdZV
R@BZ_9TIDJJ?:>aImSGJ@DP12UfPVoZ<BcO3jdEC>RnMTk<fFacO_]<H=h=]fh<n
4SK5=on@M2[pG^`@ecYSDEL4h@biA`V3FADGNNB=UoiPIk621`QBXn72>NnCOUKR
>PDK8M_bgo4I2f9cFnXGMSDZ7XiTE8QN9b5qhBGJD@Em:FI16Bkf2P]2gCLc61YP
WcF:9QgF\L0TkijJe7MbG=Q0^iC:4kYNK=9l]aPWUJ5ke8;=@Fhka@CBeCnqU^m5
1fD$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO13T(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
3QaVVSQH5DT^<:PYVXOnd3`Q`WD`0Vj[3FO]KPpRkZWT7bdc3dm8hL2mGSMoi2\E
PDp2NX3k5397SJbVEF[FZB1U2X7Ja@WgGYV[BG2ImZBZ:bNNEdoRMBl1<l_T1U0Q
=0mpQfEY?6q[4ecC`MJN]JIDe_OS5kEU?PCGEVaQ`=LnU6hm0H2q\FYGE2lFCU8J
O<9a1]QY6_@6hhnQej`hQmqBB9P^Xk9on`K^S^MXG:9fJ\@>mqQ5Ban[hq\CX1Y=
pJ9M490YjA:EbbUKck7Z=;MfeFoiHVJlE9\d?57hAo?W;H6Uk\@WG?=c\2Kimi^J
jJ1QjGTh:JJ5A:5^^T:H_f]R?QmW:ao\5]\SZ\<GYkbK9T0hNaL\VldJ3J>h0@n^
Y>LL5DTp0>gO<_JmYRK]e2AfF9b;2^YM^;=q91V33>C2P_7cX\n\e0]940hbRIkb
d?hA[Z;bEgG2fd9E_aE=MF6YbRKP[af9RM6Y9^:MM7bhmcO1nT<dY2Aa2j8Oc0]c
]>?jHZ@N@4CF\Kol]AK_1LId=K[P1Z\>D=bM?AL0[4qPh?UlZ;2;fDjD9`c\l5D\
0gm@@9cU?KNdm3TMhQ^@E:VL>DcIkdfoGFU80XNEXG5Pk0OYLlZPKFhb[da`GeUn
;a;F]35NH4=FmO@`I0l]7el[BOM9Qj@hhBhCVASX[?a_0njCDp1bI?8JRa2@dBKm
WRe2V\Y?<O8<W68\ABG@9NHHhZ7e]X;A^[=hH1K7L`o?K4F2QjNIT<UAlmm@2^\g
YN=afO^]9HY\BdXYkmY58gTHHZN\;]L^J7\P6?n>adk99lY0QRL51iZ9[PK?pSaA
Q5Q\84kFM:8UTaHimiF9?k6]kHPN;\nF0^iNLk9;i79CfKRZmI4d6ADZ_]ZnAg[S
jA<fo>QC`Z0BY5ZVdAfm:Ql8XWCj0?o_j9i4d_3R9L1k;I3F8>3C[[UgZan]Mj`W
A0Sa<@=qR7An9e8C4aZj4_@2]aneHR<?XUdf=h<nZY<[28NeYkOFn3Gq2a`jSXf6
TmJmiQ?54AK_PCZYi3J_NHO:8cA^WnA;`MWRNRHV1I`]ADeBEioc?L2T21\I3mm;
QZl4Uk`@G^?X2?LM0U1Q\YaETc2Kl:KkY]<bf7W[;DjgaSQimY@=O832?\c\NJqO
Cm3]O]f9G9;SU=XF39>oocSg0>9>glUKe40iHn0=O9nGLkVR8ORLQfM7]D4aO7]O
c7^8;JNL\Ra:g?h1b[[TZWJBQEnE@hR?ehJADm>BCQm`CkWP^oD8PD?dhiaP0n>0
@NIl9pN6mC6koNJ:eX;]03Q?1J;jb0?AT3;Io24B0U>aO]NcYUmdjk\VT6kd?M\N
FEeFPoN@UY1SFO7:Dgg6A?T=03W2qXJQ4a7q4MBV9IB=?>_@h3V7?3aUgTmaeZYf
bAO`4\LTO>1GXEWMUHi8;TZ62V7EaF5Ql7iRRDB8PUhcnndEKfVOKe:O6mfp01n]
>dQQ9e9a\L0Q9[9SU`=W?iH4jMg^^nD?fLFb8VLE_RO;_lG_X`i66COe>ANa>o6\
QNG@8^f43H^a89`O?BIqJnKB??H2\410gmHi\fAZ:01]G3[_jfl:]Wg?bN2@qRi2
]XONJDAEAFG`H<dYmE09e>;RS]=FN;g1FIC>ieFE7a@EJd8hG::Z`h6THdRV[FAI
af;\>U;NfcDOdDEnK9CTpl=5jRYM$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO22(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
M=_5CSQV5DT^<LmYGT^j>:=4eS`^nkIUmeSaqSETPae3iC[J^GC`mbePfqQF\16C
=7;MAR1Vd7co5d?fc8<[d[eQpBe`SnJq`d\jJSnS_PKC]9mR14OoJ?JK\:`7KLT1
bMp`N=JC`d01;M>FeIiko7C4Hdb\[g5c^6[f1q<LgRNAd^fj3<_o7P<`ZmgCebbd
_GVBpFN[Akko_XFH5^PZ\UFE[?Pi[8W`Rmk37UmqXOKRbRZ;EnkZ85>TW]Hj`:T=
;YpQdHN_[Mqg9FL>=qSU_@TJAYVi5Z3e2_BVjm1eMh?gk9OSdKmFBJ0Lg[3kTk?>
aim@Xo9N6oDfDJ5ckUSTWXOeLlo5_6^ggYC]NmgoQ<Mm62TZN7cFDm8P5HKg^MC3
j^mA9mg_pSW>J4H`iaTh5C@WXaO7^;Y\Bp1nD1Rg5De9Onga`IDT2gWhBjB9KiH8
OIi;8YVgRNNEU?;lA>VMM2oGj6VegRVWOO1KU4\bV;FI\PlYEgCS2\_TlZc`fARB
V[P;<YHcBM09fjDVFniZ;oSmp;iTiLUHOLNI1iinTjFT]7@DM20lA`oN6lW;4=Sg
W<nPfoIg8:\G:1hb49\UP`0C?;JN2hA6LgGgOhllKAZ41fj4`gmUhQ1P[:WV<ocX
6R1]=`W7`D>B3dCqX8X4a8Z5[C]E2V6bNS_6Ek90FO@BCh0@`0MBF]M@RLiTiAS0
geWG\@ka1:][YX>XXmBKi`aVYW:@gja[_[LC1Iq@l?DcAD=M>_oJog;_?E2T@`NH
7>:fN=Tg8]7UKI8En?dj4DkEh@I>X?nTj8^c^nX@Le^TTX]gCNH9:]03\CjY`E:Q
7ea_ajg38]mR5>k6hFa^7lOCVcR31p<1Y:<6eRBg7FLMq4NYKihk>5<Sc06S4XPI
jlb@UJZg`ClmnAmohH[EBnoN0EN0j9F^Q5iW@jE9<CG`54XgH]WV?>:034AA6Kl=
GaA`OgC;nkUW[EmGN61W@Q?5N`Xmc`XKn:1pHnX88h[65R6M`\X93MQOHgTb_k]_
PVfYZ;9h@S:CO6boDWS[==VRkZ:C[Y7Y`W1THB8m1`EQiJIAOXODA9j8]kgo?221
Y]GnJ;b3V0lWH[86oJhW5L;4Q_q:dWZg0HEcDQ_hRMadK1HNEj@65cfijmW7i1ZY
<T1cbg3FF9LL;?eNXj3ZFM`31eP:WTK2kW1i`[mMKPD_D\oe2po_jncWUAOQYIa;
mWNVTjBg::GZ:\OJ^_Yg2ne7DRj:I?^X]L:ohG^okBDMH:hGDDoX^MlG=2f4?B7d
Xh[`SkOO<3X<J6d:;k>gRZ0Hg7AK:iWcSkScZB3Gp];U:[[ojZiVEhW@g6`WWLTg
F6H2A<053mEGi]MCi8Of_5\aa@PB]S^fGmbWH9i22]O::G3?JHLknAVL\0g9m^=W
:WTTA]gF]0EG[cd]I91j3Te_\lhg6D>q]c8JIjnJGEI[F2edRH5;?00_@SX\K?OB
6WlHb6Ld@9]G9YchNPDSd]UcZJo7YoIZOPiD:SF^C6KelKiW=o0Sm=:?JUIK5P0j
n9Mo>6@Ab5>bPa@ZgS@30\IOBXp\Aa@jd`DeP2_c2BFHLU<BgeaaL;^__1lgI[An
6WbXZhk2\mT=^L6F?RXBE6O\BkWo`EbO0a==Na4ZL\gQ>`MTJP\FXplID;m@4X<Z
kebNkAGW9_jK^:6O^H_hI6BgUVFf0KLZV\KQ8f92gM_LDd1bF8[CRNl8dCg_<`EV
e`Z<^;b[gD25=5]CMkl:2[PgIQl6fj_^SjINb<_b^<>cq]<G:;Bo=l^jYkC:a6An
`p;@M[cD_5fB>[dmB>l@OVZb<IAmC[eT51_3\WJN8g>QS;Ya^hmZ8GlPS1Z@7BWN
G5Wj^m@543HEL^ZNQe>0DlIkSj;VR]5H@E6F7;GN;Hf\0Rle4JOgP6cS:IB:pU8a
G:lUGVP3G]]N[c`CElkfAoU8hKTmP[3`YP7]]hg8Zo]k]nR77R7mdRM78`dIc`b1
]R@ZjMeZlfZecKI\G;>kdYOHR=hTOGAoB\7IZ_>F7=Oi\Rl:;3K1f]cqc6g@<T0W
B6b;M600MQK4]gPgO2mlYGlEjGB7aFVAY:;]D`g2D@V:lUUP2Jn49DYB`d_me<ST
<16Lg;LY^Q<h;O<Oe0qoNOJJRp1b<UYf;$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO222(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
CW5lVSQ:5DT^<KBRDfe[2UcG^3SknkIUmjKAq4g:G:_BV1[mEba\^J^nY[Y2DiW`
f94LBV\@h\<i4Di6YEP`I<7cAA4NT?ST=UT1WbAqjA2haSe8dHg2VM3aSDj83546
;UTeqjM^C>bpcg^ggljDX^FHdie0O]`SZD`Dmec0W5]M_SpKTj<_6l:TYcC<QH:g
i>2Do=S=H@DAJ^c>BqiF;D4H3MCkh6EOKeaC`0MZFcTWLH^IF6?gp:6i^1ldncJL
a;\J23W7N4`Z2IU\iVJR5e450gcN1pjP65WY6Aj4:a8`X0aB9Q_oiDg6pRW13GFl
qNPD09`pM_55oToKiRobgEed6fWkGK8KDSnd]LA_OBbWhN>Zjk>XaC;;[W8\BNo>
8UO[d:AfMLe2KM\4g5WmGRZdKnk27_?\b@K>Id\PhBFWQXlF_VQGTYdPXB<Boi\J
?elVa:;6M4M;:M]Rg54IGRZdL24A=iq1]150577S\^XbWZY0cp9QW7AVZdAcm1k<
9WBhBmn1ba<NcX3PlI<MhQ2fK]Hf@:dCHMMWdg;_?1bEh==eYb9H>5fHaXM4lCQ@
ij^WHZ0TIdgkTm6mfa9M04?b5SD4HAA8In\V]>6M]ejYmOce^N9b^>[H7?M4?CQ@
ij3DTWnBpg\5oab]c[hS[3R^^ifGlH8\mC8`kOKEhWZ8N:SoF:AWe2;J4<kd:bTN
8@:`]9PgdgCZEIDX\C=AN1:<=8IM0e@R5MWHTWnFa^Z198Rf`0B4WOMU]LUDh>2R
T5_gNiP_Ag3boMD@SC=`m1:<=6G3HXbqc[a6jJe[4S0@VoNHhOQhl8_8H`3m1X[X
=2TFh1@GmKA78LmDLlm<2W3:[nTH6h?[ck2^P:fB]n8nd8C3GdcQa4c:7`E;=;4>
k2Y_cc64hKU9bHO2F9=G`>mQ3D5<\hM^cRVOI:PB]nond8C3b^_I[mpgM0iE=ZaR
>\F?EnWj0Z]lfMGAl7MAB3HWMQ?cd0TO\^0>bF8Y9VUlBI83^k]Id>XgJ3>ghb:6
AX4eUYNoKo;92UG?Z9W_TAWVMh61iF7^DUY4ciNXMZARb_]8bfV=d4hg`f7\hBV6
A62eUYNYn>DQCqR;RYGnYcidO\UF>8JSE7]EEh5O9VFEKJ\1Ag_8\XXmafCg:ke[
>Nnh3Q@?Rm]^`Zdik>`:=NcN9IFoWKKmLm?4LbZ7V4YJ<Z85KID8H5f4d3DX6LBL
?e3`XdaF8?^Xh_niA<`V47VNkIFoYKKmLmd<Ef1[p7HTh_1@AO:IQ=ELhO`9N?2N
ci9Y]o>>6WbeM5l[WSjV4?NnW`OAAhU<M`7Y_gS;H7<kdSdE:EdEJg[8:0IeW[2;
V;fF[I_h;TbWc:5I:0UA?kMh^hHGYW7<e2gNY2S>i7o35:dTQEdK@g[8:oVnUoip
iglX1=Yo<4@_OZS]CI[amM3Wm_AXOB55S6\d3lGO250TLelDh7lVfbYa1AA_4k5`
ioCX^:j4e=ZXC8`CQYhQk8AC_fDRogK]D6k5<e9_<bIE<ClR_`PAJXe^<]HeKkAS
i`:\K:Gie=QPC8`ClMK<OYpeY7lHUV1kBjCg[cd>=30U\?=1]79hJ^bIX<Y4`^83
UPDD`ellf^^f@b0=5T@kERRjd9iXPA_q1kU`UTY=l<19d6FYHZWI=\M5e2E<4=jR
bFeM6T:\Z;8dQUd=naN\>3EZQ0[kn1B=1;<Cg_MICR?XL[L]@D62kPem0cP1b699
WFIK6RG_J6F<<?g_LJfI<i1b2;H`S1_317K>`_lJCRBXL[L]KE0nnOqB2@W@lEnE
HR@bTn7nP0L@Q4XUK:>>=c]`cMhFOTH9^:UbWGS8XZ=`?\XB7>@IXa0B]XWlf86I
bmT`9If:;];oDpb6jJZWJFd[PLR6m:<Jf7:\GdHT\6@4meHj70:D_=PA;?;NaEZC
^XO]M;SW=[CUoJbENdmh3m\Tmd8XK:NM2fm7ZXgX`mM64G:jMGW;AN=EUmARF`JW
ZAVGX0H\DKbUGhb[CJOh`f\<<F8XK:Jb9Ye^qBH`4FL\8;E6QonO>\7UYjEX827S
MOflc[>`9>PYVAlfH<g@=]?EoHCj\K9RCKP>UB8F4YEF`Q7:OcX6>A=LK_]FPTB6
O\4fXl>aYENG_4C2I<50`b2f0R<f3W0B2]PX<BH`7:E5RQl@9cX6>hATUA<p;6j5
P2D8T=eNBm[B0oC4SXUPn;6X@06iMlD;j9NBj;@=oZ83l@Qg`XCb__Fo2=6k;3Gm
04NSJO<>XHjCIA:BO1Tm=RM>;i_^Ula8`2k>AbfCX:kD8T<]3aRL9S;U4=E:;Gdb
c4Y_JU@1XHjCHAlF^bp:<0J6`JahIA35>liA4X<d[j4eR6M`cH58acOfjFH[nAk@
UbcFak8Z37@cfWkOO_P:W519P;<TBU2L@S=cHKolcWHQ:F998:?UagKh\_UKESRe
Cc3oW?;6NGn8H0lLOKF:me0IP<_T2;_L@S=aSa5SnpiQnHf@MeoZR`CgcZ\YccPj
A\I6^o3IJ61k1NMQJPh678_=\hALO2c]B662IQ\KYALj?\Q]mYMc\IQTZlbgafGU
PiIEW3kQ6X2JeDJQB3ohbl>\Q5`3NP;Zg>0`lFnAIAnj6FQ3RC[c1bQYJ_bgaf<d
3@58qVL81aC?cR7W[=Z0fF1SSWncb;4C<a?R_Rbi5mnMQH1nmGeETnmCD<_b7Q?@
g3S\j1l<B4eEj?b5Cm<U5:^IigKAS01_E?U2T`cP8mn6F]?HCLM@==VT6_@W`d1m
4g2@kOlcA4E_kjb^fm;GI:^Ii?`kjLjpYLF9Qd@T=W]>E=3O@3Oh`lT;`o8LQ@hf
DcBoT[RR@;?llG6XU4nVKESPDQ=TV4[dG6QqJ0E^WVF7E;3HfSm7o^27iKbMLe1d
afMS[3OHCI0jI1h\R\_]Oi7kEH;Ld2iQZBfTJah;9JNN6CV]T:I1U5]I<1;=[VFL
klkbX3j3O<]ToO4TMQTRDe7;^GfH1TkGOBWBJGTD5JUa6gPAT:I1JABJ_IpDLk7n
`DH:fBgg]NS:j`4kK6lbmFn1?iSGPlOi8e8[O?Bh:bP8P:`Q;=bkZJ0HICD5iQKa
N>B^PajA;41h31IPER>8IkV;4:Oa<YdF8Sj4nO6=]eS>6n5PYfa^_O]R>2a7i\[a
O>IDPUBA]>3h31IFcSja6p4D2NjlZ26=Vl:HKJec;LRe<4n^Z@WZe7jKD:16`IeE
MZ1:E>ja4YDN1^0]gW\I[>4Gl8hQa]O9_I87HPI0cDjPhN:^`Bdf948KRc3Y59`Y
HYQZ;?L50i]@aa=207kIe548d\kQFkOiUA87HPgF9b8kqCmmG^8?B1?YjKhM:oo4
HhUULno=2n9baHK4mGMgbSdc_Ab3WG>X0eP2DHnhcbdglCI;<_NC6PEWeNikoSnm
<eVpg3PGNF7dDIC7R19PN<[UR6Vm;9Ok77oVkhCmQ381IX]CZ]_0]E:M;6U0kW?2
7CRhA_3aU2BY4YFb3Z;UJ65C_AMJ5ij<\Cc@mF]ld3f1iPk7`kWBiYh0Vcf`k7Q@
:\nbe_]7UA9mlY][3Z4?J65C@ld9MBpWHT03Zed3C0i?4Qb1@3J6KaD08l2XB0bl
l04fmBQQJI7[`aDBn?<qNnmWUYQ>dY0^mU0\c9AcGdX3jNhKU03J2_SN1_;U_SZL
PK97LDLDEC@XhNCamZQn5fUUb?UZ6::7?2KGIEc?PX27Z:ecHVSmS[0oQ_1dF872
>52<>^Y_EeDjo^<ePEg^gf=^bNQ2^:mV?2X7IEc?B1IJH7pCX^6\X>J3nBhL`3S_
O9_DX=6hfI\So=3\mDJi7cenQ^8Sl6Z=ooGCFCK4=O0m\MeP\=Gil2c:aE]9ejnI
:=5iCTW2020j3ZN_jUKS7dmG[TjFangoNA2Ajn24RR2d4P:3\gOiMV8CaDm9eCMI
:=5gVS92^q<o=38d_VO40D8lLT2I]PM;0=?W5gMfj3BJ6W0N<TYEM7^?8]=7g2l6
0:m=Lk?YF7<l9i4Fcl]oR9d[m^GkQXYSQTSU_KUK9VR3[k3NX[F@1@Ne8Y91lFcS
Xl2d9PT1n99lPm4[:hVo9=d[hEGkQXCj76H9q2KJ7:GGhe:RhMGeFh?Mn16>jhfU
TKXo=KJ_;21c>bJBLioQcY4b`:gleF2?YUT8@EV;if91KiWoVEbaOAXI5WeeXgJ:
nLV[jAgml31FL_VE5Xg1bTS4XHn:D8HObdeiL5VYEfZG`9Wd8EbIfAXI5EMSLNcp
ZknY8=lN5N;`Bi][A=gflh9TFAeh0=nhKmMlSCN@jK1hV_J`Nl:3cT0YHHXUf=n0
@ET3d7]UiJ8]iY58XX>l:XacW2Fo9R4lF6_13C8A]5R1BD]4Eb0Tj8m[dO0eY_9B
5EJedL?FUJkNiYe9XX>lLe6EjYpW_JJ?4PRmni:@:f4;8f?[f25:kRa9\Rcl33TV
K0=1b25:VJR?KRk:d[mBDh[AIB?WWIWUXOcFXjQE]jeO3YMG@8f<SJ\SbKiJ3ODc
Y370=M6Q^;9bcJ;DfHdhV00MI<aWZan>XQ:FXEQE]jeHIK@H1qLTJBNgYVYcPOUi
^i9A595`BA=FgmFg[;G1MI_GVFH`5i?0iERA@98T@W:]4mlJmh3?i=SH3SGn@4>V
:6Zm1EBHYljcQh4<mSWN^QXG`FQ8Gl8:5C7gQ9H?8eB;gI8faDg?3[SZo;Yn=E>V
BMZm1ERG232Wpi9P;ajeRj?:WQ]HU_DLjVg8_ciRi4KC@NEmAbXoc31LXH\dUIQU
Wmmo^]?JHK2Y?NLBiOC2Xjh=l21e_C\m1mJQ>@kSmU?5F^8D;eXT3CO5fDaVVbjm
1@ed[HCFPIaLMbL37OleXShlT215_C\m1908VD2pYB;2:;kmh?2\CBdnLTmKXS8[
NfK9ZaJO6E>6hf;1TGiN:LfopOmRI5NbVU:Rd?:?^ckKiNhRBmV_\TPUMeQoD[G0
lKd12GE<W4>G>8?;YSncG<Bi?U97SoEbjF\i1E6USbQd4ZE7I8Rq=NRLL2Mc_UTJ
RbWZO9N5TmR6JI<9:<4lUERZljgU^CDFPU1>X`QAcPNioBeaQUUfBoWal?j4@<mD
hV>_Z8[2PeIS7H\XWUea]9?^2jijc92Yk6XNnC>Gl>fj[eG:JOo4LojClC;9P<QM
hO\3Z8[2ZaJe:0p1;j4`e_1^aa_Yk[6c[oBNMS[SAg48T`EebeFSU6Q`ORLUoeG6
7AmTC;nd;56[hdaH;kFQR4J_^Rb[dOiloPTQHc8PA`n7:=3?P3I`bH1[`RlK_kkN
7eC3acYk_IKULQY1@F@\R_n_ia0ad;0l[3LQHc8]ATMkgq`mY7Z1;k\;hT9i>84o
Eo@e4g2e;2?9?Q9Z6blJ;6ckT@mn=Oe8;=Y5^Z>J]\7UJCl=hi>VEbXd0_5\JiXc
HAIDT0DEhno3in_438CJWbJbW^H3ZW?MjfO^XfiO\iO2gL==ih>JkbDdAk5B@oXc
HAbh47O[pHI;?99?16i872kRA;80XKICeeFaXDH01SOS3;63LdboDX]020G>CF_1
mAGBgK\omf5>jSb1VnbZXel=HWH\Sib^]]=04ad4:QkXDX6_PW4>OM^fH57C=8c0
@J`l?fPgJe5F6S0A8ibmXe5U8WH\SVKlWADpF_Mo<0H^90la;K\LM]IJ4DC=TKI]
\Y7=l>aQ?5g1_H=3W5J:`mBX^@G>d37=:Iof?hhWRUM8LKMh3\oahn1\A`n@Y6cP
_abWd`C8X5gBAAb3[6nV@6:oKPj1nk1U?EU7IhTbR4=C6KC83dLghn1\Li1j59q_
Nk7j^T5RlU4K<KB`S2`EhUHX\kijnWhP479kNCpK3DQcP73GRh\]NI2JIC5Hf3ZL
FkD00;WIcW?aJj2UH1LU_M^WYjdcM7:n6h]>2UiRE75N@15E^7=>2_j?\L1WkTbR
lD`\gjVdQa>:J`ROGaElZ5<JTFHIkk`00lGGhIfbE>fNe]\7^Ro><QD?\L1B5QY?
Cp[TcW:<T7f0n]oWA]9iNgaNP5JGJO8`ROWK3?Na5;JTQ;McZ=@ifanZ1AIPSR[f
T1Bldd;hIjgW801<\;k[UAXE`gaO`XS=0SS^C0_aj;;E[]^<1[eLhSJV3oWKVg96
;Zcl[?;@D1oWB6102[k[UASD1556qCA]_G_AIOVDk<PDI\m3L9ao8ma>7THZo1^m
0YRT\NX<]3ca:j8=\W5]c0b98HZ9nE=0l3hAn\PP`3]Aae`>9I:[laO[Dn87VDac
k1RfRB^gB^Cfb_2lOCaeQF5GVY_HS_=d<3KBn^P\F3QSXe`>9MIVR@dpeZ2Ui8\n
9^biXg2plho2nd5WE3U?o7J\ZE6[XYNg5O@5`dL\@cL;V^0n]^BRLN[m:]FjD8GO
`>6EI@b\QlSCkQ27fa=G50]D_5NkI[W]Qi]B6kN:AXJ<i^]c1_[l@>:m2li?:>4K
>BfERj7RRl4Sk>0ICaCA5T6:_5NkEB\T1>po4cF<\fFE[f7fSHjF6BHQLMDOZg`]
iS]DC4KZg`nR7VdEG=?P8L2;bAi=>A1e65CKRhcnm3Qe6;]K=DbhEeY:EK^VNpPg
oTdk\5@:NIMnE;`@9U9=BjY]AK]ELGLkFHRIA>NJaNn9L26\fViNnO8eoaS3:W6j
mT<glC^7j8Yd;P0dMeHNXTS]AKLU11Z2\UVI7h8@a0;N\3cfaFXfXgKF=;Q=R1Pa
MKngUR^_bE[dZb0dejHNXTf15kHIqja;oa_`MV?DR`iF7<=66lNO_3FSg@@DZh_m
5R=l\Ji9@bSiHQ_;J=:eeiZi^AUi<7cNBUn3nNPjWCMg]5eZE;LbKTFGMK5]c865
mJOP\cWnA[b;B\m@I<`K2MO53LI75j]8GdnDmN>WmdMah5eR_;LbKe[UJQTpfK_P
1TBiF^;mIE_7_[h7_XG:EJ9;04JeU0Y2a[fN9Me>^JG\4;j9U2Apm<986LdS13dE
1m7P4;lfD0JROI5Hh9>Y`MH;F<]K5MiNo07kXMIU@d\mbj9BSl2dOH>o]J989A`^
fEfBEkCP=a86[Q^L@U]]fmU4P<TB^NcDOTkW7[VC8NfUcABBHcK69HEF]j8^@A_5
fEnlEkCPc3Y<d6p69nlo`R=M]RV?Waa4H]HCji[aXAQ2Ml]eQT85A5aF6h]7VH^Q
EmL\Q?eodTV;BhOaXI10L:e2>alSWQeUE:GO]m0acGR?EfJ7bkSRAQ51N[W]N1Qi
DgTdIP<;[NV61f3NXSo0`e0[>=_SWZ;UE:GWma_E9q7TKjAl1E^Vf:UTb4oJA<62
llY=n:R\:DZIO^YXOFKP^4[Z4Z5<@83:l]ka6meEPe2;7COhk;jdhW1`mXBMK;RY
WNU=B1UD2Clc72\W\\8^ALJOMlN<Z;ASDnn_NV@?U_7DgCIhNBjnfVH`[oBM];RY
WN^Nh=;?pd1LK:Chh8h`m2@80CEd6ccgIH?k6dG\VbCcWDkR8AZmb]h:R?6n;7;c
\\XfkS9[jLP3h3bClef7X>aU>SELJ0kZV8a;C1H5XU^;g^kd122fFCP?Q_549YEj
UW=ek3H^8\PE`3?XM8f>S>a?MSELJ>6b_mmp13M`]5Hjggg;aoLBH@DE62JNYX8R
jYReF_EB4`SQm<[0V_nI14QAPBF7TTASW7K6:3KJi[9l^>4N^KfY<B39l@SB^Ioo
BC1eOU??k`:8:LOS2FQWBH[D<oBM?<La?7N]g3[bi`H09>Bg^KR=<B39GmhWS4q]
?;?_gE6l4Obb8lMA7gnb:TWQe6d=jD>oK0Vo\dILD=mOW60[kGC^GQUVd9ogVZ_m
^baU;jn`b7I^PDC=GDA`d3YmeCR4hDYO73A6[2_4Ta58E64X>b`TlfJjN15Lg[E]
IG`m;Sn`Z8ZePln=GDD`d3YC2ko:hqMAh>8P@:7G;oo?_5=h19B9[VC\@\Fb6k5N
XN4nid7KWCOijD99B]Ngl2a\:Hm:UI=dg89DjiX5Ta2]kDE`Z61R@;`\A?1OF8dT
<]2VK1Y0>LQ4hK>e\QA`@PdkahUH]MM01?QD1oXT;Ej]C^E`c41R@;P8>Y1Mq]b6
edD9NS]_NT8hAhejiPS`Vl=;9;h8[7Sa3`=U@MVLN<1K4Gl4H7HT^W9WP3hG\hbd
=FGEn`U:1c9k:GaRB;YFeaQG2dnqdd_OCbJ6JnVdi^8M=6Hp13N9GdTGh6a>]>R_
eU@jEgM<?4U?U9>3f]@nSg5S?2>R2l1GhVXdIcOC[Q\0UQ\6oQbXCP04OOg>1S4m
[QU?7kP_R4cXPh:M4dVa36fNP\g;5dlcXSmo2BA]bj:k0Ho81Ke48P@OO1a9LSU4
[XD87kP_ZZOVRWqO9m8bTYZojU8Q4LS2NZC]`JlmlH\YDCjA;U<KdmGW>^38c[6^
^:G:<TXRAg5Z[aecZC[C10=N@i4k@7>6BZn69<n1lL?V39een\OIJk6YI^3J[gSe
k0bmPT4[^ckCb<mOaL`J1coNJ4f6@Si6Uf[69<nn@?L^^q\4PD;A?JbYObC?;jiT
idO@2jd1FVNE9KFEEQIY<V?HALPPWCkRXN8LfBHf@:Q]H69[fRlMNQj4X5ceeN9O
KcfkkDa1FA<R@\QR6bbTU5gO3j0maU9K?]Sb;;DHJ\o8N>\kXQYMJEjOo3ie`^96
G>fkkDSQ[UV6qe5aeF3jFfRMe@m8QLF9if`2m?WEmC>nAm4=3bNR7WR`:0Gm1H`W
36k44Z0gk8P\UnSF<]ahh_NYX?MmBKV7m_Bej3jR8:g7l5D;:hNoBYDoZnofIdBj
I2Ue0[<Wa0<>Q=SUB]Sj\fN[B?`KeKV7m5<3go6qP3IV>f719W`lkXfpS@1hZlTi
;Bc<k03GY^m8YPjOAPenZD]Fo093NOd`mGc\I8L3kjF8aFn[4FkjAJ8L\O\c1iYN
0[^2LeJjUa>aGS[T2PIFoRah>8lFG6HVKWc^eXmEcE`YSW:f>jLZZOY^SLOBSii=
08ccGe@OUKa^GS[Th\8n7mqZmaS3mjF_CXWmo?1_GPL8]68m_m2ZGVZAE0Y=[B4F
D@QFE?iI04:_j9NLhInhNRGhf2lKN_jVXY<OBfIo`Vb;[YN<_nPiK`^4=[V=OJTL
;II4ACLkX[gMKA;4k<_:bgnZl2ShNM6V>X[FB>EoSbj;[YNlXX`j<q?QG\8W6Q:I
=?SRS<54?L[nDJ;ZUD=?CKIME`T6;E5\5<?KNS97[J67l>9V\nEU0^a\8Tg@oj2_
JbBiiBd`E2cKgASZAD5kI\]EUOV8Em@:5YjjBH^M>@f970WLmUg?S3?WWHi@Sd2h
=Bii1Qd_UVcKgA8Q6;cXp8E[VIHh>jchUB]:;`;8\k:=Qhg;_JUCkdb<cZ2VO=SE
QON@[Nn=T2>>`8]?5:niRgd9J\J:j;RLceAIgQPlHelL@0gL0@]h2WRg=fklLGeU
>NaLQTVi_XJ\R@KA7@J[S8C2TAJ`M;Y`OFA4\Qi:YelL@EC9?o6pWo0N;?S0DBV:
8l;0<[Z[ba2ZWKQ]\XWj:\[=WofC>iFD1<Gmc6cIX_m3Hh\ji?1Y2RU[<5MN^8N]
M[_ElgV?dmiMoKfeakMO]J<i\`CBB\5IUR8<0Y@i_RbSOCSkmoNQWcSf\5P0^I[i
e[k:l7ahdmiM1?nT4jpVQZ2V=JWO<4<G]MQm^^17^983ASddH3]0BfnEEl0VXdN7
9^\c>2o163Rc@RlFDFOO>ECB]k\o^[2SQQTa45njj?lnVKMj5q5NJ`9od`IeXDL1
IU>UMYhMGX7K;lb4P]g@OkdM62oWh\;?_neE4FCYBWb0<pbHVGE6qFYD<\6C$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO222P(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
e;`0\SQd5DT^<C_]XXM<<?]UaNgPAh0^U1hpok4Od]?d[_c\7Qb1L`?o6_5CYUjI
m[Xpf54PY5BB\`mZYhRnlc3<Cg7j=:kG8L4J5`h\@h=goj<R`3j=<WT_^:W=C_8L
RU;Dq;_1;D2p6h:MlVMWiO?1@@ao6h61\0]PFAc65g]=LGqKGeMn;1<[P[JAo>4k
5Zn_D8FQ_G]L]IMUSqjQ^97iV<[KYYde\375cZi915A50P[6:h0dp7dgXmcS9D]3
E8=Tn\R@`iXIkC;1:o\29lKI@abN_qJZH<6?Oj>9Be_=7k;a0imUHT@7qVWMAK10
GP:\ffYW9m[FH_L9dZcjN^X_dAWFqV^_B2KAp8GmX;Cp<_LUE9aEmQN7cnNTgU?G
<3PYb`7Wm6l<mGnh95Vh:7XfA\DLC3AH`\9?@dKQIh[L<N_V[_3MPOmHjMD10G0h
YjFXA>:7k;S93GDPb687S?QRiKImN@KLcAWQH]lJghV7<XKnN_dIPO6WjMD1T[aP
HVpIN^kon`kg7<Z]]DO5YT:j5UonRZQQB5HWa25Q4B9[@T9Fm3AK1M5Ai\XPGR5]
9_=IDhU1Pa;<oQhn^1CL<XJGS2c_][nglehOa<hhP<?Hc\aOLLU4L\N>h\I1GK1m
903ISdUPPc1<ofZn^1CP\bdohpAY1WGRPmO4\JBEN^C74g:aSK0SOZOjCBnP>m_=
Fe<PVBSII7mcAA`8U^WeW7LGj^T4YVEb;IG1iWX9JEPiH::ib9ZdCBfUeT3?caU=
FeT9akU>=iOBB]P9jkeNd^I^5aI4D1EDgjc1mWX9TGPiH:9l<5iQp[N9V:bIM6]c
=`A4F63DA>CPhP=[?ANfXC723@5F_A?2keek9EbUF04M5F425C^BWZQbT97adAm>
;Wk2[XR=dGKiQGjiRTE[cN\M=X590jZnBaOZR2Wkk<OEaRn9_^aGnbQ:N9FKT0ml
iWk7OXR=dEI`H8nqYYFiaABDAB?k=KJR9d`\f=Ta6F<\eB0:eQQ[K3@5R2@@T8oB
e8R=D:dU2MRRMG>WVK>8Cl?SiiVYfbCg0MC5?QN:eRMTRbhdGZKDH3mn4iPLO]KI
QEo;Sb]l<@>Qg29SCK8?C@XK[iaCfb[70MC5`gH>Hbq13M`]LH?gKgoaoLB[@DFc
2JNYXHdjY3TF_EB4`\Bi<H9V_nI@6QedBFCT;NgW]K6:3KJi[9l^>4N^KZP<B39l
@ZY^IooBCQeOU??k`\8:LOS2FMWBH[D<oBM?<La?7N@g3[bi`H09>Bg^KfY<B39G
mPc\4pH_DQf9XWOl`QhlKd2Z<0HYiH_0V`XbVKSTfD^=>fYE=PA@GU0^kNA:kOqb
2WRe5^0L:]?bSk:kZB8M5Tg;Me\?nCIDdBN;FAYH=@JST7POgNRTE1XPXeEk>hmb
GIj376al\RMA26M?aJ`b`4beZS@jdQEFdBkMJmR7[mQCC_31a<GIh3VXjBon>72b
ldnE7_6l\<MA26Mf2F_U9qgMeX`>fTTiMIU3l_oOLE;?WXNggj^`egm9_W;jk^F6
37n@Yo:l=8L:R[T6=S3l:BgTETDFI4D05W@:Cm<k[4FRL7:@nhWeSLI9_WREoA?Y
hgY?o[Zgn<F4@N0T0B[lKjg2cMkFiTD0LC@:Cm?VS6?PpP:Go>HFKQXRX[c;Z3R3
?=\hF=QT>dQH2HL[^Ee08NGSX6\m@UQMjNoeWlQNXZ^PN1CXjl?WC<enUJCMiLo\
8jCj\P<QMhV>_ZgfN3e=S7H\XWG`n]9?^2jidc92Yk8P1nC>Gl>fj[eG:JCoHLo\
8XZl4:bp[Mi>gBSB\XWhC:I=e2YiCGm>ASo3[`SUccOOm92F=:he6ZhRU7FP4]d\
a=?Ih_^R8>29fBn@PJ9]Q\C0iP;gAII`8<p6Y5mV?hPSJSbQWTB=h4b??h;8TCC7
e[SLoX;gYQ:\bMCDCAfE1TbRdne;;gSU`hm6K\BOo\jkn2Qe\T]hcFh=;LlSKBLa
]T^aoFgh`FB2^g82=@g8:Kc\4;C@EO3f`gF6XJfLoX?kbBNe\T]MLa=QCp\`Kg5J
YQJ>Uejhg]<5e7[fbKkn4gGOmcq>[Q<\gaU^==\8h3H`@\ok?ZZR0ElfYg44KAKJ
1Tbng1flKZbZ7YT1;FRZBgIf5oK8b^k??]Y:W>L_i44d4<jLFUTKQ2Vo`e[iB;mH
1_5:T:h<Mj85l9>j9^o84cFMHd?abam?HI]0W=`_WRBd4<j9ednnWpnj9nW<`E=Z
HFRYalU?<8KY4^a[JU[AcU7[l:78g0]]Ua]]B];SSTODF^j8CW1J\a[]`>TkGA?B
bg=6miOOgRLLQ=7W0QU_ji<Uac98JRZbEJ8Dm\Ji3P1>ME3E\eKjF83]3eTm0`2B
oG=ZUbOOgRaV>lbIq?>W@H=e5ZnNM12gP1g0iWVWQRU_B=`6\9NaBfgGY10Z_@E;
ToVfD7=Q5Di_YfD8B1A7L4\?PX8UGm8TNIfB^I6I@;_]8O86VcFOPPg5oaolPPBA
88Ren`]=QV@fKONh3iA2o4UMR;8o3m=KKIfB^OL:?9dpH0o`:Th<kAcJ6;f0;bcZ
5<DZ\JqVl4Z:b[Dl0BEBI=B9;<XFhM>aBkjAHH`=gXH8ZF0=VhDT55>GP<D@F@T<
8[aP?bW6kL;lMRgG[DYMLg_8DBWVD<H>=4H?hXJE01OGZ7jW66fMZPB3YMP6oPnR
alIO_kYLkeGlE=gB[1RMSEK8DBWKdILacpJacEbKaAS6E2_LL<alE05@<NcojDkM
Hack0Z:Oe]19PUYbFja`DHa`g_95gI?bh@F`]I7m];mG71dC5^KJc:I4me;hOBbT
QZ>8?QoORSOTn]_^j^X71JQA:hnBgDlYWF]`^H7gobfGb4dUmHKJc:\LS=2Xp7;n
Ln6ME4]ZPkP2Cc27ed3TY2lbDV7=C]nb]n5Db<HGGd<Fik[P]XcT]gSj]0n6D<Hf
m]ECnMF]8gFbBPJLE@IghDj1]D8U9Af`5H5VMCkJooJZCl7DkZ949n`\NX>eJ]Hn
c];co8FdmgSiePJLE_>bAm6q13M`]5Ujg<g\aoLBHjDJ[2J3YX8R:YBXF_EB4`mB
Y<H3V_nIVMQcdBFCT8USW]K6:3KJi[9l^>4N^aZU<B39l@ZY^IooBCQeOU??k`\8
:LOS2FMWBH[D<oBM?<La?7N@g3[bi`H09>Bg^KfY<B39Gm1cj^qQOWhc2P;CVHSd
>M`M6iQFVBB95>bM<ehR3I3i7b:@DnNN]hMR^=4VDREd1HkB5MQQ9EIYlCF<6cnj
T4JlCW9WY]^`29Wj_gVk3T?To7oQHm[=0>Y^iO[EFil;>@JK5Y[QYYDllKN<ZI7j
T4JWhK9h?pUeU\XI0d?M7^WIQIPHHgHgA;aW]`[CS8Z``L1Tg1FI=fmDdG>8[JAW
@`a?kAKPmfUU3P\Y`A9`im<ZM?1Lc457qf[TCYiP>QZf]0?OHl=HaLeOLXThQOYV
o2LPJ9<5HXUJNJb>V:72mmJ5:GbjRRm;O>d1n<CRJl?c<X4ac4oAQ2DAWUTGD5j8
Kfbg@h864JfJNCfXKkAmNO=^hH[QC9>RKfanL@C@1l[f2X4J:4o:e2DAW45kI<hp
WQfJfO5f[?Le7DhXMn<QMhKWOF>kOQ:DTH^@\`>N4^aK4SWc7CRcQ<J8h@a3kh\<
REh6l4ABZ8;GO`:NAoad0fTNUF]ilf9NU_mmW?_hQD`UeA`UZSQ>^jfX^_hd\Gd^
WIj414MEZ^2;]`HFAoQd0fTNagb_`AqmjfR1@Jo?>J5\_\?AYN;g38]YAUjCc]@_
`K>U[3l@TVfRCY8^6GVmK:koo6Fe08YDYOn=PUf=_KKgb`>nkm:Ddha\AljHi>D1
3MhFOZ=aaVEeY5PE386WFfibd6k2:o<mAo4HP;@=jJKFbLbnka:DdhaHUYdd<q3L
;3B5_2hmimbC5PH\XXF4:VkfTJUm3aP:i@35KCY`=pM2_0]`d:>Z<]EkaXIY^iZ`
TW[foIA`o_8;emQ6lW]DHR3gK8TSZDBS4gC0QnC>Gb5ac[7BSX2V\NNgR_N9cCG`
MabfL6;2ToILAD3:d0KNO`V_4oo1YdBCdLcc7jM4[mMC\HRBL82<:PFg3fN9@kG`
Ma2P340Wq8EhdEFMNJfiR675Vm50I]KSAWVEW7^XXXJ=X?GoN91N>f^8niY20UXO
Ob^b9^[LO1>f4KA4ddG4d>^GLcQ5jb;0l;V?0?Yac6jP;km];2@>R_\bL8KQHamA
9`IRZn20e8Qc23A<EdZidD^BQcQNAb;0l84^hm2pa3V=_3eY6Ln`fnXbYXW`]5NN
N[9PUfC_E6nG]MK9BCPnB>oj73DQH^ieiG8JAInjoAD1@[]]fN2EDlCg2VJ:`FS`
f[]SYJ^>WcQaYWDDi:P>D]VNBm43529hQimbi1^YadJ`Z[XOfmo5ol\Z2V`I`FS`
_cJ9HMpRD6Em1WX>V;ADad3aC]_HIc?6PbPV]6f?QFQ\C^m;kl]LX>ah_?nW?gd^
iM82MdCfX;o4a?T`]ME\kCRn@[EF=L0>PT2gb8B??P:WPc\0cloA8SWlP_[=e9dI
DZW1_GaR7Yl[aDi`9efPkQgn@UEF=L0j:f<\npSM1`WG?DJUC^m:Vhb=FO@j=?G1
?2\1836mLY@X:KII`o:5@aI<Fe7HL[kB4XoTAIC9fmBW>N4cPYnF9aJTe<QYkUPP
2VgXY98lKlTX?N<c:3D@hXnlT8^0mPdXF[KdM569;mB@0gkc;2nFmbJTe<?o6god
pORoEi?iT^i1d_M8Xc]Lf\d2GV>oGj4Enc29i4N\LiAA=BO1T9Ng8QaT9faaO0QL
k_6Mk^9cSXX2JnLLK2fJ6c<bPh@dYHXOXjH]PFN1XFa>e;Bad:TJdD:96i_Mi?XZ
146ZA^gZePXE]nL^`2fJ6VCg9L>qJ3f]A[[d3e0kF4BDF^W]cIWiQ]:k5NO]1mpZ
mb0h_gO8]MGG9W<[VYH[RQbZ7Ej<0O]W]iJDG:Zob<fOPn4a[G7hP`l0NY]]M5iK
XLB[5e0nUBhmU8T_Y`@hi]?hmqAdDbCoWDnCEo>0ieIS1eA04AMXg<lRO_]\NJ99
`0d@?_T]W^DAaP0K:Bf>IUW1DS957JC7bS?j_c8UDX:SiJdC1F:XgXVD>eHEQBF;
:DT??N3oH_DANKK@BW@[0OGQK>AO@2P7<G?BINlUj\:8O5dC1FTNMamNp?iM]>Z6
Xh:`YeaC1XiL\]YWOC]AIIhV^D3Ha2C;WZ@HDdf=8P0KCciI;FJUVJ1WJS9oJh`:
S^3_eVa3Wki3DR4T]O]meaH^^9]3TT02[3BLi7l0^nm^TX]8a<L9U`N0J?0ih1`F
6^O`YBa`XkX:KR4T]0Y_8^1q<@iK\hPcH7Ca]GHGoO1[I1YLef>YHj2a:=80h6hN
l[McQVnHhjJZ\heUQ=mSPaHLQY=Wo8bdCL[ibP7LQ^3E>YJ`ef0Uikm4AgGh=8OB
fcRBQk:VK4GdNCIdT1ZF4XnC<oNE58U1CWR]3PRlQ^DQ>YJ`FbH6E`qC[2JP1a^>
[Jg\`3@80=Nn=HTN;BL0V`i]50@6O]JL=62c^WGLI=obEV8_JFZ>_<A^1F4gkNi^
Gf3KbEB]4ScB98gY;<H\k_7:[aOZ3Sk0S6=`7J2WB9j52KWVjHaf`NjCdJjBknS^
6JG[bFH]EPFB98g:ShE7hqo]C@VbEnToYI5?A?I<HJ38h<:h`3pbU9DlLGi2?Kc]
\o=HZU49`O8EW<bdG:1BOEWLU1<]APai[KK_Qh2fMABl>JDNV\6`@95;[_1lWnAZ
ONmT2`Q16Ik8WJ2CmO1cg;_XLl5468a=kaa\QRIS=Q`W1m[Qk`6bl_l][1WlG_CY
OecT@f016IkGOeN<Mq0FiaN0c4A4AecJk1<SBKUBo3b9R18ORoSOP\];CWWQNP1L
63lJk1OJbaNGZSj1ElLFDSX6m520mjW\W=6Sm2Icl6i9>_G^l`WhQD5EbD0<oFSY
[lD;[7ePY0Om4RD^Z<0D@Z@6Dg2ZAkI\C]6g[lIcl6F9XmGgq[bZ?5`Ma01aB59j
R?Od`DQ>@mDTgdoThkQE_gWc]FD\nZ]K\51`FciQoPFOGeodbL=OR?S>`8MI\6kP
SG?D[0kSO`DkjYNnbeKcg]ZI6i[\HT<bl@AVbaoC3=ma7E?IS[E9J<SDK8M>D>kd
BG3[X0kSOn>BL1>qaWX3bBM1i0@djdZJbMejPkhXjEPC;Llbd<Beb1EiWTmB\WYD
7aGn@dZDgE5BC^BM>0Lb3SKBCmaGZG?dAcHU\RTAJEP0F8gkXkYB]E<=AAm@17J[
NTIh?f6k<8\N2j?Ca5bChSUJC_@7LGDAADRQ\RTA^Ic[d?p5TbS:ISg3hFU5He<L
hmdgR4a`cRfEd>\FgoEEnk3cDDiK7mM8NCAVnn0SXiYXgn_8O5E<PfhBR11RVH\J
aYT<CGcec<W>WF;6TX\m>JgQWDBHiReHl4=\@k0OQhBglh?56gS4P1IBCKaaVQkJ
7XV<CGciLWCgSqTg?9Ygk0g[o0XCn[a1hkmk^4_kOK28LY01ATJko;lELX2AR1nY
heI@STKmL13Nek\?n0O>h2:6C\g_\aPDh7>SjVGf1ZE>qIKo\eHl^R@0?h^:JJ_Y
:N=6JW`XB22nOHThPGj]IS7UOLi[0396SQgdEo?TqCHZ>olm1_\En9@^b3bVVNi`
\_YNC9cYMHadGhhGLRNWfEJ_XogH=d35]H?J<65:UoX8OgHD73JnATOfkPfNBg[[
Z3YYRU>SFMR4\;5j^LTDYj`2OOjUB:o<fO6bM_ChHC9JljHQF3nIA6O?=PfIEg[[
ZQ`dQ\AqElO5^hlL`ID2II[];ULKW^n5@H>]idFZBCaR>h]VP?E\\;BH4:C6m5i@
J>\G[?`c=0[cDdH?jgn3k5?MohX9PK8D^H>aeKjV`8MCF>dV3ZlTKndIOm7g`^@:
lcdiFIi7EnBWNdo^jlYoO5e_ohB:PK8DHG^YEmq_Wfb0V\H7S5<Coc;Zgo3b9`dR
jK0bFUN=\4UY9kj6eho^XZ2VVFil\2RO[jMLIg6ZR;bDZQ:n5eohFbmlY1BQMIHP
j8ZCWYd5jVe29AKH3h87K`E8K=jeS15cIGUYe:T_=8hGZ3lnBfeYFi5lYS;QMIHD
ZDZ?4qaP`kQn7<HDY9n>K5aC5:XkcRemHFhmcYGZT2g>]4l56Pdm8Fo510o0SiD0
g]PlSd^Zeo4D^dE8H2cj2m3iX=]^K?cmmELeEhEPZSG_^]lRNS^LC]o[JLARDdM0
b85l=_aaY_6DTBE\o8]j\43iHT]^K?c8`:Fnp;AFi5IXRDHB2<Z:HAb7SaP2oRX7
ijE^Y^GW96f@=1;@DD?Bn?cZF\QN8Tb><i61S^=>5n[`WG4SfCJIQaLgh<k096Xe
f;B7coW^cY73YFRCb`WcR^ZL7M9@AQh>E5FM3;@:el[[NGEBgLJjEaLQM<k09PYN
deaqJBUhIRhc<XY2T2_T:bTW_TdU_ElT^BmIOB?P>Zn;lTUIQK@MNlnT@\jiME@[
G5\D9<<fI^qBX^a8o_G0RFSgl]Mi9I4]nm5G]<K3o0P[GVBgnAaS0E[iS_E1NM=i
c;PmlKQSAAAKm5Q_CohknobI?JO8R1=H1=BW]gR1LH9H\^5V_bOBQEL8gAdBlk`H
4bDGSL?WmoFBn41YC<<k9@8j?ML8R5JH1=B=nb3o>qF8>e7@Lb1=Q\0Jj:c0leJ?
0e^lUiF@O;iGhA3fL`4[D0UMcOT3748T[0M9U>NcKYJQ1CT6JH7O4Z:<0nB?KW;b
MROlUaMn46K^SPb39AY8[j5i`e5aJhg]T0U@HY@`28F8PTE6Oh7RQe@<@LB?Al;b
MRhlWkg1p\3hUeSka_l8me9g>P@Lm:GWIK0AD2`l>];O^Hb9BBX?fJAeZ0P\K4Ba
h61ZnAJ;84cnL;?L]Z>a>jRn=@ok??8DRB0AXMCZHB6WNlfSnS>?k=6ZIeXAoObA
kBcn>me?4\P_d9?[>ZV\^7RMB@oWl?8DRfj6oY>q]bgan4MO<G_7Djf_7IQNKb0:
Um2ZCEBnfX`WZ=[@oR^_D6<=OKQ5M9?Cd=\UO6EHCnTafXJYM3n\iT?12?Kfgc8]
Ym2?oTh4ka^9J^eV?G^1\;]5SiORN<Z48ET]]AC5]Dn03XUiMc_SjTFO2?Y6gc8]
@^[IMQp?A\`C44^lRGC[Ie47;\=9R8]B\okJT?MYDJ`j<H;OA_n19AQ2@LYC0=G^
MmdH]SPR5aN<;n4Z9`i2\Q\`Q[D>aTLEn`QIop]=h1lVKg40@<Ce:WDOd1VX1KgB
2jU8_dP68LRnS;NG;Z=N\0`CBoI[cPSBc:U4?HcoU2W]GXB];=]mQSCdMbhAK0hB
2G9\n\Z3gjK5o3B];O0@QJ;<hITFkGHHCd\PVU]mG0N]@CBA@1UmUSCU1=hAK0_@
KG0lpO`EDg`J`<QKPObmh?g?I@GP911R<De[L_hd:f3<JbURHJQ?=Sl>aCPBVM=O
`gcjH8R^N[@GZCP\Je:BcHAaabW<aa12<0fX7B4S39KS@Tf7cB2[6KlgEfD3L\n8
HnQo6O4PLO@mDCO;8>:n7H29SbW<a9FnTmlpoSf;n=:N:>M=G9D]GSmhnnKYVSg9
>L`f6a=@RU[0D]VnAWBbPc?>>V`TmW>A@dClJKYRM;IdYMQRFcXf`hn4M9diZS:n
XjcYLZD6UUfUR:HHKQ_PXlF1LGDDS80f1eaCoBYQP;kPYo:>Dcl``fdDM9di4<`H
RSp]Y]4>=N>BCBD]Nc=LI;k?;6B7>0n;6Z89G`XjmJFg@:GfJGa0RG3aYf>peCQe
AdH3cXEh`[::[34N]L=_Kanf694lMFTYn6RR`8A>YOH?dlL9oJ7D7B7VZ^DD3akm
n?Q_i1BTgKoYOn:l0Hk9:aPFAoQhFdOnW[nj:ek8@aImPkJI499Qb\BN^L6feJ34
`?]3iWF>ZKQcOAaU0Hk9k1Q_eSpS[cBU7QIMFEPHYB\0mPjm<:joHc@bK4:MmD<7
oBmM<^IF_ZY@P^g]6i45UY>]MmC8VZE?LO`\c1e][0HDPEOF1K@lHcIE5@h:2gQB
hcLO^X=^5cb82c8J82;XoDj^Fe1SC6OPL@U\9?Am[5NDka0F1K@XFn@M3p_?[7_[
keLOBQU]@Yn0_XfBaB4g[YWCj`Pja9LT4m^h[Y2_HaZ]OYQYRQn6jHPFXQn^lXb7
k9Qk57<BfelYWF]HnUcgICfGb4dC5^K=]H94:9;hOBbPdh>8?QoORSOTn]_WjZX7
1JQABhnBgDl?Z6]HnU3P`3KmqXPRXI\=]BJhkHSZoiA]7FB<o>F5PLUGc<cnoJM0
6aO1F^gV83]PJUeECj=M[2j0K@oGc_W>VidDg@Qj98GeYYXh1_F`MN>0YEee[A9U
j7<0hNk[W@0^9=MBF>IJ[k\7GX[;8IWfViJhg_Qij8eN]YXh106U@LjqZWMS=@HM
Hkh_gl7iPmTJii=?W?1eo3AVPB9<Q]PJZfo\OCi>_f_IHMZCQ]C<7Wbj=71KkFXl
4AmHJC5P\<AODBCBE?56D4[hf]Z[8:;]Dgo^@<l<^6Bl\>UUS5;nWnn>ZFLN`FIb
4i>H^C01\L_lDBCBChN<8=q@PF_S48aRegAh1Gb<jgpB8?c^m@T6MGG?]U[DXPUa
kX3Ym17YSM7iD828@CiXh2klbgcX25O>d=;GH^3;N>U2l0Z4>2@`<FQ9GfPoNOi0
Zk=Rmn@D@k;dA_`5GA=2C2Inlf?J=E9>=WogeF6Rn=?BSgdh>R8`<PYcGdgoCdO0
Zk=VGI3OaqVIaDhU[XBn[5JC\lAl<@B1Sn9j4DTAffUVKie@IX89d8mH4H\Td^ea
hiLPBYk2hM;PLKWeNimE:4WY9>kbG]6AJU:o=d?HpQX8RZ^qBHP?S:7$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO222S(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
d@mj0SQV5DT^<oRbTlWAe@JXH[gPAh0^<1`pHAlVFN`FoF0i>g94F17h`dDQ0nDd
\mAo[N2X@Xm`8B7mQiefOoLp7;ZchLYCm7Zci2]82J2mZBEc6G`HK7Gql;3mNcqE
KbjB@=A1KAdeADe\4\LA>;?XajVAFBoClp0WCV9i5h7P@UmEAebGIJ<;j9<Y]@om
6S9<qS`eh3_oM=9CXYRid<H6n:\jNfa1@bjf_M?j48gU:S46`065ihk;Vk5LD8HG
Zp[gR7>A0M5eGEQYJ[eJOQo4Q5E?<hWUKG:Tql9_nXRUj`TK=4gPi;DdYK3i1l3K
W@\XdJRHbe4aIq@3`2JQk41eTbo_T^d:iU3[b<>WqcKjR6UOpEPA7>apXHF0\Q2b
0Ci>YigC?GWFBm4]l0:5gSg:A`7`c04n5f^;kjmJ_SC8\d;FF1Y]^k^CXB9lcobK
OgZWmFjbY;3<2bH<LSHg6FMdV`^C=;UO4@?iS2kA?Co6Qo]\RXP9Ck``X]fTFoKE
Og9WmFjbNQNMHNpcF9f8Xdfn8jN]9ON18KUGK_FKZSVePJYb9F_]bM0^=k;m\j\[
1YQ`d@>C[iOa?LmcE>fj]Dddnk6nEBNbo6D8QHgX[2FD>;@S9Dn\EBWWWQ40P^oY
`9_bb?gli4ji?E^cFZ1c]Njdng6nEBN;I<Ba6qI:0B6Za5MHkj8Di>Gaf:SiXZjS
JJ\GW96fX=B;W[jN?0aTVaJF^T;Y>fOCKleMOFI8mlaRDN93B1g0_D8gnm1Yb6NS
Lc0AUcVfFO=6iF16LW8lTL^1WW3K5NUeW]EM`MICS05R6i93KSg0_D\\X:I=q]TP
h_WQM_dO1jEm;I8]PE2OhFGomI^E4YME><h1A8fOYRl7LF9@Q\G@`ebBp=RP7==7
:MLb347>gkQHPXia4:bFg_=^W_`g;nT3ER=FM1J^Dc7_3Y3X_kndkSTmg=^jmnVi
im3eST4oVRQF?MA=mcbmeKN_Za`l^;S=H1gAL6b:cn[ikNin2U`aCVTCg=GcjMVH
Jm37ST4oVoEl@[Pp]:lEC4BHHJ>CB^1f16dQM9BDV>B5jJnGH01G\=lNW_;Mj7_a
cWDdZM;5dJ72nj4J]2CcEW=4CFe@aUSLO8BhCM4;mO8i3XoXY0A@md<lMihB?oUb
nhABFBc1Qe8^Nj<T]G>00WUgCF`@aUSLP[ZWllqdQQaZ?F1T9PWlVZFk4L>MP[4c
kb7QHmX]^jUU>0RRM=8Ha6LZ9Z7>3ZP8cPQB:b]dBLa[llDhJFN^>:AV5S_j<:i`
ClV6]_e=^]nnPhEEQ@]4_gAYLnGkBTKCGm6A:XCdMCZ4l;DhJ1N^>:A58X1RRq:G
KX=7OQkLFLZX=KlZY`S<Uo\7Re8cm:E<Q4li3=oe<gfCDRD2G9`KNO:n6SY^a5:i
:SNgoYJZ9_AC5RInVbKWi5OoWk^R9Ue<0QF1f?<M_@aXdc[\:32DhHSNfjM^ZH:V
TG_g;YJZh2AC5R3f=jBdqlbOX0>``A^DbX3QQjE@=B[Cl`3:fWnROF\X\Jf2P19g
_XGPV`4GEfG3D2\VZV_bmlnaI1L^mo[JLA;Cbh0be5l=_aaY_6DTBE\o8]j\43iH
T]7[d_m4DLeEhEPL<G_^]lRNS^LC]o[Z9A;Cb2aOD81pZ=fZYhCK6:IX?ZYH;=1<
lXn[\[<d<GXgNM@4QQ@M::6M\ZaVEFo\LbmFbEH\i@8eZj37j:fV`AgT=5?Hg`29
ZeiGNJ::`X<OSMRhlUmO^fUo[3B1\oEh0V:=7fFc`@3fZR6LH:TL`ANm=5?HRF:Q
>7pA5\fhXk1ja1;5XMNcB`H[VLK;h:YH1ENAZ2D813W7WV8]MR@nk1C=kB9K`1nG
b0\AQefn4;350<:VS91PkcF96qXb9?9@F[CU=8=ANbkMYhc90TkgRFo2be<C0<^M
G4Bo9Cd8lq\mPJ3Ud6>Zd9FcBGk>YAJMVP9P0D:lJon<c27X@IDX67QlWIN_MO0J
M>fe2E<?fQ\PGL05\DEEBQdYFZ?g]SkN\hCKeh?6mA\<87De:lm3g`3PVLOo7V;o
6CLY[_e?ic\fjR>5@?EV[ZdYFZ=UCo76q9<<<JAWh\I@=PgdP>7fRj:I?bR]L]oG
jTTB:h_X964HlnHMh7`ogGQ:Z:ZOS<cM:9ZgH8g8E_N@9JJ6?37Uk1;55ef@D;cR
BiTB98hE8ObIj4Zjci7I9i767KaD=KcE19[\EUg=4_^jZJJ6?SH4lKSpX5UflSHI
23Uo<B0SfE2D9D5WP10GULFoc4=CT45k;K\L5cId8[10I3M5B`l?k`NFXS=7@An<
[0n?@FhSWPF1nk1U?E67IhTbR4=C6KC83doghH7Uc`neY6cP_aKmd`C8X54ZAAb3
[6H5@FhSbgdgEUpYUO[_mE`O\jlghY]3]Fk`2iHcJCh=CD5n:^]4cE[T\^?iS3M^
T`j>i;HG?hLXC>hYcY>Roa1HV\7Diem>:0jmh\Q;lBR16Zd;:^jHb:?4\7iRcT5D
5fRUlL<VUlABC16YQ[Kaoc1Hmh7DiemNCG>inqZ?a5Q:;BQM[lmj4TTkD;CIMWVb
:[J@`7=l0=C>RU;a[UQiJORd`P09l=l<eAo\D]Zdl7BaPnBYQ4<k3afF[BdfJdfE
6TBR_ZclfGck_S2O;_ATAgNa0M6\46Q7WQ3\LQZ7H_QaOcB4hV<k3aRY8X7Bp_^@
Ff?QI1gAYJPA3HHA3cHblDCQV1a`FgY^Y]b1d?ghdmJBVS0`6;U@b2;[fWCdC_FA
K4Xdj<]3BKREgV`oSK:GieJk^C^Q8\YhQk8AC_DDoogK]D6k5<e9_<3JG<ClR_`C
aJXe^<WHeKREgNX3hkcplHoL`6_>7X`g>1a?Y6UGGa\7>N<1RH@X@IPH1@JcKQO5
egMcWocUId`20X>mdaYMlWKkWXaHaTQCIBDXH?BX5jZ4ZX<X<Gc7_IU`N;j5aW^S
AP=IhjU`9h^[D2om8a=Pl8C9YX\0aJ^@IBDXK[F;WXpbIkC`f<NDG6^PRTb5KFFC
iH3:e`88EW[6;]4moA>SAH5SAhV8IVkVDAbU7H;@WZoOci_Z4kfjM@[dWa7hJ7cH
@2kcANN<EcZS1MUVo6hV5c^7eO3A`C<MB:@fK2F_oOnmcPXZeP@`MoBdJl2hJ7cH
CK@:CqV5RUBmMGDH?Q5J3O2lSAH_n2P5F1m[ZYGESZ`EjQoFROB791XiYMG>QhoN
;n>Q;nEJqenaafk?fooE9501Z5a1Yl]98b<MPBa1ADD>M`KAY71cmkcXhF3e3V0K
j56J^9^kHe:X9XM[f36IKIPXH3f]eTg[:A<LimdYXTDd=Sk^^k;Go_Tj@R6b0?<7
eH7>UF^aCejYg]Mb236okIPXHQ08J>Wqm]8WJ1g2bRAlfK]m\\P3TU^4Ba2KLA0^
fT<7RWY1EUAXB=l48QY6=^gFDD9MTnY5mXd]84CcIKi\EbhROg1gP?peX:T0_k@_
1YEUD[<L;A[;jQfa`G9kNPYAW\06B\QomNQ]@T4QP4oEGLU3`EETXQlL3>>E]<3d
]aHNBNDdHdG<j>df`f9ld@DPnUIPZaD>YNT>BXGhbDSj;h2bRUD4HOne=`2T]7Dd
XYoWBR\dHGb<j>dFXaV40q8AN0Lm4DkH<UUQY9`AUIoQDBX9A\nC1F`8hKm<^3Pg
9@X11VZh_QeA^7V@V^DAmUhob59HcRnNYKSE7lRHkd]lM]`N86SH?fY5FWG<m6Wj
Km=4]Ro\`2kIo\08cKHM>lcoKV9oTM_NM_SE^=RHkdG1OnkOp[B5KlTVjo>UbYJ9
ek2@TDSdj:nR;bZ=ZIg`\L6dk4P_2FL295An0o40NEielGK`;1_7IBjaFGg1:B8j
CMn6:N7nVEmYNBh[DnCPLk6]KH?C<8iIhZmkmhL;7FLAcHHeR2_OZBXgn9g;6B8f
UMn6:6edfO[pJ=\8GT`VWYKCJ84E2kKE8VSn1bhTk5=dEGQ7YZIIXI<dN7q;2:2?
e5=o3T:;SCef52PF;e5A30k8VAfnMJeTUob=;AdDg5n1?OC<JY5B06\N0To8c@^3
AEm?N;0`hhJ`T715kZP;NV7V`KY59UYKU:?\3^b@8@BM>B1k6UiZO9SVQIOHc?l3
]5HDNK_`hF]`T71V89X>mq8c[]jAolDfl8P[R=De4QKZ00nRnJE<ABVDaAlCGU8g
XGMc3_F:EILVF_CoBeHfG4^h0j`b<206G1MB>J\CE;>bC?U@OF7EhmU2QGACjUV7
D4?dgDCBJCh[j`CS3:ji4GSh;=`g4>l6LGMBKK\CE;_W;dJ]q;e>oM72m6N^^jFP
Fc7;LK:5NWjYHYX__KLPUeVCmV2dWUiTWI^h>hn7Dk`Z\IfkRHo@^H9[Oe_3Iaa1
DQJbCI9k@alLPo_aS37e;8VBnZdnTN5?<K98^MXBKRbL[@?[4Uo`nHB?WU_RDaae
<QJbC48R00dpN>mK=8Fa`S:\W:^@?W3H6[LYkHRE\heRA]bKfjKaPoM_[_5aJC<f
`JWJF:M]M8I>N5W;B<6E@7\3IT857hFLW9[S]G4`5K>P]]I40h9n>cX]J?k6TY54
^=K6JX>2=80cNSSJj<EC@7m>IT85QUIU;TqMZMc5KFCd28`OE0KA9d8qoZ7gRUIX
9?>Nchi@L^YN\kG>T\<XVd3l>iMH?DB=1j@3f`<_eAP6=fhCko5X=>`T`6e891?_
::37aTM7h8?4SN=`j7X3EjE1<1;[;DQ@U_0C20VGNMA=RKH=lEG?1iSAj6VT92be
7:D2aTV@h8?4bEO78KqjehT@<\h[1TbCD:C_KDY71cmKoXlb3BH:OSDK1SI0E2co
9WUX`]0@bY6gKfFH0I;j5B0LLiLS^5AJ38V\JLY>A6_\o`jT:5F_O?5BX<VnHQc1
1[26dX9Z[FF`O?Xg0VBj3U=MLKGS^JlJ38VQk>n7cqSG93LDe?G2L8`M[>L<U439
5@hlgA??4fN?=lDdeM`cY<j1\FUE:O63[0B0cP^d>gS^kSUiD>WEM@IPV1l=QgNI
qP7]G265mlFQj\5[`UI_6dj2Dg`NO8P0R;n0aiMa6A@lTCX_JB2=`eG3?CGiFe[`
OSX=`B2]^lo6:Q@bkR<bPG>H[cJSXmLgYP^1=7MKS1nAG44B7j=N9mHaRggmdZ3=
G`XY<BjC_6o[XQJ`:R<bP4mH;;dqliHE?4f8A3N?9Q<P0E@VBcX@g[R_Q?N3hb[_
LkD<WHHE^2T6ab[\ROD:B=AZo[;Uk_G[Zk<f61cW3U[TH>H`EN=3I[G[o><\\1Eb
NaYV6HHnn68Q2bfO4:\NKj@L\CGNlW6TUkIm6@NI>Ui`H<2^EN=3fK?^2^qhEgHi
;Ea79lIi9c`d_C`nbEc3Afol_7WmAmhH?Z1NPfISLdCH`YY9`=gMlkMWlj<<KPE=
>7T<;A0:Qe7X=A<Z@Z6]Yc:JdFndn1j>?FlF]UjQ_8;e]E2X]WX2ao2I8a=iK=M=
Yb91;c0:]QcX=A<;gNkO9pL0J9@fL4N98L29]Q3F\9^1TN53^^BOAX8kEKeTFQ\8
5cUHAdZ3Gf7=f<iA@7USU`i]@JXmc^jo5:_Jn?RTN`ka;oE;OfjD4nMA<imTFC2d
ClJ;0adW_=JK8oXeF@DY>17]m6X1kn?oUH_<RHRTN`O<<NIepc:?e1cJOI4Wf`T^
X<6qWT15aZEIbFo2_jBOCJ=l7_UeBIlW5b>VOlM8H9[QL:?ZjoHAVA=^H@A<]XE<
1jWbBlk[R[R`K\`2dCC4gmoo``n`\fI9O:6XW@hVE95[ObC3OIncmdmUY8MJi;DZ
YP[]Nlb9R<6Yk\32d_Rngmoo1P>O05qmb>jB[WIZiBTfnR1W:SbII8KQKPh7noM^
=IF_P8LDR:E7i?43^?6V;S>_cC1l=Ui5?1:VKBX=Nk[N<a[k>DE8D1i_f27Bo^]_
Na5=P2_CSIToM]QZHR4o9DgS:79]gQ]_?hNVFGaXNmiNY16k>DEojfXQjqQDm2KW
?<;CF37=_0NoQm2\><DKTlCc\a3oOK5O_LEKo6>12AChk]X_d9OTe3=`V9FYmYX<
T;84;:oQ_60:R>3KTWRX4MBD>llfc9IOKdcPEo4d8T53=UA3180_UaF\\aAY:eX[
?Y@4=DobV50:R>l5fl]lp?=E9[C[_0o@6F6QA]8om5dY3WV^U20BQedlbCmX^VPh
6U3Ie4F@>@FMl[1TbEd>>?5U4bAdG\oafTPBHRO?WBX<VnUQ=11[26dX9Z[FF`9b
og0VBj3U=MLKGS9JaJdMV?J5>>A6_\SW^TPBHH<0`:YqTjQ]RRVR]G[TR5Ba_hK8
5=XHZS4=<\0:jC47c1XLTolm0=5R;BjP]ROnE?XQ=lb`2>Jd<3Y3hiRHnX7HT>B1
_FTIGjZ<_C=?S=aei1On`USePB16LA]@5[5D:oe1IMEd_>F[<C32Fi_In4SUT>B1
U<_moYpHg5E=>5LoGMU8Fkai<Ye\:4Tbeo^^lNc2_MFF3bg=JZPG=]jfZ<Nj_c8]
KZ>KjZ9Zd:A_EPRbO]BM8JCi\TL^EdjMbqUD2>NY8S:lF<S8jGUTWcP=k8g_M2NU
iZXRg3n@n:>17Cb^<hc\okI9[3XJ7kVEQl070JlVfBOdk`Xej:NTbXRFcBL_^joF
XSY3lKmD`iN_7XkI>I41>4LD2J]TPM3?j`U6SV1VC_OgdYDe;mNTmXRFcB_Uo@og
qS68Z?4EecAJNV7m61j6RbbW0f]8769=O8eG`OonHOS48\;n0hZgo9ASl[AlTX7:
cPX=J^mBS>JgVeh3SFGNP]S\f8]9CLiK;]MX[4`IRU5UNJcG`Q6HN3;m\F9^jNN;
GSQmb:m6f>Qo2Ah]JFGUn]S\fhU=WJPqZMdh7^[C<>TcSm;OfOm45TnAY@[FOB[]
pg6Yj:m0QkH>>^Q8OH@58iU;<nnPGM94hHH?CTi0B7Sf@PMa]6hhXeSI>TL?FQfm
IdlDUMPj_W`V9C^]S51im=4cQ0\=ZS_nBP6MOli0O7KUON><\4[EPYR>dkP8m4aT
\>lcJMN\Xb`KOC^Ok51imOe4WOEq^8@l;5iI4hU[:BP9HJ9o0:E2DANMf=7j5gHC
2I3bV\;RL3a7N85X4SaBWYC>3<R^OVk:57j0Dc7WVHUK>FkM7fSPWANmVX8en3YT
Dil]GM;39Y\nO8Hk;li277BW7lT\^VK?O7HdD^LGgHTF>FRM7fSPmQL5?KpdH^D5
b5Pko2`l^ZSiOQWDbn5lM=[@6n[KjWJg5mhd4:oAQJ>e_fPDK]Pf>VZOn27FJnmJ
<\XKX2nbDHP<A5bhHo7WM;CR]?DEAO`<G1RSML4n;;OO_4Ym6e1diF;PTZYdfZcV
<X[KY28NDZ]<AGbhHo7XHM`[1qI8Oa>YC?Og@>EfRYDKIaO2jBM8;k5=a7ocbiOF
dS1`U<V_W29;d38Tjbmd=EUHCNj:Ta73[KoBKN]A9?MgW?SM`dg8?MV3EMG0nO8C
gZdoOlPBA^iP8Y\NgCjCgRXKk\IFKhI3e>ok`9NA[?Mg[2SM`dJ0RDb^pIMD;dd2
Z^L7Hf1XlNC43S8IoAGG>ol_G096HF;m3^dNnP7O;<c:BWe27KUb6mZ6i7O__oP]
^k=fQ2[?:8CRlehkF=GKWSEJZ3o97NS6GHYNeS5@jl4\6876XaO6Wa1N\IKAE5PE
Nk]77W[598C^>ehkFd]NeVJqAK`1UPgf0n6kUX\8HT@JA9gScA8D[olSRRkdj>56
ePa6biQFjRWj=jRMl]Q\=M0E;4^fYEOB^QgI7TgR1U[^[cliHA=lQUePoN0V6F7>
YAZbl?4HiS<M3]3Mb[<mh@>MAEaYGE2X^>9^NTAC1UK3[cliM>Z[Gcq8lF>B0S>=
XhSQ`[UCOOOoa8SWUoPGg5j=d<=OIMQBNioeoWf`B3cX3Q@3=YZ`m=;A]DMcWbV;
D>EFj8G0mXU1GKR3Un6`KdZ5ibOfG4GJDVo<]Do^;_j<Mj`M_`;eYO883NCnWKW;
BhUoj>K0mMU1GKRSD=@OQp;J==]>QcQGc<c5J;Mocmk;jph]:Pj_^?8AU`<XGc:W
jDmD6W[F:hW=a6>TMVMY40>ZVK323C=QAJeKlQh2Il=OPbTaBnlN5Ag08VA`4MfS
<Qf9b9dIn?JOq_W1mR6CEh3kjnQBC0EikFRQA[C<kk:N<;jPNZIm[=2KXi2QNJF?
664LH<DZIZonGbgGRkhl[LlB3?T@8R3[Eo1E^iCG4F89CDXh1FC<JjK<4aU[_7FC
DZZJUen3[_Tf:_\j6ch@DLNkL@Te]RSMho1E^Q2A8\BpK5Vd=MFP;gWBLdH4f7li
MK35_Pj_7YS@h_bBV\c_oRj<X=L;IRQSVIC6XW`C3VRDVhJ5_O1EM8LO60mHm8IL
JoB59PAid6\kOTMZb7Y<2SI3`WSoJ`^:G0e>1OJ9GDKiKB[@SOXZMU0O909lmgKQ
JoB5BZDOClp\UcX;WMeh@FjB@CNc15n5l=YcKiTD>R<Y]b9B2]:V0nfc>\J`@@_0
KELc<2[hNI]YOd4`g4ndbEmHZMk1W`5_NkN:KG?]jMP3QcA^JK6]oB;Cm9AFYNB0
CnO^e]>VCHf\77ZFgEldbRd3ZRV1jo4_NkN^<4OQcqE@9oJcmBG;==M[IaHfV_:e
\PQG>hJgENL8oGXMdB7mkUGJ@kJR12l[RoB:NSiddJ3ed;go>COIZRP_2^6K7Mgi
]YhgPV2E0@6ITaKMNBTGRN;QVg=dRf?H0TB5FUjG?f?eW6g\=R_IN1PUgi6K7M@<
?cPJqUlhC0da7eRIc;YFKSQDLSH8Ehl^SfkO4B8jMiCEW_OmVRUj_9[=ChgOTMV9
Xi:<c0OLkm^Tlo^:ZQ9_PKQ;Mka27alCa9DE2IGiA_T[^jVmUCXn7bA4PQaZG[fn
03<m^Uc]I]^]AoeS`89ZPK7_Qka27M2VoneqVL@JOk]^n:TC^\?R`Th@Q?iNhAkI
HI4[AK5BlYqgINBD@N6VoaQ\FKe]B[fmIEe6V3Tc^OGU@:lTD2bHPE\4`iY0F0<M
ULX^1d\=HlGSo^He2<dY\d8SRVoEBFCM5?n6VAF>95V2CDIRaP[]89bJNmL3`@JR
EVlAB>Pl;_:gmYMB2]eYQaQ;RBgEi1DM5?n<od>9Gq8BI91h;1VBQlYeBN5;8Xb8
=0M;=0^AYBRgZnfb0>R@T[DEIQHLNkC2U;Mili0E2Qc2MhWCaUfGD^C8PoeU=Sk^
Vf6;V7Qj]j;L_QL`WZAVTPlVXTJY<f]<4e71Co_j^I81Q\VC?>fCQ3N89ceSiWk^
Vf_J9ck?q5E]SMNM>AS=VoW?k>9_XIXV4A2@Nc]58\@g?<WLd:HVJIea_h`4iCi5
j>@bC5U7:l5a7T<`;[P=@gGKV451j]T]dN2CJILXA4Y4LPCB2T`4kI>cHT5bQ@go
5[>Uf]OTo5Tomb<:h[j=^UGMf44A;]T]d>U25J[p3OXbKhN^8Fi]LMSPp>4gM1c2
gTPc;Y66iifMF[cjnZP9jdXb^Rjak73g4J=E0=H?C;[\nVfUF5A27LGk6no;l]YS
_DoSW3Y]HP;:XH9PQ]PeK>7[5N_jDJ1jgO:cNX83DS<cPmjKlRUOG2F7D>GdEAYG
@DXY=iYZ3P`TnH9PQV^Lom=qKYgm[QBk][[0[X7\WV:YV0X\C<6>^4R9;C4NAl8H
`bmMd=Wi7>U5B5a6CjE3K]XXU?7Yj9oX^QblcE[4M<`2^R4dhEJgobp6ij\Coq\L
CP^GL$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO222T(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
4NY]cSQd5DT^<RlRoYU4PC_76Q6QdD@m?mF=PY<mX\i??h46p=ldOUmdADP[DD<c
<X2DZD]I=M1[A@UZUenAj;]5l>E;1W:EJ_gDPdgH<qno5Yi2YR<f3W[9bT>Y^6p4
[;2i2qlbDlN4Ol[gGenG<S`<j?NM[A:Sc]hBN7Glq4OG_\^E^5L61;0fSbS][16b
nL2V56ZQX@0qPSHT<Q`>f^7FXSG=E1QW;iXd1XfnT`2E_Wq[:4igjhRG=@4U0H47
d3b[9VoFY8bddeWB6:]=]:SqVdV`eDB>]nDeK^2<A?K3=R<nXBjLIU4H0DIl1Z4W
>:QPXg:Xi\4em\aqLfkBSA2P\`f:4V4V3BdB_YBkLDpTChHXBaqLjNHX1pK9cLKF
gY2FVS=MI\M1imS>[OG?NCZ3oUek3J>MhNH7m99B\eQ;AJMmE0Ej>H2_kgT<dY[m
37GaNNYOMe0Kh^ZYlE>6ZE;GlnVi\aeM02E1eD=@O8DbInnEY6`UU7Im_Yk<85[^
kHWan0YOfY0Kh^VED=51p`IYhoMLDVcYe@IOoFn=]X`ELo7D@Tg=AY2iIF>4?AVe
YDHl4hNM><GFkH`Z=A?YoKMH]:7<1MJ6Q1T5S78j]iC^3V[HI20CIU]<84>==I;@
B_oMkB=U[GeeCOh2MldG3jMm^:l==DJbe1T\U78j]g^=X<BpAYY?U_WbYY3:e3:0
3VZRD_P0RAQ?7aHRjXEGk^oY<[HaWSKWnPeMcLdT3nFf4VQR>719AR=iEJ35m1nE
@TLbNXid`<=b510GjMC11^oYFd=a`LOZO7f6TV\AB71G=dE<R7IZA8b?LJE5m18b
@TLbcS2VJKq?SfJKQnHPEF3Yfg3:a6V9GQm6ImC:Ie\]XXSM30kZdf];l=JdcHc0
@fR>AE;Pi]]Ma2@NA=CMEW_<nogi[1`[Cd>G_2g>J=^]EY]53E5Oll0>dW:_o\Gk
a0l`M?mm>mM2aP^NQFjHE4S<n\\i[1`K3CE[6pfL8Hf9YBc7l0M54@oD`H[G`d7B
[D]N5im6:R_Bl>id]CD`SfFYNd2^S\I9]K?eLEWJ6Wf4FWGiXikam_9][i`caZ>B
=h`O>ec27^HB0A5:RhFZ55BkG??J7dL;gmjL1:mJLWfKnC5idYka^n9][i]IDJH@
pU_@ECmQ;MFIG2geRI=>O5R9YF:KR:J8N>CJCC`kLGEKf\Hh8V?I;3X[8iS;Tp?Q
ZV\O^;0?Y:2MZJjG_UZon=_>R65cPeUFN[@OYG_4hQe1H8n?dRmc[?SYU7cfJk<I
bIdng^cE^_3O97N5[UEYNOS5@jlB7m876XaOCGa1N\IOA85PENk]a:W[598ZR\eI
l0dGKWSEJZ3O2jN5[UIAW_=aqOd876NIM<5^I`o>H_[DXY1\2EDUdXc:3f[G8fZi
kUI\Uo2CfQ?WBmoc>oS0b@Qg5Y[C^V;McOPJ0LM8f2SaN7:Vo@dZ:eO<N78lkTZH
=g\RBW6BnTnk3gH<VJlmMIj]3H[7eVh1H8P2PLMgR2SaNC7BIjBp5\2f=So[N=[G
>G_k[giOBi\3g0PWLlbKE_=me<TJ[eACQg2<32jA?P3KlK2dijoKn8jWe1Rin]=H
]ZBgfeRoWXR1N3kZ2j0UUCA1@<i_EjCcKG5g=To>Gc7^iULhMeBmL80?eR2la]gG
]Z`gfeRobVlKl0pKeDVkZQEB`\MdYi=m;BFCX>lo?U?`PbX]6<]2_DnnON4EghT<
X]DY`2:UflYoaCSk;1B0?1:i4U2B4db?ZXKX>ZbCVN<_Z;K7YYXX_@]bHNEU0iUZ
kf_`3i\Q;ka@<M@k;`U0II@k4_>B4`5?ZXKgTeCZoqd9YASQ@mm_WCB79PoWVD57
S0ohhOg^I44mc]4Cg10JjP9l]@6Lb1JQjHR:]?KB=1hbk?U4^38m[X7b;WO3LPB=
iGM8pCcmhUJQdIBQ0U[HJHoW95XAQlXgC`=8lXEXbqF?AFL=j31Z7ShlU=50heb^
3A3ClaLHF8Sk[ZoajA>8i[M?RW7mULgmFKnhOonhMNO[b^H_KlQU5aej:OMnjYSO
4NR1XYVY`JQAe49a[ICZX8@e^eNkdg:TmWiIX@ILN2<[J3H`K:VUgee]A;MnjYX]
WMXEqlffQ\OP@TR@G]U04@H[c0kZ][TfiIQMN2eGo30KHeO`gNEJ9QUE?k4B\^\l
ZV[8WOF78FP6D?_kk_\F<5b8KiDV5Chj7MYXDKL9M00l[CnKk:?@QfogT8[7ITib
Df]ecDF]cF7[d[_do_QD[5b8KIHh6ERpVcVbdOaedmhj5KAXK<Lkm?4fR;0?gJGU
kD[H=ejkaFXmV3KZ<=\WTQ47aU<kDV`WWdo_?\QeL6Df4YSU]gcKP96ef`VF6nQl
iP]65eeE_3i_a4]2nd2mXHjO5b>m>Ce\AdI\?YC@D6dN4lOe]gcK6N:0n4qaQX9i
PQXX]4bgXKAKnWj_ii6AjmfZXQD@ca::U1jB=`3A439l0[4QEC3cC020Eh3oE7[g
fBne16jUFXXZj0QJ]TXbJIf2Wi=5]jBMUCgigfgbOo^>:fabKLo?jJAUj\\<Em^g
M4Go176UK6XZj0Q4hYEG:q;5b]de\B]@?Fcf:2F@`ajTfJ[6C]Uc0SIkcTA7m0eN
]Ii6De?lbff3?:<b2M7PE;R3=j5^eW>lFgL3VWM[k08e=jlIiQOgH9T9LPK700jP
jl?[Cm\0<Y=dmR>n?ZbcCgP3Nj5BkF;l;HLVCmM[k0?T9[MCp1D;9HKf80\mELW<
e_7hbFXC\Q825POYIfn:DlnNeFTS9hIZBMZhJFIADY]PRC2_F\?_19Jm\J=Hdm7@
4dUmNdlFdV;UFJnf7TSD^]n8U4XEDd\21jYTW8jnCVDNG\7mI4?c@9?1O:=4WmKP
:dUmNP@J8_<pO;30C\A:X4V<8XRc4]WAlhe@aHn]HXBnJii?Y;4eFF>meHXF>UMZ
TWjmdfghJ?]L4_I@DQlo20JkE_NbbJ5U<g3FTf9N9G2KO@2bV;>I3POZ_=`;GU:X
GJQR?CT;mG;bF_CoDHI=a0S<ER:ebJ5U5FgolJpDf`D8PS_^WiLjcCZ52Lg<^<lC
_DC1FmZb;jRJ]h:9K_aUX14g0o^F0=H?Yn[AJRhSc<X:6E@?T8BZ7gAciioRFmB\
dKdK5]G;dQ02]n;IUQ5DB=S_3AMQT:AeN[7@MLM]c72:mKS\TMBZ[eWciio`nJ\C
Ep=OK2g79R@9j44b;kZ<ckX>7kMP]I?94LC7aBLlcFYIQ\VJDkje];8E7?^A<BiP
GebQ6M;EYkHL^[:?JInI]ZYeP;5Oj`MN=U>?ihDlF_YS9:TSkjTKJM7Hol2XUg0f
D9iQO0;hLQ@L30:fT=nI]ZSgWnS6q:YLImfQmoRIRa3gFEi7P^a8OjMf=EaOL3fk
ZjY]2@4p=VOD9bkZ899f068PUXSSliWTHMBobQREUla0FBk8H@=9imG?9a0NA5Cl
_ESU2T]F4@ebhYP5c=GE:]E5\C`RfJ1]3mpe[BbkbR76M3Z]8WY^3>?Umn=dURib
DDLon:^oCIH^^M8LMU`?7Cl8Tn\0g>BCabGT>VRcPGn3T:`lWcjCCaU=X9=YXbK=
3;ec=eZlCNHI2g<@5UN`?19Q];RE5^D=3XTI>9Xc;hijTIklW6jCCaUGTgR=`p9S
JIJHi1O5^dMY6BWh9a[\IQcFKbi5@Y9C_9gZPjldX0V:fQ?WaEoiMb04IhfKfc6;
AA5?Z;gm`P3AY>YL\I><mR5MLlFT<IYnf_0Z7K[Q@?J0RCl]]7TC:A<C699Dh=O;
d45X81]mQ\3Am1YL\I8ILlC>qUae6<c]I\W3g;919;NC2OG;oS4iD@EgMZ7?3H3C
5V>glJFcW8\>0HJMF2YXX8_l[l\g<k_4fEmn9ZEnM=_l[40OaYLkofSMfV\V8D3m
PYEKEgoXf0XlRD`\JHCB4akeGd\Z2k4E:^mcgZEdh=_l[jA5RDbq:^^:W6[gXLX?
E]Kh<3l<3JKA8?l9CM?mU4Ue3J>9?9?TdZ[GlCmZjZR25NcM>MGcCV`QJR0fN6@H
XY6X9[1b^OfXdVETI12eVhV9MJgk><4moDUV84F>E<=F41F<4A<B7VPcJI\cb6RD
XYDC9[1bH3TfPbp4U]eW3>;JH@RQ2GRffT_oR\_ZPLok<8i=7G8^hof77h?ae`:N
_4eCZ>PNn:UaaDnXHbF[GOf^n3>MkKTd]4ATh`G1`J5KE6IboOnGh_5`N8271OLA
=QY=Go^W06>C[2NAH>R[fF?`nAYMk=4d]4A847`bPq`^R4?S<=K_kgiREA8[jca1
2An:Ng`Jg]aWWU2J];\;9l@\?Kh0Qg1j`C3<7aPFB]Rna\>b\1Kjc4E0g\YCn_3F
Gg0YMQa@K9?6TX?J5Q`4ASY1hZnFBNA8Y>KD=[G34fonj1>2eOfj>4E01jYCn_Ge
VXDGq8SRGe^K0JLiID5lNNQGSFGNZ@3FbV3J4^=3?NlS^g9SFeB1\M`:K=826Ua=
m6^VJMB\g6i_?f]f8oRh`G7]i@=g6gS18=@1M`4k]QlJ;WnAU6[jHi2Q?FO>ejh3
=m8F86BL36?8P^]laoR10G7]iZSjakXqT`UiD[Lae3acoEHXI9=YV0QfKGVUiM?:
d[96eP;gqH94lg1maY7IBXmT=`hOQ1fCQY0Q^jjQJ_HB>922c=_BlBhPeM18DjDR
H`KCb8l@3j1j0\?GOQ1d2\49a;gdl27m__e1G^UN>_T\dC2eXg>c[HLXS54bb;mF
4Bdc@YKeGf1Si\:B@g1\@\4@a;gdlBh6ACgpJ5>6d_BOaZ8=OF?VA\jf^]IIX_2X
A[fZ6:FXCMYYM9<09XBI@O6S@l2Liaa7NWg@3B8>>3WehN^L_e`2YG6RDMJHFQlG
CH4UKKkO9M^Kcl5UTJ_V?`M1G?X1<_e`;_8TABOl>QBU7N4<_e;GYG6R]?0674q\
3hUe6ak_l8me9g>i1L0:GWIK0USW`lT];O^HbbIBX\6l7M0o9dM5F?\bm^MNKlR]
YBeR52JNPj?0NDFUYoeQ6@T5IqdV^6d6>YiIfXknXDfDDg:XFZ[0@QPPocQ`JNHo
M_<ClGJQLh1Ak3`SXQY3><6nId2>\k`@WE2eASNJ::`8X`WMJRlUmO^19Z[3B1\o
]h0V:=7\o[`@3fZR6LH:TL`oNm=>>A``LEZeiGN_5]`8X`Y;Fjo_pk7hWSFQ7N7G
48><MmK2]Hgk0dB]iFn3^H_1adohWE=1\XiodNZgU]X]_HXJ_dQjinX@8?=``GYd
3]b=`jKHClC;3ehX3LFLUIda;VoP2lXDa\<ITiSa9^_VUBJ<a2^?Y@XYN?>_82YX
B]UE0jKHCl0ST>cp7eiOB4QZf@TTjNU6KPFV32U;=WZ?9B^ld7`6O0D^9MVpMO@e
YB29QOgg1=99OH6h\N\Db3H>`JWh0T=jABlMZb8LiK9JWHGd<]2a=d1XoeN<85Xi
YY=53ENX>2?4[LdSMn@`F3oCC]_C1RM`HB8SZd@HCkDRSREgHGXeJ84TaG\IT53U
YU<hHEbe>>@`[LdS3J^_[lpYm4WcT<bA<[Rn>Q6]JWKo@TgegT=BKZ_6`[D>]`JW
N9FMMe;g@K;k8Q0NNRb:`Lm[C;MN^of14<FaLG`e5OIfo\eHh__H1HoiTTJS]F_8
gC9IMi?=8VjK=5CW9Y7fhJ;FC82Na3>[4mbaLHQe5OI^eNND@pJPL6Y`KcD0dI;M
fe\PiY7i9QK\SZm7O1i1Vo<257HAHMKE`cNd`H>kIUQWDkjfaa_c]E`ij1MMT;^i
8[?JnV@08O`d5AWUnV4U8h82HWM1]\;=IoiiXne?6[MLH<6l5emcYi`UYL[M9J^c
IT?JnV2oSdg`p12`bLGQa=8F=HKa9oD98b?F_CdaX>U]eVmaF<d=SlojC\_\?NjN
?Ojm7d:U3XCF>8N?ggYCTVXU4mBM3[eoJ8E2jGV>[0E<QnNK5fdkAh4m_6^Tm52Z
TjaW_4UQ68>jl]NBgg[AJdXWLmbRc[eoJGFQkMBqoGDZAcRn6S58E0V^Z>n9d<LT
m<M[5RAdSiC8B_DG6EIcUSKi:ESK;02UDh:0d=qD?O7D:`^\RC3S[;jKVi9G4gU0
=?YA3W@6\HHHG2J[;1nNIn5Y?Ien9F;Q1SbdGR@bX<75R?kmSL[4_V5hKd@<IdSN
^l>a]_i7Z@7VGdb494ooo]\F\6iE8Q^Ak4>odihkXVh5nWJZS1W4nYkhKd@U?jFN
Npc<H^j[j4]1Gn;TSHjemE^XY]bA[0c46]neGh014>Y\<IY@bW`iKG]BS6]kQj6S
T:?WY3e\n8Ug5Q4DG44cF8`Y?UVk]bAKQ[Fk[981fmSCK2W8TbTKJhGkL0dLHn5?
RHjW63eL8PYgUS4<KU4cF8FlS5:Dqm]5miZo8FBSYlh^a0=P:Glc30B:i=MAj1B?
k_VZ^@EN9Clnl\Y6BUiniNA4E6>b<5oHSbM;hjl6gj:Z2A@OMI5<@FEOIcl^L7WP
`]VG]8]`nSHQ>bg2o0RMan2\`AB8mOoEdb4W30lVLjKC\A@OM>N2\`6qSA0[=^:E
iYSX571kPB2?T96^j@_P0^_c::KaKEBEBY\@9a<gij@5qjdM8gQa=h18aS5L@JBb
8IfU8WMeRJJHGPY?@KD1Knn:9TU7IN8LLX7O]4>XATd?QWGae:7SYa;AUE4bO\[a
<O\<i_[p?]c>`?J`eP1ImPIjZ;W8ZZ2BEXicbgDkGeG6geA<_M9`<jUll1@QoBhm
oDU;9gkl2BDYCAj57UJN0LAOCI<iol<Z=X192Z^BT6F39V=mMQ9``@dJHa`?`Jal
J:dhi2SV?DVi<AH>7YWbFLBICI54ol<ZV<GNREqB6ci<o_gL>B96J<MYj:fkH\0k
WOeb[\mO@TnGT[nR_nXLI?o\IKDoI4^[hQX^2OTeZgMOSkSD8FYc\?45RXeL`UIG
WW2dG_98G5M0;IcTWnkXj95mV`Z6\QM`jDbMQTVB^?29SXbDbDDY\N=5RKiL`UI=
mRo8mq08Sje<^m>JkAkJBQU@HUHc9AD@4543cJ:U^CAckQ5G[PVX`[JaIKj>kelo
okPe\M5VW\OZ1nR1BW66UK]kFLeIFM^\HXlbXfi`7TPckJS:]FnbaZo78GWJK@3b
ODCF`lTV0gOg`fB1[S66jK]kFLbIUg0:qGIP]D]FSIM^^LIRheSDK3@KWYndUK`h
Bf8YcR>IgO=VJbkZ@P]70R2hDN0mYiQA^aTC7<7BPeNZ1PSn538lT<oeoNmBE498
eI5lb]>\gUPLNjEKal409dPW9?nh2@HV@2T]R<3AF9NjdPS0R38lT30LE1AqkY]8
H@Rd674L201iY7T=e\WkD7c03@iKngFgKPFc^6S0h^QX1>XF2ZFdHHAoGPZU7kU8
do@KUOAEN95H;OWU1]72:7Xan]BEKm7?49@AI7ShP7odKSb:6L<`\B^;BF0okN:V
lo;TU_4MV9Hc;OBo1]72mN>XQ^pL_=0_UQ_=YQI=]2`n_0^C9>SC`]J20K\YcOfP
CIGjA??2F]fKFAGFB@Z[c@P?J7jFnB_1K;A=36a`ehV?jBH<b^_MFAUO\FJH^26S
CI50\BS<8lKWdciei04S1=Vgo;[hn521]bBh3YP`eB_?jBHohm@\HqQ9?S<BCRJR
O>F3fZ7V11;Zi9nKH;Y=a?gbaQ=ZK>V72ORiJmSNV^_A6oN7^Vd4XU2l[cagDl0J
8C73X`@WZJ\WUX_hk4EXLe53FdXZB_DW1IPUUdm2HNGl]c;kAdcVb5^lQJao@>4J
8A73di@WZJZJ[\CDpkc]M@f13GhQ=Lmb20R0BXJ56QVVEAVg_eHL?JA0XbmXf=fZ
WINfPoobYHZ7clE9A6EFQS;4AU:o_V3Y;k@Jm>WZh84eMJ@Sb[n;;CAhf4ACFCbc
nJLLChWR@TUdD6HXSbE=PSRI<0:_GV3\>k@Jm4W@d<Tq>7`L7_87io6EocS=kYV8
GB1dS<YneJGAel=7[f54hMVDA>bHGaC\JU;Q`dD`ZB2XOH6pS\Tja@8LS_66j4FW
@@8XKY1F?5Kd]UAP^Nnk2>P6U8AFOTU5VB=TRjbLZ^8HMN_:[]<4i:XSV>>2kE?A
HJhKQj\gH59fkn6cC6Y=@AM<CO?CHLa`h1?\:U8>64S^_E\\SiL0U:M_VW:WCEb;
HJAKQj\ggdh7nQpFX_^41JKFS`m7]:kF?MnoF_IaA5OfSCV?GMjIkc1;o[cPKNKk
G?DJoQ39E[GdTZMgZQ?DG;mE<Oe]ES7LOZ69c4`P0H3;6qGR=j64WK`4l@<AWneJ
2iTf<gW8NY<]gGU6ofXo2X`9=T=C^V66C:J5QF=<]I`4dCO?=FdG8QTBfmn07f;9
PSmEX6]8M;:AFm\Z@4Egg7W8K`06OFh^fPdfE:b2fAUnkMGQjLRG1ST93nf0a3;7
WemEX6VGc]M`qSn7cnb6EWUa]8^\819ETbW6egi`a4WP=f[gl8I4Sc[@7T]SHB?3
]fga0o9Y_nAgAJ5XKWI^2GEJagAH\997Dk2;L9i5a5J4_bLJLOaQJao@>bNAe?Dd
BUL^QfXE:jjW5S_9KEIcGG=f<5A099>BTk2;L@Fm;:hp_ceh_@eYNfPRmhM`bA<C
5fC?>@NA2S`5^Go@a5cIBa<9RcLm3A;TEX01XlNOL1:5J4ZCOci_Z4kfjM@[dWl@
hJ7cH@2kcANN<EmZS1MUVo<hV5c^7eIcA`C<MB:@fK2F_oLmmcPXZeCA`MoBdJ82
hJ7cHCkl74qPl9Q^dWFSjHh[GRHmRBM0:EYMW>`>L=hc^cQQanT\4cQm8@IO]9[R
ZMdQGRIeH?61B5I\Jl4CU6`YoSAcTFXo]]U6GYanR5`:>L7iaDZ@V33B0D9I0Q=F
WM1Q4aa16GV`BNB\n@56UHIYmckcTFXSjbGX4qGUl]3VDQ8P<jZlB5?@VelQmXhA
2K3\@UfZXS1Dj8GH=`Okj?3]:C`jSIYTd3f`KB^2@Il8dOaMZ[1jRi2aX7doO5X<
WC]NLEE;?T9D:QCC>=AEQPG8Jg5<FS:;IJo_W]I2\OlG7UiME=17oQ2aX7d0O_X8
qck5Lj@\1MWm5d_F\@kPaIVQS623QFcgKU?FU`YhR6j>BI4?Q17BL26Q4>K_Dall
J[^EalFGAn11`2Kc@:DS05XMKb23hQKAhn6ZE4n`;`j>25`Fa5NUb\2ekY91gdTD
AcGS74FHmnCmKLK^[:o?25XMKBfKnaUqj15O6AZn4;]eXBa:;3k?[`c<]<nX3Pbh
XXF1\h:S139>>bU`i4lAU[]oM_d^JT;9K8Z^2\G398MOn7ofTL[\^TT44<1_P\bG
Jn@FFLai=993AWcHi4D=Mc8_Zm7NdFM=j2Wa5\lj9fElo7@PT3cc^TT4J:nHU^p2
fT4;L;Md0AJL]W^n0jkNQf:VRRRRH50ENGgR3KjQC8B=1i8Z70HqYXb;iXQS>mU7
laRPYhZI<OiAbVg[2Ri8a\a=0Ag?eCfgSbf]Jn48k_oA8X7D`^@1I^B5Xg1WgDg7
XeM_SQ;C`0H1Qe]SO]@R8=GgNA0\RYjN:]8RKdMk2o9GM7^aak>T_^UAXmQZ[DDZ
XHB2SQ;C\j=>b0q>VJ2EXTOQ>K4>MMDkEMYD7^=]3nn08o9A8mK2J@H:IldTV;Oo
WCQYKeNj]EEF^l:4\7DVNi1o`@eMnKOnEaZLS;_63Em0>C<>lF^oKAU@[\]M^n2]
n5f>ja^<EVM61AN>gUHCN7Lo6KiSnjRnC2FLS;_?J5RM>qKZ2Pbgn=InM[BYQ_j?
NH0SPDT0>_iWSCHYoo<DJWgd`\UiJGf<H?>6H[F_iZ<0@fW;Anff2P?Lkb2J^c7?
9d;S0O;@[14dq;6d18`qaUPaKZo\^:T:]mi@c7Y<E7WPeX9<=f^giD=RM:DNh?2X
MenUB9OD@nKZd=4SXkDZbi8q^c]3_6c$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO22P(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
UAVE3SQd5DT^<_4i8E]J_>k5Ze7[HT^Dh>iaC4>9lYf?>G:hbdJ^Zjo4GBDFLop`
kC8G\f@e]6Bo3]]cN2:YMT^nVJhH08kAEY]VF@9^Me?6>X`YR6p=jjN]\Q`h0Qci
]ZIT<<qY5ZF91qYnc3f\^bMI0ja?FKVQ^9H`d@4d1[7DBHT^qD:FbFH1G9jNATlk
KiJ>88:QD^I=P7bHg9<qS5WmniiDU;KPdNWJ5S;4md4?A5O=AjQE@YqShWYKcCbD
IP4fH4?^dneUN]I=1pX;bTPK_p8g8SODa\0GTEi1Ag>O1QkM0fATkPAUWmhKPEU^
^O?aAEYIHZDL4eH\MlWBp5X@TDCq3X4[F_:gGg9D>ZTl\`d9l;Y<DdhajJDeH^B0
4?7FYmJ:_1kMMXaFT669D^<C<?aP3iKERF:f:>R>ceGfb:IX_O\l4KKnaB9gM^]3
h7A[XVfjVQClBR=DoPpKm@9C5291PMZnKb8KBa?@D55Q7Y@VSZ[VNX9>gX2mV1Co
CIW=ldY;YYDMfm^<3eGKkAL^_8[m^E?YGB6nYBolLGJT7HWe<d98NZW?eh0oQ6gd
RGH>`GJ2bq9?l3YcaFTecSeA1n2@E03IT:]C_Oo14FOMWo=P[B5GUeS9S=mTIWC2
0PG=RhiLd195ZC5^EkC7g@]TBZi`:eBaQ:1BeQU5FhfMWPN\AkJ;;OjfViVObUZE
q>LMW4;MIl=BYbUMmlSVV[bJ2P>CQ;8=_g=5>9C3E23`B5MlClWI^\6;iW=h<hDM
^>60b<_e6j^0H;DYJR2>452pAZVaZe@ASI1<26b65Egga;SOeb4@dng@JLXodfSn
^881E9T^584IINba=GY2hicZAH3>QMn<^:l7XMlcj?T9[J9KY[=[:=@omL?jQ]gD
\ZlMk84=K3`3?1p1l63M`0BCheQOa\`I^BM]ZkeGfNI2Lg>Lcf1D<1[^jUaO3m>\
S9MAhBocOQG?`VEpl\l0MZ2kc?^dE<[YSYioCbW`f73Q^SPZCJOc\QEFX]F5DBo<
dS3QA?@dF36kkI0^lLg_6UKEU^;\a:0Q15BTlUfZU4?A519ZJJHQF7ABKmTCm@Pc
:5HVo=p>T`Y[JUUnBjoD\^QDjN4^6:J`1g1LmGXB@8U1_WFm1=X9PO;Dak4QB9ET
>ERVg?l>7l3_83h\=MiAf1ATBR_WogJPm9Y?[<jf@nJEMA^G5ok1Cm3NA1ZokqnY
6W`H:NQ5`Y<m>ZfcW^>A300EfeXCc`P<Yd_X@ahTS^0]OnJZg8AccDEoPNXoFDn3
A5eM1\ef6kkamUD?@BS[q=^<oc:]AEHjY6GPH=dhJj870G1diVTV>X93[[UJ@:<P
F3`5:;PUZTR_bc9=Z2T3M51q\Ahan4XgJ9LR^hkN7TFk2^TSFiBZ^?>nNFIo5EiY
_m9jOFZeQjDA1kj89S@6KELQg2R;1k<ToaU2nhB_DKNQ@DelFH;;hV=2R0RAAEHG
M5LdNA>:<OOIlLcgFYp[PnWSO_Z^\:5AcRE[e[;<bo\C]6bQCh;2f_6;>7Ph1cW9
QVP[Z9RA7[;YZ\K8ZZi[Y4ceZC?6a8a1hkg049HD6;R`31<?XdhTfaZB:[Uf_JjB
Pl3m:E:Fbq[okFnBkd:lYD_Y[Mk_6nL`NeE<8ZhaLcdCmogJ?Bf6WX_madQlYKTZ
0PnfHQKb6H68PMFGAH[Z=HJdcj4K8KOm[LFoOCQdD78^kJ3JaTNYEM6`iPDIB[OK
>aJgqilWXDE_645<:A:3k[NLbfHUN5F@360B@LT]j^_pFcaJBEUgg:2<C6aH\TMC
K]@V@[cG37cN[9D@B?fRVk0kF1^U^CdX@g:fMcY\>n7;;PSfh5DcUhd?DVoV86YN
]9Ui`hpEC?;nE6`Jg0k[DJm\Kh4N<5XPZ8:RR6][a75JTEoGo`bBY=1VZ1BWX_Bc
EWjna0:E2HXMYb@limT[<2:eMV>ROCmiRgEe=VB5a<jAh_<:b]@hVM`\ICZ@Bq4?
\34aMLiO2ei@IT`oC@heDDEPia@Hd2QQcbT3UVGC?8l69A6NAaSU<X8Egn52cRV6
MF:Vm@MX>?Nh_\3hXVEn?1hSdQPfT4d^b7m312:`dV1_iaEFPE:g[iMlqIOaY3Tl
V?ZC>X12baJFe_e7V`?]7iRaoY9I;L`Sj870Cc=cAYHEHYAI@`9ge<ecd9OCad^5
M2VMIYHh64c=lQm1V4`SPdaQeRH`KM`ZXADS?X?C_2dSX4EomS4p1Ska4kZ04A5_
Td_FW0\Z85M8kCF7kNN7R8=_g=ElnC=B23`BT;l9iWI^\Qn2W7hXhDM^>60b<_e6
jCFU;DYJR2=:;1q\MfQ``p5RXMhC\H<QghZ59J7nD<QkLb0=OIZ1C`A0>J3gBYj\
h4mIjK0JJLTA0oX1pG=DkZka$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO22S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
;fkcmSQH5DT^<lWX29PD=<hh\gOFc[mUbe3TH\c0jajMNlLO:DN2dN9HkAAbOe3h
nI2JV7=WH8QqJ3mSDM6N:0_\^6M\FNU=a1@_1Sqd?[hbmli76l[\h=W=AB2GeBaF
4TUTV5AQG_OLN8_34PdFiY0GooPl_>cCP_Tb7GGpEmWO:?qkcRCgo2c8ARNScGCe
`bjfkPQe@LA8L^DA8qGP80ge>U>FbM>m_UEZbBX^Ej@=dfSgaDaZqA98`0VB@6ll
J4Mk6e4NRM^:Pfm>j^ZBoS1qF@Y];\LWMRSmSIh_ghE@;>X591p6JAhdj=pQdfYj
mq0aD;G]KEB0P^ccR6@kRWAQERq^IE<5h`4jV2kPMgT9OQll^TJnnMOY[A0O?_KA
nJG4UDLjK5j@WNBA;olGM?HDf[:^Rh>>?YUhWJZ@8SeWU7?Cm^2N^KQLlD^;?_OK
T7WE3j[HJn[SbT5HCpOV[:bfLF1kTQgfFF\7jU@Fh1RLLmA6hZ1YMjX[^Qh4@cMT
7;QROUFj7QKhUKYPE5OiY6f2o\IH<Hm>:H3^GHQmA=W2N>ZZNb_Y`mb9WQ7]lKLF
a0iD2Aonq4NYKi7nA5jS^06k36P?klb@U]_g9UlmnAmhgL[THnoN0i?0K]F^55?I
FjI9YCG`54XgH]WV?>D0Y4AA6Kl=GaA`OgC;nkUW[EmGN61W@Q?5N`Xmc`XJnQnp
5hWOA0j^Y;1j1k2aW?k8;jdCPjC_?6YFLG8@T8`AP1:YWYh@M\WoPQC`8MloCc`3
50J3O?WiT83QRXo5F^UcmQp6i1[IQDX0Z<4kgcjna6C\VVIbh\7j?mb>QLn\1[R=
kPTRo<hJQSKm2lDOlMp21ZCeiV6em?Kgk3PSHefB<K5g<bL>MMgIF5II@HlR^;5D
4bi<N^nb_1M2PYca40c2;M>7L256k:FXJV^EjU6MN[PR<eLFmfQZFdVEfVCUVCXh
f=bQoc6G7p_fGki_?A3E:55jA?[iKGU=>fAGRbEjTj[7>9ZG;Y7gMBB`_6J`>O99
e2<SD`9KF\_9U:Nc6UA?1SeVn`23nf=c86KG6EO?OU07@f8XO6>JCOU37dP1TZEo
qnXGk@5ULX88AZX?BLc13Phd]D:@bK7`Ol;M14Xof;C<>4;DYT0GVaiP^7EA<Qel
anhEVHcE6UHCHZ7EW]0RXWPZLnk0:l6UE?;]UW^HhZPoZ2aM09Oi7B:qPMR__XC[
nn_FD=Ocm3@HYK]U4K?^ZeOb]VbgN6NYnL]Z@`8S4=KTW7;<faQ`HF=PPS6cTZC=
lXIQoEf7FMT55Cp?4;OMC`375Dj64[9_Vm@3E_F?RioX204dbP:e5VakFbIag]__
5QVjbB`XSaBIPVe?>OBkQY:TR`niWdi5o:EaDC\9Y_23i2BJbgH0JK;W42[QaLR3
BhKkTqcOgA7lJH@LQZ8hSAIFk6F^`DQ2co_V7FSi6Tg1^5JoGIZW^Ao>9d5bkO_d
Ea_7]4cj5^P^gW<O@c7IFhZPWTOdV90h4MjTYTHiJ>KWEK?fTKIUX_=OXNk2qFj8
2:F9@C:9:RDghon[YF<nY5cdTamI]lARcR<ZXDCT<nHAf53K0oB\fhlV6a65lHbM
H67TpV3eZWMa21_WO<o`QDDT<mGF\M]dV?Z8jUJP7OR`T=KZ9alIDS21?o9Cdina
]GhN?VOS3f6iThjQ6S=Q4YXFR`>W=ZAe5JdEFiJ`>`ShhVCY;k?J4h=i\jSq:If_
lOJL;:BU9o:KAC;D<XGcRkjV<Zbm9F]ng=_JN1MXHH]j>bJCRD[=b9ha4DFD:TD`
I9E?ha0nW\Ch]f6TompCB4h][PA?ooCGDOUPY2Ac@Vmb=g04B?SI:Ta7L?MC5\:`
oeob3F;D_;NmGHoZP15C0G>mW1ZU4dOaea:5_g9SUY=fWij@N]Sc:n=<4^iWPM_Y
;Wa_Wha>IpGKOgmjbP?;V:Tl51ogb<@d=kBY=887bcIQ7j6@QjERjWnkM<TYNbV0
Domdi\_<Y>P=Ih[[eAGklPG1eAQ0HEFn?a59\EHJaYES>C4@YGI>HI@hfQYSlNdD
59BDpkOFm39U@EfbbkBmnk0J6CQYcR\eK_SURWQELd3S;gfo5;dWe:L4LF0FkoW5
j_CohknobI?JO891=H1=BW]<G1LH9H\\IV_bOBQVa8gAdBlUgHG6FfeCV2mpc:YV
YIPn=JP^FKY^8VVg8=AK46JX\=f0Qm_Xk`FMVXHGgKl]5lTK6Z[85nO4XbHAcAf5
5JF_e9c09DdGigZ7Q=p>1bHQCqFL5c<4f4U@KnQSMP]EP4<ACGD^>6lFG3@`]kXJ
b^<^G9[R2j1bV;pIk<19ES$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AO22T(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
hkRJZSQH5DT^<FDbealh17dIB5A25=p0f3N9ilXRnW:8Lo@d<S9KB<c>b:k2b<Ga
d>WEOK9TFJOm8C:XIpmm]h2mQ2Bc06EJ[\UZ5hp:lfPAPp@G<J]:9?E@QAE55fc8
78^`m0WJX]hen;9Hp^kA55S]h\Lg[dG1EcXN[N[iPQZ_@8bOcV?p6>eb=AT=XEYI
lT[7GB5_4_caZ=4cdkB0UmqnUAjP@n[4=hmHlT?@KbHjOgX;YqE[0;EgMqTLUbY<
pLhKgAQKabam5ffaQjOAD2;=C_VhnA4[`miOKmfNG2J9S:dCAkO_@mIFKTh^BP<B
F`obmd3CMKbI5OXFKY]Mn\]c0ogci1IQ\`[[m:fGGEm<;eWRV:m6O<J95@Pph9SI
WdDa1W?lMGKVaMMQ0gHgJkUPVoYYRf9W;Wao<J5ehZi]Ed]VL_AGR?\_h:Flf=oh
CZg5Z6]F:HE1mkloMADlXTILG9^@1Sm^PWa8N^GHmF@Y75T30TlOU5qRnH]J_9k[
V4=aG1ZaFO:;DEAQhVY_;n6iY:9Cm]emIR0[CP1KXZ0>8HUjC=WLdPW=gO<qH^=0
m>9W9Jdh=d86W:7Q3Wbb;JOiI5c_h>EcJGm4hXIlIEJUoCMfGDX:M\o26Sk8H^@d
X`lC47@T6YmPNQg>7K?E:geB;K85H>EFRe[\E:5bfn^]NgQH99p>QFAm>1Pc:GiA
3ED2faIC0kPOWH400@HfSZRKOTUZgU<79WHaP\V4jRUaLUi@9FJ>PRCSm0Y?5M:W
OLeoUO`>2qiT0K3Ehd;;8Hg5MAJ@ED?IU]J9PTT9]0B2KB1W>9NH8HCG@;cKN9e]
0YW0cDF>aiTGW8lN3WJToHI<ojMe]`<6m\YEi]NgFBE^>[>WdjV?gkdfAf5m^g3[
oaAbpT;2iTWgC0^5FZ`\]NdJ_\C[PCWKRAmJ?2=YWJG8@Mm=h_4NKjnA8SS3X;CN
A3DeHTMVDi[^8EEN^S4Al9[@YnS6lehV:6emCd=;Dc^ieP=[3BYR2eX^T6^q<25e
YBfGjD@H4?[RNnIniQoWK_bnVlL<^E];:?Md9So^QjZ4DhHNXQc\2B6:c[0P`FN9
nhbLm9?D`ofA;C\=DmacPaT\TXg\c_eUF?LQmc6ZK3\RYKgZgM:E>CqoMA4VmNT?
YS=e_[Cb7ZCEMliRi^aLBjn\C?NF6Bjf@=S0l1Q5fAHY8C7ZVeWRD9D4Nd_T2lQN
Eh0>Y=d]\5_accQgEp;nO@WoM4DQO5BXTEkTRX=g=QhmhCJ4g@n<aZkPc?mb[[c7
3TCCiRLaK8[3a6Mj7T_UT[G2[7D;k[X:MR]hNCB?R^0KP>TUY7lISB`PSXjK2ENQ
TD4dAk[L<^^Wp5GIXH6`1e<0dEcZfeFF2makn]b[OHgmWNRRSRCNEiEaE;8>J91a
9O<X3<W3:\3UKm9lClTMfZZ0:P_XX\O<odH4d]N7@hED4k1o?9CBM981cPL;;HZ?
B:1[<l=q2gabLla>6PX1hIn\O\G4Am=\omkZWAAhWCKnUUaRoa@g9mRNoUZXQ8=P
p<L:YYS0O9kPXICm[FXZ8R=J[GhWF0n`ZXLb^e93VX?0\e6GmC]VloE<>WZU<GM_
IT9JUM5\N]bf[@c[cUKi8:B?0U_RDaa1]QQPUc9HfalLPod5e3IP_2?mRI1pd;kN
lb1;8\g^8NQM5]?D^^:1CDBLe0Y]?@eZgX<6[j>DHM1[[il=?boWe2Ee=>n70:Ia
DD31Q=Zn5<nl]76f=j`]lVphHM3\:U]2d7nCB\6lk<ii8\W:>SGK:>fQj_m8SNjF
J<T\aH[E=AFKWFBXML07TinCb\]Nm9k<`I56`2@4j24:EKe0@j`hH@VY<Q\bSn?<
[GF=FbjIJl7C^\7I1pJe[949A@?0bI@@`lF<iK>Wa^KlNb_RICe3bB3kgB8n\a5]
l1n8E[BhTlP8`7n8HEUm?U:HK3?DP[7ZiKVL^\=Ah?NZ0KLd[5l:<omkk;H>lclD
4k^>V@j>9afNq?YZLMWGNdamc;UmWWPDC5A\a`B\4\6=fXEHOKf6;6F4ZKiXc85l
E:kBT;<T:A?FH\hcJP\H^Y:DaL2fYj9>lh@Qol;C@_9Lm\Ten4f\4gTV[FZ`f>k4
J\9;@\NpL?PY^^_8@ZI6\84leQ0a5=Z`h5WJU\VFnNk41GTQihNoBG5_AjD0<`NX
^gkF_0eJ@6>2@KggOk^;lm6L1fN=XXNe^]q4\dY7>p5n8R`Z:3O]1BNN:?l0pIAN
WXZf$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI112H(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
MSa3`SQd5DT^<oQRjn7G8AKAKaml?;lJQQJNIdP56NoqlT@M^IC_U;hN1421^cPf
>_BmBf=gjTE`BA9We@7S;`JZe87T_[8IVBp90k^U1PGkmoOkK?_0L8hUGLiMKqn4
85cnqfR@e]kWlHX_?AUh4=i;3PZ@Wha\VQK[4E1pKhQKZ4JVBTd=54XmiY0@?IYO
Q@Mc0[3;maaUf6Aqlic[gU^[2dP[MLH_3i>f0X@MXQgBmX:TUD4O9LP>KY>`^NA6
JODQI1oXMFIR>gO^Q98pa^Hd^6YpcPBMI^qJc`Md[XH7A>0m>Q>_O>2foa3@DmlZ
2^h7QAHi\<Kehk5OBODPLLWJBc6IA>;2`H7J?122]oELAK0F73RUbR:N`aFl[k7c
<_`<Q<HfFQBQomoGTC6kdTKZ:qnPO9F9B>jgPRV4ocl0cKXD?YJFK2_hnM>@h7n5
1`D8^TZTd12BCo7JW0p7gUK_8FYdmdEMM[j1CU`ZU1k@^673Vc<<iWIK^J=>G;_G
a;YliF3;n\SfP8H7T\]7=o\KJh>Wm:HYhY_>:UfD]VNBF4[529hQiEbi1^YaAkVZ
ZCkcjL4b_qcNG_2IRK<O]niiO9RS0ZbXl;]<]Q1OHAe7KBU54LfL7j83JS^R;WIg
=d<ChmSRh:c?:QokA:2O;_A@W`?aE16\46Q7j`3\LQZ7H_QaOcB4Q@<k3aRY]4^A
qgh62iK:MZjBdm30kM4NhNFT`en1=k0ICPFniTja87`B5nGhEdFK?NlZ4[5=hJZX
BgFQ[UkTjRj3[?FY@HOOV?5p4e`kETckgb[58;A2?6H3\JSSR36o?aeNQPId6m3d
fUPLakl`5VRZk>f?f[o]Ok5l4ACDmRY[EbkEEU^;`a5`^Rl^?Pj39;X]HPI_V]@i
5AAREm];Zd06n>q3d;:82ZeebT3C>Cd4bd[@S\pJecn<dPlF\ajAHBP4S]]:4dD2
h^eVS`WEC2jc6P>8?0HO6BlYS9EcXCmf1K@T=HAJ_573C7eT\037?PZ@BMGhKng<
Fe;1R1NUCd`1LHGJMjcVS\0BnTHdDp>GkAaj;E4IOa8@cUb9XHZM_6SO^Ek?;2F[
]Zn^Wl`XmBoLdfc1=E]?QJY[Uh<L[@>HP;Ag\4VI91i`OCm9XP;YkZ4?S9A@mTB[
QVM`UbUh3V`2HcRFoDA;qM;J[kWa\oi]7cWHR_2F=a7TSVPZlbhc@enYP]c@c]4>
N`PVmA8Nn5DM;W=GUjk=:MSK9ie8Pgi7Y;05Jf4^aO4pK=9hk2pNM`b8T]@bi`GP
KX2MG2[7Z`4P2iBjcQ?e\Rf19a7eh19dWRFV@k6F<YhhLdBBJ`aNSMVB9a=Fi;G`
50Ael1p:kFeM\f4f1ML=KRd]i8LPOm^\RG@CUMenA6II^cZiol9F9X<AR4\LQO6c
cXR8]`S:0<;PC\nl1Cog4K@RJjphQWFgXD$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI112HP(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
L:N=MSQ:5DT^<e=:9Le[;OoD6?>9b=m7MT9[4>S6P>8OWaXYWe<f41cHpKg>j7je
`EhdQAAd2FoE:OTH@aCq6D0=Cj>c1Ni^_jlaLVB`7OR\R]T?Zn5R9L=[_gMmIX??
[IhA?8189LV2_[?oEWR=B>QJYLAp5g:CaDq;odOXa=DFT04amW=K\nhoSbDdhf<g
FLBV?pa?Q7kg@M9C?d@Z^YOg8E2eY[54R[nW9[KbKU<CAq:P_<OY1q_bhbL?q?1J
7?G\i_7U=HCRV7eT<18mC51Y?13o\hI7_Id:Z0FnY?Ml?lIFQ<iN@ck_6Dh<b?;0
k8RA?077P`L5VIJleO]kcg`\KZo9aHIO_81EcY4Dgo^8gLiMAc6p\jlDa7eVk=Z8
ZFnaDMJK<?lAfmmO@F_bBbMh?0M?@>Q4oOFO9OFhWk4L3^P_bDda\oaY=F?l^=j?
_>lJB8JHL@>1jM6iom?X3bWhNJKcW9??];NgU_NfZdqX\QIKno`=;BGDbak>CYH_
YjlRO5c;`]3PS;N3IVW0`]g^fIU7inmpQL[]N<4GgJN^GEX>g2]OJR^gbL_?6_2M
9SL_mdTV0BY`WHdk4ITS=K_E4>RCF0HhQ4;e\oYO>J3MSPe6\?^3b5[n<P:i08J3
fSL_N67deK?b^I`VI;[oWKpF@Y]R2Z0lO:JSXY>HjTChaBDCE0=O@ahC14MK:Wk\
h:H75L49fRJ06i;MY`<=B_YF<2ca_0FMO>_SI@_>HAR8Rq5`fMJXcCCU?RDLL5>J
iHTND;YSjjKUEej@l[njHUh\YNRaO9jIf3O5akKEPI\Tc65oMB>[NGKUGN@;j7nj
jFcO54Chl7gj8;S@S0\dQi_N21;NZVQ89X]kp>j84=QFNgHX8J?C2BQTn[n]mPA1
=gBn=jRNl;91<CSaS^<n9I6c3JM^8>CdX3cKe>;hAcPlKmHH8UZ^5Sml0afR<faX
O@mmi5RNlF1LmIT]9DiWBIEjOTlq_L[f^=cnl_OTVJgVK9J_dZ[GmBmNSZ<6STW^
F0bCoQQORPLoPiA:25:SLIdX<3cJ_g2h`k1Lc_HijMDn[3JL<<3Zejj76FZj;TcZ
oJdm:<6Hdc?ec6KDI1p?jcn`e]80[YcoKI:[QJ_hSZldlgm;fJ^;a8e9LgXQ^0G\
^48RPFSW=Cd0BVoam7S?Q_SW4<U;[Z<FD@Ld>4VC1qMN1Q\nE[neEJ;AS80nQMUA
6pJc0iL7p]Kcb@I69529?Wj9ilDMOPA;?WIaLcCLTmARAFSA1;d@Y;2ERm0bK;Ui
>oRXODb]X]QfhkOV>@2f7Sa7j<7\pnbc;XAPjR_7]P<SG0>aXAc52MgEBoK[k8^4
HodCP8OO:iF=?i48EQ_hKXM9BA4<fn<:^FG3XT_T9bI8mEG9pE\E\03Q$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI112HS(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
^oA77SQH5DT^<6[HQ=JDSC5;LJ\1b6i]VT2\P[9g?CoRJGOj6Tb63Peb2j\D0<En
^a@I_ApE\`328bBO<ZHfF`aY_[b8`94jL\G@@2_XN_ASmF;ZHHC[<9Y]RJP\Sd`q
I00ihX_UKm6XInfZjK?>e>;NOPL>0VF=@d3I6i5RUni13dO:YeGbq5KL^gTpbKgF
n<J7oH\mlY>?iY@kZhm2BR5Yd2Dk6<pCM15QEKo_XV[4b6IWVY4Sj_\oPbD8bimf
XcVc]Rp6\n;MHCpmk;DZAA^D0B0L0H=80?c=n1>_JZVB9a1?X1O?5NKc<=Ub`?8K
>pcdCDXlpaW];^67c]?H[UWlKTdSGX:?OSlJSfhmgLg>IT5KoFG`HcgYE5E@Ml83
CmJTcC:S8ab<n<3JmL?k[ADEhSdj@W[_Q@B^9UAW5fg>BL;Mfc9N1DEnKm4=<[Bp
l1F^2@F2?hXdm5aPCM3R7=f<n^N@9:WZSVeZPS;7EFfM@RC2o2Dn9cWQEVd0Z663
lWOhVloYbhYcdmnU3\3iDnoD<S@1DjaX^VL5=LgUh:7WR8Ge?M@MJcpW6Q5F>=k[
50;GX37j=SER6<7a24W3R<2EZKS>?I7JE5e4S43bTPA40SZO2b:IDXEWQEFCKE;o
5O6<@gSO7E1]Y4bmWX:jabF:ZANib0@T2A47B:dFENYW<pdb]:NAi>iQA9Shi537
::ae`:X24E8ZleYoE^i`dUQ@5_5GIOo7TOEIHjSCbC`4RQdHocKn2L@QV@2g\8HN
?[\6q:f7[;0[Y1NYjDjMM^5RaPo91MMUDkX7TMU:h6YALd07G4hC<QS0=H:X[0`E
889YX:Mi>eV?^3NdcVS7_@_lAQ=AKcRnTOA[7^U0E9CCe6FiFV[EE2]<f]6pcQSH
>`KfTWFPiloe1;91YfLA_6LHFb^;kemgQToXDW8c;@^[@JDl4YU]Gjj9m3J1cl_D
FT7Y5Wo<>mZn9Z6LXkdagX<72O99CeMMbjO;SULKdK8`YH1jbdqB2_:0W]XMUaX`
BPI=Ec?e>DEaN5<PAMABO=HMe=ja>8;NgJ843kLBBkm1?ScXYOSBSWN54^Q_UUO6
V1A0[c8^CDe0AYf`>mM6O7o[jGBXIemB`6CR9h2mQq9JB]H3Jn1BeH4P_`WG?O6O
>MZ>2f>Eajk0<eDVGHP`hSMc>qKMAJjhbQZi6PB?8JfY5]3=m3JL@nPRNM]idR4]
AmBa[UKQARP6oaA51di56FX8nkKYL0n1QgFiJCJEe[Rn=oUmpElZUBSpg\aW1[Mc
;]UP[D?JANEo3a37OJ2BiT09K0=d?3HK;;j92GcVflnd\RkEfO2dkfELge8d27HN
[gl]L4f5OnMpdI0J\]<IR4ffN5N6=6ieASX^76LGlm<aB4bYSiBfV3nDK5]V_A@G
SX^^TMEVdAN4d_lQJ9@D\4I_K8P\Zn4qSM8[Q0V$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI112HT(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
Pd;EPSQ:5DT^<JCHL^OdYfegp4RG@SDT>hS_Y4L2U:lXLO;>ZF5?lJhN86G?LN2g
=ZjTa]X45AEWQqIe?@9f[C6`Kb@VIENFJoIoLA?CYJV]dU^KHR2RgI=30qA1SRg2
peEKHP0BPCVQdF[>5G>_FgScI:kSATERF4OpJONoMXi47o1YG4[5=<n=Bc<hBT:D
2Eh4F;mc\VTpZo269^cqaj;G@eh\5\G7JBA5EJ3Z?@W=b:_fhZ2T`_P3V:5p:8gR
m8qVDmMj8bOAknAKhjE;k7;Ch[O??3^A=;2>Z4Se4=o5YK>3;[cGPRI\2d=[KWR1
^R<V<=WME15Kka1i78^6LnKlA7Y7UT5X6i:VZ@ejl;ZWnKl]Kg9H`Ai99p`5jgJW
Yie<YdT]TmU7:W^h>[fIKV[gHW^h=Q4LJ86D^iABA>h1[BnGJEgnLf;hPN`Ci4MZ
BQP<VcXD4l48:3j]C8WbGlglYQmhU`]BYOZcH<^`31ObJQ7DpXlbdfY_ogPV\M8L
PACaJ1b?EWGPH3BG:83cdfZg68m8ncXDZ`7had^VF\Yb4D4?aXP6UnXXCEPl@>h0
@<L^5WH0SkKnG_80aV3bdUSTX^k5k83FPii9iKTqiDI;C7UfAc9h_DU]HW`JZ[`i
O>BESPKWY15ePcQCYjd:Md3Dm@HNH2ofgkf[X:C<iTPNB0Q?ncSN:F5FJF`mdmpj
=5n7:iBAe:;9Y5>cAcmC:DCY2=je9W2H]inqFT^3X2<O^mBn8<c`lYB2EIo^1EkZ
UidjhEW4ioALc1\^\;k_W?XQd6PWEJ[Yg9XJFSE6bH_i4mCf8;YC=\KXFO91\SZZ
TUb]^EmDb^N>SQhCEfXd<O2@;?qco2GiRHcZLDm7\Y8ZL1Fi0?AWnmjoX<d;4eH`
cUDT2^mKa[NXWSZSS@h6SLlh=m[c>m<OA>Q^L;m1NJfOd45a`TBiJiH:`LeL4POI
9aI:T>SeGd]X`T`2BpQ?k1TfMH;iTB8_@f7IfccchPIhHhVRb72h1[Fg;1Q`kVl_
km:H5l7200R6B<3;lnQM:UggY7Gi>GQ<@73aflAJ0hH6EcNBmechCSDNfQUkJQ7Q
DiMmLiE8pPcO?K5cb>2FVW;EHaOaX0PEhH\Zd1MR?OT33c^b0RFgFL_2NDECd1^B
@0ARaMFiUP:oh^^=LA2GQ38K5OUg\g9q7eD=VKq2hcV\A?UZn^4i]dJWCl34Q1JR
R?jOFSjM:ChQ[KhncK0>OkJAMPl;Ycb9BoWSf@F2mi0\4QVon:=UV8OB:=qJjeeo
hf3cSA\[@LO5?^;Q_QCadYE7dlejUR<2J:TANN[5o;hd=V^K[BA>c70YbL]J>EQ_
oU^mS;=^WEBHB=q[?@jDLT$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI12H(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
Di6EeSQd5DT^<Z;`GOJRn7`ganP<8VjL3FC]SPq53KSghhoK:<G\<oW;UOQ]_G[3
e\hb5eBMRk3o8@;MEXZ^HAU1MKNDOnB]WTG1bg3SO=qH9<hCaC=fPOCTfJR1f@`Z
?j_[M]acVYT_2KGVGgSb[HFZg^LEVfZKAJ\9M\\q\GFTU7pFE8M\UCmSWY?Mn8iX
D?<ePeh_29?A4U7aBqiiBH@=JD:3;NA[NdM<:L6]8ULKnY]cP\pR_=2XTSpkR=BQ
mqlC8;DP8:l?Qa57pYK45ScAa7S`nJ8a8\N<gC0=k`fKbFE0NH>:9f[C\BFJ:Gd4
ZQEGlc>NK[Ag9ReWEYMe2dk0GLSE`h5dAejc8;Q;;JfUe[nCA`>T8jLD7g^;DlCo
goBAM5Kq7dgXOSTm@9e^GUI[R6CTCY2fC4`:o=@0j43=AkL61LmTKeN>AEoCg=1i
n?5JOe=>7l?jElPRD9k_S7TBa\YF^X24396CTT?cY47C<0\kE`^MafhTFSYG@`q0
1`cbXoWMlV7R30?^^e89XKYICWV^df13CL:2iX6fMDi?c46YmhDP<aahnL>OVe70
9V_hEB:ol1lSj62n^e4HW`FKCH4TYMfoCF?AVb`nI^CV7616jSU=Tq__V<IeEacM
bTR]Gd<WTh3JA\bY=0RL1eDB5QF4KT`8lT9b^J;OQbl9IX?d>62oFL_Ae9\Q=SeM
3khe73]O7omIpEIOKgIpXJ:66ZI4;n:\l;:mG3?@M<[n\EO<kD2;dlo]Y;`D=E2M
0DaI=0<aRcQ_5Y[?0OC@XK1KILAFk3@lEDbI7?8q>2KA3:]Y0>meUZZB;:XZO6OW
n0l:dV5J\_o;K3DfXFnCQ5@bDmd3mQh:dVBn]m<9>Z\TocC9h>c1fTbVSY\qH2]4
Tbn$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI12HP(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
QE`j@SQH5DT^<G<YAa595>=5G7FJH43?hDUEP?<ZEmBY>YV;`4ipP]Fj0h4VAj<=
;0N<Tc@YA]SkLX4UZT?Ld9UIMBgYZ:C:Y<D?h7KoDaQmYj?YqKbi?534HQ\TnABQ
b`KbKp;NRC?6pYWhMQeD]Ej6T96?ROOYEO]l@n::j=a2a:^q::g9g?8@6=3PjPSl
2cbB`P93nn5464I?pDEEUoU4p96CP:7qoc;hb?]:@TB?LL_Z8kQjN]D]nP@WNA3G
3N:\Fd6IO8fMC62MF>3`_FGZN[Uj0Uikob=V6F4dYT60:Ma74K2X:][;bF[93@J1
ANhNVEZA^XZn7QEmm5DlGmpjJ3^aP09^SQKlUc3kH?NUVnhaRb6df_]N6Cai9W:D
aGMCZim_kC@QWX9ee4o1N:Oj<\7`l3RQSSQZZiSb<G56Ij`?R;_1bA9X65hiPd\k
>6;?Q\I0g;LCCqnV_SQJYgQM[>>oPFhH>QT9<G:\AMGP@\?b@3gIYoF]KkCbQ@`D
1B@G5I7CDNd7[3njRX=;@0UMN1a\h\R=>0]>iA:CT7XHn`HbO@;hOBhHcBoXg5R<
gLU6qn]k1k0FAk=WjU[obZ44HJl1H:X7bmg8]dZRaKUN>dHo64Qi8AUQ>CeG4@oe
:QP:9nD0?6DLW>=d4GfjDj=;Ao>pPBI3dW?cg8eDH=D_YX;\1O?ZKJGOa=^ZQZ7e
U^J1M`bE>XqSD6:eGq3I^U@81Z1`C<T\hNjVV8B1j;8HNWF0LJc@a>D@5=HgCk<`
gOlE]l`UOJ]2bRcOFS3aQh2A94I`4h8U0TJ=Zqj>4[>5JceHOc=E92kFN\T[S7N@
W7S6H_:d?gAj8cX3IU1\AQD^W[EJ;03F`b?OOhj<IMLe:1GHIc4hXo8U]pGcoF^`
R$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI12HS(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
@JO_YSQ:5DT^<He11\\WWo<de4Ved2?iJLZNUI3TW0d2_oWJMd6<35ngRbMB7]EG
qO8iMhG8Roe>;C^M`lgC@Y3N7DIF;i1R3?SYnZH5=7DFl@8;p\48^N>gFM]LVB_0
NRN9bmhU==CCAYWVVN[eJNUlN\YSh1ZV8Ca\m[03bqTkoBamqQaC9J?B5UPSCj_?
MjE2Ie8:W3]S97N>]2@q1]IZMNASe`>cYA6F6nTZdCNCEPCbMW9NpoVF<c^Sqh@d
VX1KYL2_DJgd56MkMmXOSQYD^]o45J_:^JEY3QO1P4=AXF]KCE4Yp^^nX`dqk0\X
M0;1]EPcT:=4:_oN]GYNX]AbZBo;[e=][C;NMa`I4jLQMHg\W3m6n3RLl91hkT=l
ED0NNEbQ@`f?i8hJXA?FcbT6KTdN\e`>2NVAd`HH0?Bn93UW0Pp8`K?=Z?_Uc@Jj
B5[Q1aamTOE<Di@f]@nSg\Re2gDE:4TZHePWH0`9Hb6MW:k?1X28ZP9Cj\QJcoAF
1RP`IhdVZW\dg7PZAG=Bg<SVJ8TUSR;MRl>NB<d05qEOEF@gZH3XGbe6WiKF09>B
mZUGig0>PaMofTl_i2hYR2lfLi00ORifUNOEe6bAMqaS>KAF2IZ6OLSTC6VD9E9?
efJZYD[mo\@Zh\14nZPNm>_biA5mON9BKi<LR?]ND>aRND12_OP6J[_mAAgb9VYe
Li`JdSmR\jTZEF3GmlNZMEIo1NLdZWl3qYWi`LOiaDmDHX^OJlkAKaL20[I5BLmJ
YL6jE50;_X;Ha2DM`RHJ9EEd:1CDME?nbYUZM?`:G=m[nMAeYIPahk0pO^kT26qO
aml08763I;6;jdEmc=Cln0I8AId82d3ASoCVEmIoQoSodlS;B0AVAgW]6:enihMO
5?CQEP;Sk@OB3dK2XNp?E9`X\@@ogHJC]il91K48fiOdF`9IJh4<KHgC]bb0@K40
ho\?AG2JHFeVG;69G:0?053:Zj?YgP5aM17=d^q3>oUL9e$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI12HT(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
@0AXKSQH5DT^<gh:5cReH3i<;FR9;AAGO9`nTlRPG6_S=@Wmmg^ZZPJ[Te@K`86k
iJiadMF;B;\kBiXp^<39FPb?O4D[0\b7JDSCG52U7_;?NiLIWDPA]:FKP8`iD>\p
al;0VHW4=2VmQkEaVgmj210k=_e4oc>P42XO0VIoHS5obfT0QomlOn]nOXVS<5:N
mmqjgab4?pF\EV7iA45D`0efm\=VJKNjfX3Qefnm<nknqd>`Ud<TIJ:RiMTb[EXQ
Ni>_f7bPL7CdSqc\eK>;9qjOiL\6p5WcBiKJlW<1WQ\ah@EQ8W=4k684ZDP^NPUE
B[<Nf;Q^L_mJhQcX<=a6gb^M8g4jG5EE6Vg1hJ<3g=S6iKnhfMU;`N\<4^gF3LU7
S^8b<j9^F5T_`iP:>CCqBN?@Cbl@Xd@QK`4\P`oHP[efa0O;dNnC4NBQN?<TDo9D
7API4fg1HI36l4N8Z5WlBNQ7ILJHDd5Z>F9G;^:EBJ;5d0:8K:F>`Ng4iS1@fAm5
CM<V6BoW_6pHiXglM_\5>feN71FIU6`EcE;l9??mcHeFHBk4SX2:4dD2h^eYSc3P
K4o82o`mUFVH@8cPn0`J>j9l<9<A56AT7:kdYSDU:@a3HYPZ1:5BjPNZC4=:RkO=
EpAToXbg0hfGWCb4>?H2O8aSAdk_T52Ll=U43_2J8C_XVLAR<g7`IqA5\fh?Edj0
1;5XAN?BRV[VLKMY:3H1ERAZ2D?1HW7WV8]5R@]k1e=k]9K61nGb0\AQefn4;350
76VS91Pk`@;CpW:L8>VqYkXc7<Y0LVomO6BY>9=Z?\\aBLbm;``7gaj:hmJmoo==
8OHeARjME4Sm[_nH\4@8YE73nF50AVdj0`I;AJ2p\V?3bdBC2m1B`?Hna;kY<3^Z
3admP:L1lIKl8HNjHgA;dP]\HCmRJWK;m`Rh0Vdd\JWd_TlF]mWO8eWV2<gpkgi9
@NX$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI13H(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
N[9aoSQV5DT^<iAlDW\[]FC3>UlQRdF0qTPGI:4dNeT>[^43k3C9<Vj]_Vm5hFJL
a>?q;S]W[5\?^0@Q3<FV4il_m[T[FG4B`XR8?0p0Q`7KQq@b1RJGT2i0UWb<ce:f
3Lg@@kCOEfV0L9oLV;3RKFq9SoYbN@7mcIiX8m3KDaKNB9XGi>LdAF=p\L7n=Dep
LmISfGqWHiG:8C@kX6WeQg;8f@B;`CBOYRC=EC2R[I6bMeSj1d1^R>PiXDiT@D6Z
CcAX;f]=J9kqi6kSnW4YhAnNAY`K58PFK8@]aV4l21^@ZeFIYmhc2QI7:J3jPFi5
<0gRAWkmn?Q_i1BTgKoYOA:U0Hk9:anfAoQhFV05W[nj:ek8@aImP`gK499Qb\BN
^L6fea3a`OcCok??Z[pFR7IC4Q2dKUKf=:KO<73E;M0KTi3RCoDMV4Z=e;^2;afZ
GVfoo[l4ebai1NLk^0aF5PlIKBULKSM\b<dB0cMXnYFckRGOT1;?V@dAgmgh_RYh
T?64]oI>DYgcOcFS<OlPT@PinpfiJ@e>hH^O\^^gKCAAnRmCEdE4B3LCgeT\3O[>
L=KZmM8PhCX]Td7E`GL@cOiN2WfmC9JilBDOkh\mm=XFnOS?2ZlFc@`4TFg\0kdh
PjRKkd_ng1f[BEm\eSn2b;ce_VZ^2<j1pHXB:WHCH<>Ygmm^f4`[Y29QbL5oaqE]
C`@P2T?<fTU@4G7X9a^A9lBBff04eI:]fA>IIYl0\H2Ue2BA:_KiK9Fa1c;[;XEd
KB4@Lej<TjG129EoTWUBB1^BUfKlNP]]oGa^a_@4C8S^2V06LYM]2DP3WhcCKODK
YTckq?J4Gj_DWSc?Z8^<P43nEmOmn[7HSk`J0:R:4F<5k6AJYmaC]E5?XGcbP]\l
W^\Oo?PbS?m3TAc<UVn5LNknTD3I1d70[kZeO4RSG_TEY>BiS46I8fNf9A_4GGVc
aFXHMAlK@j1qo5K8\VUL73hi?WgifUK^@WZZH@^_>i0GZo3Dg6Xd9aDFA8DRFTMa
:?o`8WEFJnfHo4iZIMGT<3@j8G=M_DKV]3A>d[\JQRS]^o1E7c_NTSi=c?V8ngS0
1PAe]1iN?BZ\8lA31VpL>Bm;;go\8;@?QULkI6So7B1aF3BGW4KfPYin8`>8:T[i
llGLTmJd6EFX>>L@kZAL2<`hjlNl8\iQ8VZ`[n=?n>f`H:CDLlXgPG`gYB>hVEVF
U`WmjF;ieF>Y>Ylda2<Wi<I6nqS]g@=^]V<72a;Mf2TinRCg=MVblEnfO7`a]9?V
TNo[n2?OTIONm55c3E@O=FY>DDS_Je1<]e^7[`9G17CTo9IIp`1XnZBpeUm\EDF4
oc9Rhb0l1HhV]KEKk1K?><B02V\MQm9fj04=aW9KkkY3Madg\M=2Fi83eP:3GUJ0
a?N42ZY]?Z6p`:4N4cWK`^a\4P:?3ic^n^LocUF3eM:\9H7;?<eH5E<XbW@=2P:F
3=aD0jUca8pDHQJ^6=ZIR43lTM`gHB9N4Rd32;D2VilEglZ4NdIkE9NK41g0MFoW
H[DfV[`D;C=DHYGL7?HNR?9^Y7co<bq>lUDMZK29Peb]5TmOVa7U6=7D?MN4WWU2
J2BA;;A@\?K8\Q=dj`C32X4PlB3Rna\>b\1Kjc4EPg2YCn_DY=qVH>Djh9$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI13HP(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
P]>m5SQH5DT^<Ebb2VJHA_fg>U?CA\[=?cm1mC\FTSTlJIqn4Z>RF[n]6APoU:P=
\S6Y9SSOl^fMbJ^SL@:]H1@=^3q[XVh[bom6QXH52MIpolUNK=qU9U@7<J>1jXY[
SbnCKP]R;a>2RK[__JaNMX5\1^_qa8N5B>\Wg\G2R`Fa3]3SK0T:`CB9iPfMq>_:
]i8<pB_Mnb?pS74d`Ikn;`OCPa=cPCaE`4O4CdjOYV6kULHONSC2OHL2<kebBhe7
^XL5ca;HQ6F^SGE2R>b@F`R4]kM5?Eke3=?ndd>HGHFB7L;T:o@kdEXk^6OXJ]CJ
lI5=17R4^?aKJcoo?dp`DN<;lTce2Hn2BkWjUlB5Hi7T:hWFFRiE5=Y`jd@HBOS3
lMAmTcA_d4Jf<;Ic3AT`aCk4=H?N2b8@g>ooF[PBXM4hM?`B9m?U5;6d9J8K13;H
fa@lRFk_jE1T<GBOM\NUDi[?AqOamXW7mXZiGT6cc2X@RgehHO\GfPmZ]_><YOYc
D6WRTn2laDdE?lo`e\XcVV6]CBOO:EPI04VieU^H3O:dRl5_J11Q01m2[AM<UNU]
aFJ;d4c7E1oFPeUB5Sacmdn7Mb?2JRYSp]4\iehn6g>X;8S`l>JmkcOA6^kDVVKB
4PmZBVU5T0VMQO6pj^k[UKSPd@AliP7OGcl\C@J\hVeR7XSBWQX6h32?WdPRKcFI
\n?^lY:?;;Dh4Edoj:cmA;JLF@cWN9K_lmO@`I0l]VeW[BOM9Qn@hhBhCAASXXlL
P?jg9L@:PKTdb[dagSD9PRpA5lo7jmQMDg9WG[bE^eET5OFmaV;nn^RHAGcDA_Aa
k<TZfhGbn15mnIR\\PVW9>ZANgDjDdjoDjHf2ldZ;eiVj16]aQA99NO[AKl:MY:5
GWDNQXeToLLfg5A2P\Fg7hMTX?E9dq]gOc@YPLaQX<dbmKU2O7C`?\Ba;[n<GKYX
IQW?`R:WIQE8HbRHgLFaPAZ1C;=\R\]aPY3PKd:QlBC<TjWAOaW?0EMfm\^UA75X
IS49Mk>Rj[M5YUP1NUHSTGk[7N`BEJHenA=Dq<mRf\naDeBQPebEiM4L?m91N`df
\F>Q@fn=On?k9ABge]0>fp^Od7\O`TX=Nce98nK0=M^bRnFlWTiPDOR6Zg40\XWV
9P^LDmTKRNcfI47W;`IZKe^@@Mmc7WF=Vh^OSE5]bH_0Pk6@HSMBEfn6W?8I4<G[
TOU3?NJGZ@7`jQ]WJ=Rg8mjhjlbep117bDRiWWN2T>OVFk;:;:G>7en97YKG4e=8
?_0`iJBRgJhhe?oZJ77JBY>`YgEKW1jhHf6Rf9N\Bh9>C`La6NXpnLGYBhq<Z@?<
E>hj[0H34c[V^>aXfeFK\>3o6=VAeanFF^99_AkRJlBMi_lb=hMa=eNN1L3<mAL`
ScIcVAJT_RNZeXp7NniCJ]bj?oX>6oj34;4<4UXB>3G6m2KiHf<e9E<B79PYjV95
4]@_RGea96M2A3N7__N2c3]k?D^U2\nH_TpfmOgG`P6>PilM2MQ_LIRD7O8ZVf:8
dkbIQ_T_jKOU^3Ug0XN6TMH=S7;NM>8:4]TfGhhDJS5IPaX]`KhD`Epe8i^V6Ena
ZRXc2Hqa36^D2V$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI13HS(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
6?F5<SQV5DT^<6GaVML8Aia>[ki]Eon=j[<oUkj<M:oYm?i1nBfiCZJ9;amp;SKO
:`C?6V>0>nH`<hR\e<0[dS0aHIp9[0dZohb6GQ;[>A267K9K76n=n6Ub:0XM0NX>
=?SP1RAT1q>HgUh=pVLFBM>SUkag3:<FFKY=GHM6;RQlQZl<=?RC;d:7Lq\1=Nd9
hPBco?_UiC^F=`^jOkkShaX?eCpWX_7eN>qkXBF<^pC_`^d<1^[f;KdWOb\gT]HM
;?XDk7[Zegf=J@BTRI\J6JnQ_dOcFYEe0KOCB6IbmaC7kM_K58RfCia<hDm6QDcE
_@QK5ocLQa]=AFQI:^915B<6bO4R=4GVh5T<O2h]jNMHN3ZWq8n4`an[G4OCCPB`
OeMU[lkE`2?NJlR<bOnSdb@?<O8J;BO;RE\c=^m9c_bkgHKO^8C4OeSnTcO8<en=
>@@55aZj2nmg;hFR=lnfB7cK]LRaO0WKT59ZhY9ABH:>AUiSO\l4Sm6qBgaO0<Di
>hoXgTXd1[i4UjHhk:]a<bEjUWG[5<I_`dIV`AcTClRf9E0jZ>3RAlhhBG=XhkVD
^hC:9VBKVji`^HV=;]]6LHC]4W80hh:Pc_6h??f3VN69>1_;i]_N=LUIb_Yn]9pc
jQNihDX]odgAd_@0_9:FhCB5Ql;YE9h`acR@`Z7a?E=FmiVBeOijU4J:C6AWjT>c
Ca__1N`ToU\Y<dX9Pbe@OWQlm;OQ8hgcaNVG]iTl8ab`F]lXYOlNgUa9Ul65H2fJ
dMhRMpTEdmTm7Q3_3jZFJSj==KgR<[nF3pnUiUiI?X[4>Tfn1HFTPXc]204a3g??
jR^SEd^9AFSJo7;iOnOGdAHWaZI?kNk@9=nOJib0idF4U;P2nQPIPRTmW77OQd3U
UO=SR]FHAoN\RD83^I=>5@JWUmN\9g=3L`oSPoa`pFm^_PTZj=^E@Omi\>00]i5C
mmncJKAALTFaY>h4bc@k;NI9bj?:_T3;gWmRjI;ZXFgCbAeVH2^`o5=[_g50gI[B
g4RS3;GPk]F130ibgP_824f6im]V4gW7G4VB<j;H@;`5bi^q[AjFO<?1`cEU2=X:
=06ABETo?144RB]mS<G1KVJ]dWWodQ_;HEll81XJnYOXJLS6[aYbdW_]NcFi:55e
d]jCB6mI\6?4g72Na<m=Tf:c0W@:Q]?h0D?R56==j^Z>1^Xa8j=QkdqU3ZhA:3F3
_RMgdPCZg:`^hg@`DUdJaW\6_JD=XiD?6FlCRKA?I\laP4W[e9QH8\TUkeGO;N66
_dWMX^U>de@<6q@R3;mep[ga6\4GcIIKJVomlk51MVPZbH:W_=_gdFfDdCm97F]=
NdKG?4\cbK24]L5`<CQ<6[7k0392CD5bB9f:DeXQqOSIdYDhn7[=PA8CFW1GAaLH
CPQ;6d@XA3V3Zh`egT1^MAH?LFbM:lBQ9BX>pgbZl[mk7eh]Z:Mgc\:fe;]Nd^aN
oYj0NW5`a[`^Hh<<1MFP4YHKfZPji@mC::j4mg64njbi\iEfffHhibmUpRBK7e1O
1jd3aj;TJngdbUR`d\M>@:GoB;iJ@bY@@ahgOdmbTDeo8bacdD6U8YXdCR29:B^7
SGdNaRdUCoM2pemfmZAJ$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI13HT(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
FkUlmSQd5DT^<o1l;SSJ]o>Zna8Hfc2OLd3Vb];=18X^F[99jR8HimbX_jk>SmBl
I9hXm<dkpl0GL7mMZBT^B1BZ2MoQYP9BfS9]NOb;\AF;bbT]gCoq7e4ADVoii34d
HES^NR05>DngKYbnHclW9@mm8@CSA>Z_4Ln6l;0\OkL=`A?QY_CoVd\Z^1qii^Jg
HqPAZim[;Ggg?SdN<Y::Jn0VfMMf4kcfK2;1T9lTSGq^_oMAFYdhZGgDH7AA:NAi
D;``KO@;F_eqnKP^;\KpbV5?XlpHf6=AmAV7eFQ[Sc][N^9m0W2[M9<iYG>Jaga_
H]@\h1Snfe4SDhQA<O[0]1m`2R0HBGQJKaJ8e^R[6i=VH5Z;SU<ln8]E0MFga80X
8m:^F3m29XOKElWahWmZPL=h?OdB[FkFlpPZGd4HXCHed;Y\[lki<P?NjanJ61VR
3:05VZ3M7g4>96Bm`EmeN;^GDb[7T<2FNBP=bT0lC46eoNWc14?<K`dDHl?nl2@^
hji5AMmNP21QUN^5hG_>a=6ETSo7E`Amm@_B>bIYqZRFN^SlCH<;OL?I<NH:PQM4
bIAd`b5R96n2dA96D<RjfWg>[97dKUl:oZSkXR69gZ>oBb]^6c<525aBLm`:ZK\R
N1cIfe=jF8nc:8753f>okdFa:ERF?e2H^9S=KAFYmGG[BO1q]UhomI>@`:mVnT:X
gO[R\C;>??Mi>Z`51mlT[BEDYXonFRX0Zl65e6lM=N8BHnV7]j]lW0h>::E5eJY?
NAaNM;GSXROF?d?ETm7F2DCXV[dJBH3G5Fl`>J_AbRXF^klfD>DV[cpfhQTLVPZZ
li``8;BOU70<g\KokfYVSgQH]JPkkQ?d^X@]3892^eQcBq:2m@c>R7EC?^OiQ6JL
nZM:ZbJ?_\5P^BS5c?g<50Dc0_GU]>iP[?mnaN1HTo6iX_:g^B^PZR\CilObGDEX
nNRVVH8TM9B6i2F5daOhHAhJ[<7OI][omc3=YKGO_BK:a1oGMnS=q=\NMo17lE@@
V?<@W@KHD?dI23VCX879RORL=][jbRLIbVk`f6Bi^ZPLlHKPeV0gW=MWjL5cf2@X
i=B1?75HjYk;O\_5NDG?GZRaW@2Yk]]Ca6@J1EL11=OnVg\?bP7_FQhJo^[pJEX^
^QCW51LlDlJ0VOUOO7mbF;nOE5oEHN91=AXbN0fIO<0@h_;I8B]`FOj3KW0fJhO6
G0T:11gGa9Yg13Jj0O]FMg;]60@hmN[]B2_7DReFU6k]OX5Z[7_I2OPYBIPGC99b
W4qj15O6AZn459e4UKCI3SGm<4?@SX?35?Ka9jBTV:]4]KWQH[D?6iDVCh8b?U5]
Fd=j_YH5\Qj95];nH5U0aQ2]4p_S<6QCq>01l^6VD>h;oQF2_]53O5Olk0RG^DPB
P1gdY1<Q>BU]@Ii?Ao[AlhIMGdG0QS4NM>Q><3NGnSQ5B[ih<KD8qN<AgBAN7]SD
\nAgao0]5Q=5n73k07SKjjb?L>6E\P:HVY@:L_N@PJnWb:ZN:Ril7NfUBa]7F4S;
JnWh]UP1pBaB1iX5fENNgYdL[Fi_E@CGQQ_R1Sm8=IRpGmJ_X6`O^S1Sm0=2IFBD
5:alWaZKZRBm:oVJ:?TIT@`NAm>KiN`BRnBeC1ELk?l6GS<Q4V:k4Sn0_Ab8AW0p
\2MRn6T$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI222H(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
UAnA2SQd5DT^<hWY:W3bglT:S9Np@9m_i3@dfT><\0?o0WJC`V>[mcP=W?AMPcZm
<Spm2@37WbB3PNf:?]VGjg[1L`nXHG1^M8?E_5aG8do=X9TcRM`21fpoWODS4p_L
^i=hcEF7g?Z_IoNDS\?[OI^GS[Yh<fi1p:B:Yk\Gc9W<EPj@>ne9LmU@aNaZnf5:
m54pRHnMZ4i]46RSOi;JW=>B=2F?;M7_[g23ADfZIWa3pA0fZg6lQYLh>9_glJUY
LfIf\T3;ClM7I`npK12G[gBBZW_F:[Cd6K]go66b4U_THjUma:`k`mYq4a2];i[p
LM1OE8pG:T[oo]TFmL;]o2RVRC>m5`IeKI;jAl2n[3b3Aj6Gf@Ch9gP`Ch>@bX1H
@?L@n4YGDJk_Ee2jma;nMn<KRC7UUaii:@<S2Wfo[22OdF2lKFNchcj<Q:^NahD]
OGHonZ9GZ>kCE5OjmQjnMn<]_idS9p57[MYIl^A5?7>6m;B]KT]3j5aB`ZQ2Cm39
MY8JlQ@WQSkCGRi7l[SBW[dK^Ee0OE5Xc[7SB]K573KKQE`cbEi6dPmdnUSMbel9
0h6dAI=gi4o11NGM5kIPH^6LA730:F5;hG3SE]K5Z3KKQE4\dYMcpcY0D0mnDdnB
kLQI[b>8Y>E^bnD:3g=[oQ5UmRomHTfbdddo0X33Ef\n[H?Li?TSNcEoH^De`JnZ
A]>YhUD8jBAdZc;m51?;`g5i<I:XKihjUh1:FFlcN_Hh8L=FQ[TO2cQ<H]DRVJnh
_]>Yh[=CHGJpco\1NGKPM4E;?Jj4<[UM@L@2BIPW0^Z=KI5jPd:UboMbgfo^=0e`
]R>YGhR67XQZcgJCT<n>I4^HnkS]J[Z1;F\;Oe_L]ZcQ?IKEjF8aC5X5?Hi]ko@?
jk]ZF>1GKXlBcSj@i<l8I44HnkS]LL9]HSp=aW;keD9obcLQI8AnYUoJSmNCIJP4
[neQcGa=ZOa9Fhg0Lbo:^5`jmAkE5mF0Ok;O9EZEmpAA`4^NSQE\D0TK[U2Z:NCH
nYEc[J4gkkW0=gJ4Agi0Z\NiFHkAQ8H^IU4\Y0f=:7AShJ<Dh[?\cSjF2Gd1CFR^
4eAi>BCB]c<0=5mC^o8j[mAa\<N`WOKmGdH`6=J=h^AEm=0Di`?\CSjF2Gee`[om
qR;kgCGh[B^PL9lA68l6\`j9M6e_K_B5k\1A8[`U0NU?Y[=JlfnQKC22Wk9IY_P0
;RTH4U8U4EPC[hae>gC@h8<\V3X[8=;<Xe1A2hKES:bYj>EcMBOadf`:j=3i8WPN
@R3@?o8[bEPG[hae>K?fcB[peEKHU^1?9@lLJAIeFhfkD6ooT7ma<_AYej>WXU:h
@;n36\j\K3k6aMF64hiEeGO3eS_H_l3fC@Xl7Q>54c>00@EL\GXcIEL]ej[P`VfN
\T9f_T:F]e4>J0>YJRDW]Gh4e0=M[l=NC@]H7Q>5<LL8j:q1gXNl:AX?]o\`c4am
Ze;KPb2AadX50OTm0a7Gk<WV8lD_ln9i=G=i2ogC460N35618d]Wnk<0]m\=6190
Z2IP;_TED>3PSMab06?_OnJj\?BGRQ@A^NX4;Cnj\UL93^b1fG]SnQN0]<4=619l
Djbk2q7?G[14nVIlE6Za62T[l:1L_=PDXl08<i3FYUfeWjS6pem07Be<:C;S3I]A
KC70WRVT:`eG]^gHh_=GbY9H;A74S6i_FNEeio2k?n2iGFfgde]lS:3C=`;Y3M8B
=_a0FNhHDSR95dM[U`=<?ne5h`?:AhA:eKb_\:hU3Kh8TTfYmebanb33<`;UFM8B
=UodA@gpGKOgmd]m?9Eog1NI76i9DD<;aY@`8XNalaK^GN9WNoR3N4_b8AM_H\N=
56>8GF?OG7LTdf4o[9SBg@8_PHI4E8q8ZDh>j56;N9[8G315bSWOPn4^eGP\P_lS
@UmjW;K83AjAo[`bg=L2klBQVZVCiT?8X`F=^=WkN<0`omR^GkL:K99N8F3F0fGH
@Um@?1nZ5I3MUT\L0KSNn=[AL9gei78878o_^J8k1E?`omR[50AZmqKN]ie18<o3
c^Zhm9]SIDfDdO`hEW;4[eG5_fE8Z9i@\E?8gkj_hA1[dLIWcJhFJ]Kf;icaNR?3
Ggacec3hMQo@0g\K?C\Q8iY5oefBj:^2DkLJc0^0\cTna^clAOoF]JK78NYacV?m
8<acecf:MBY9pHhVNDO8aPB:PSNfc`WUdD?;<eIeC@Mg2DDL3@5GTA`b2`0^=1Vm
EM1bK<GBl]8UZHgNZeLmoYBg9<KT5`\E26`6Z>R<Z:EQUCDL2A1]e>ae>:`03j<4
mf??@o2l_`8FJH=i7>L4\YEX0<KT5C7bod6p2:C0?[eY^llhoBFj;G4Oaj3QibUH
5H2nAS9YCCDD`SnhZU:lE=S5fR83=BjlD2iA2[2?QPnO_lP:Q[fT`]AC7YaHBbNd
:PY8ISTigP^FLeh0>6EaSGIJZFZ=CU;f\2]j2V2Q0P\d_1EPQ[fT4B>1gYqaLOMU
l4PIHndmAU?R?;5R39l6Gaec_9?\6>N;>A5iE<7I@aPLD\lNQ5:oYF?d6nna8UH@
cXY\H>eP[Xb5<Bj9FZMcGM2lJEB@6gY37>@G_90VQDM0UeCd3YOQZbkG6<Ga[lDE
c8A\^JcP[XbJ[XEUbqP?MEnL8][8^M3i_1Zo2F\fB4?ZnJpH4_eMS2[on\6e@O>b
NJ^R1Y\K4iboiPjFXlTLU?[ZO>8QRn4BNY6Bo^=P@ZFice9H_D2^<?QDn<6J8SF]
U:AEE7j>4fCAFONLXOP9M65SREJ<RjCQd0M\:3WZ1G[`c[9HiJo=<3LD1DgJ8SFj
nWce`p6QcHWdAF2e8AO:Sh`MTMRKh=2fNB2n\iL:1:HgO9maK@1XDj==_QJeSH?0
N3bHTf6]M9_BE1Se8ocDK3_aIJol@Xof>`kBZgo:f4VjTECUHo7EPS2ZbC]?MoUZ
EQ3HoW69S?RB^OSgagcDK35Wf_c9q7JD;F3jdNS<DY8KB]EE<g>H<Sg96jTMZMY6
NNZVZ323C=fKbeKlQh2Il^=P]TaBnlN5Ag08VA`4Mf259f9b98FSHLXbSB^H2dfk
3hPL=<aZXF>eDjD8D:hedl9Tfh[0RWN[0g<Ue^`\SfS<Qf9b9XIJ;gCq`md;5Ul3
AZP;Z:<A4eFBj;6AEM``;Da@lC0U0g5UMc3_<nEVLVF@CF1FHTG[^h0j`b<206G1
MZTh\CE;>bC?U@OF7EJQU2QGACZ^V7D4?d1DCBJCh[BTCS3:ji4GSh;=`gmZl6LG
MBKK\CE;_WZVc4pH:fZ1`\K_T9H^4\39:7\mhDZ[SaBhY`X2T2bgV@@1:oYB0HFA
m<XhZQXle@@mL`mHYRi2_OoBTN;GSiVVV5F>4q39\]j30\=;Yc`k917RgSgiQE8J
J>\I:i3E1h^Y5Z700<RR43ed\cPnSfbk^\H46K3EZ3Q_HLEl:JC6?FZ5H0<J@@KJ
Uh[ll>iETK1>Y^]XVO0?BCi8k@gbdfBBGaS4aN3]_EY_?0El>hC6?F96VQG?q\=^
LEoZbd;g0BBiYl;O>nmRBk;@M\fhM:Rm[Ii<5[dl1^gQYRF3]a=^D8iJ7p>`J^M`
N=0M@Mb6@O62m_]D7WjYJlYjgX`nTCe?QCJO:I9dlf`Q3iY;ZDb=klicZ4BWHC5>
3WT\BY0kb3^Gh3J^D@39eBQWiK85Nd_@g^`HEaZK\5VCCI6X6onId@KfZBcWe?5g
b1\\Yj0kB3^Gh3_aXeg8p6D>9\`ClMf9U>@emYaTX2PlG3K9R<eL][CiB8eMHA;G
EB58SYOIGD@?HHNXo4T>F?XDYb@?f=WCajcm?@m40J^K?FKQ1T4mVM8;O;BMImiA
6cY@Mb8[9>e^A]1Go2VKAaX4HbDGT2WRijcJ6@m40fQ;`Odq13N9GbijhCmfV:bQ
nbe0C@b5K:QD\GIl5FeW@[\67C1hXkgNZRg1gJQcJHO<XHOm1>F;8PDjO;8U1[IX
8BnPk9bm^>\3Hh2H4Fa@n6PZPX<eJd`MXd_\JBl@b2iU[H2P1b?9bPa9O;I21[IX
ASR]L9pJ8eU7QBhl:F`@[id6>9am_]>ZhglGG2S<_o4RZ>ZFj906>MCpTW:1`;?b
1^KiJX?C<?LUjS1\j:R:4oLNfOhGXU?[^VbF?XSMRlWW:_cGQ9k`alTb[9MPhW6l
6jjN=TB8ML<NXUH7Uk6C2Gcd>24DLYM0?@nZf;b6l^4WlYl2<nQc89TQR91Dh0`e
7jM1=TkGML<NmmY:\kp`m73JhI4GCiOYcSHjkjmIGU=j6=8URZVF:>_AQTU\FDYN
hKD_;6M]`OnCN=YDgWE`d[<`C6TI[R9DP`B^^lkBTPOh97K1_6<P:>_G5TNgZfch
\G6QP9YQR4aWgZD8giQ`H6UfC`;I[UjDP`BZ7^<F9p82dI@?^Dndl[FZTk`HY;OO
CYM?PCU?cCl3ZdlEQh78HVF=U6`MCDmn_l<g5gkj?o8`D^@nW:^LI0N65FWAmh4T
oSf`W1KH0::36fKfKDP_?JSbQ[:OicFn1D[kTZAj^d8Q:_Fn;I^LWMN65F5YTAL?
pR>76Qdi\WNBh?V:Z1GdZh;Of3NgM\H9]N]k\L_lnLTcd;^Dm:30V01X>^1oWpUP
]\IMUjWO@hU;>iOQCN<OGK:6W@R\Zab:bHElonih]QFB\gBdkH@=9R>KCMJGUPU?
YeWl8lK6J:9L[noJhkF]4>TQ_j8^H2S:b^]RjXPlkblR^?4G9:ENe^X89VoGJOUj
^YSl<AK6E29L[n[A[Ri^pGX1C94=MaU:FoKi_VLcc`8aKO@amZBR@E<\f>Eg0C^W
I6[3B7SDe2I;71UC?jUj:GTFC360`0J@Y3J>69RXIJaC>AQXE5o4Zg<LR>ohM6Yc
_RC8Ufkkk_2g3n3eZaUC8GUjGO6VU0JkL3J>6BXlTl`pBnV?1R1cIVlM[7AM_5c5
ILRP[_N7jSIU>;;9X`ZMWmK@cCE`F1A2]A;n69:`]5=LB<P_EbiDj2@bcoAahP]g
^Vp;]nfE`?@UkI:2hCT;TmNcK<5k6E^[CKF6eEJ^lmK=<]I4Zd`KMgm6\l\`Oo\S
0cS;=^WmDD6;kWMeg2aVo88Vgn@Wd7jJ6f7hedf`fEebTW6<n0FGAEdkGPkT?Amn
0Qf;jbE^DDM;\3_eg2aP@l[96q`ih]hMG1oeEbUU5X]=An9c:gdhBnN[Oh`cbI]3
gY\2j^ND_F>>5=W@@NA\VUo1:U3HdCXRV0L@MW\=[Q2C4[J16MmN:2<C;B@iFb1W
gYHX?;3eZ6fQQ6d=JSdT92N?m?3HRFXKPU;@^d\IKG2C4[LbX3F2pN5D\FmdE[2]
YancI1noTGm<o[Cb1_cW7aJQRWH:k20oS`Ynjm<`o9[bjg[`HiKY=BLC<bdNlojK
1gM7j<NXe1F9Ff[X<F0;ok1adi2:cdSVkU;RkYVYg@knK\1_UKMOoNLB^bJTN:ja
^g3_S<NXehldS:=q<KFHnaE^hMRXn52eP_SOWT7ch@0YoJGJ:YWRYg=YgXY]ee8b
Q=;M1L;HCfYBg8lGPBhOg7q=@2]YNF\iNBT^O`9o;]KkPe?lDU`cS]I9?6BOS26a
NPQ18]<:^WkNb<@>^R?@@D66Z^G4L1>\AWoPeK[9]m5F0PLWKERhA58=mUP=9QSl
f4\OAm>\JVlcKCBZ<63SOOT\ZL74BM9^A`@P<ig9]m5\\BSEnqcPlc927_1ENGL7
i0eLYP6GP2boeS@I`2iAU6?HM9\MOL4`mb`]\[YfV_kB;Em0=[CUoJbENdmh3m\T
2a8XK:NM2fm7ZXgX^\M64G:j^GW;AN=EKIARF`JWZAVGX0H\DKbUGhb[CJOh`f\<
<F8XK:Jb]ke>qHBFUZ>\<UPa`olnkHm]NjGmdL]K7]Z`143[D8SO0bL4\i4ReV?\
c5o9C@\8[P=MkTb99DA3`lZR<C^Tbli8dQno?GZT7[lGM4nlZWEbRA9F3bH7]UFe
o3<h0=OohPoUiKb?KDQ=i4ZbjC_e8li8dk8O:gbqL\@o>3C8Qj[<i3A`TLVKBm>@
]S4S;`LJDD8;f825VEH6Ye?JYI<4D=GkT9;PH?iNLIDoGiYA2;kcS<VUe7K>`_lJ
CZ?lLo3ODDnUkPem0f8=b699WFeM6RG_JDNP<?g_LJ5I<i1b2<H>S<VUCo0M1`p?
6o7]D6^8LhNo[\]?f45;BQlI:cmA=25MHMW0@=3^5oW7biDV?D`L^fb\?hba7@`?
Wi^oHZmK5Y`37?4]IdbBYGaZ3l6NIck\H4E9HDiD[eKdIccXAABBVhe`g05B7oD?
U<7?H[:KSPC37?4;8AP2Pq]]>9Ed93dBN@Y1CFbPggOhNPlN:0?]E]oZ0XT^8@NF
jbDjWA>9>HCWOR<B0CmRZA8DQW??>Pj3e_cl<US6PjJT2f7B2U<L]>FCen8]8Dfa
giNTQhamcVHS;`o=E9Ae=a<Dm>?^_753C2c@1MS6Pj?lATQAp^\68f]4U7m?[]Vm
4\W^NVSGA>[T=[@4GcCN`2i@:g@`lPTW?1WkKFiKRof5=C<^@EliXJ>qjm`5fW4X
_JRLJa6D@DNSXC6e9lB4Z3Fm27^^ER4;`YU0=5Fkb5@6CMCKW5fYo7E1a`ajIo<k
K5[@AUS8VdgnK6TMgbpj:HDKbOB^VG@G5lkh7]_dIYPWCB;=J]\Q4dMRoEMYOG`g
T\4?CN;<PF@HjXlDQ7:jG7MRQ4gPJEP;>2al@kmG\GCiCFAhfZK:4950I4n9gKhN
VmN1T0l]f`097n_;QhKjJcjFQ40PJ:D;>2a2H=JdWq\bB[_MU4C7I^\NEUOkTXMZ
f\40B7SBCQ@[acloe^:i:OO=^oeE7m47l?4mLlUf^0\L5OH2e:h]N\6TKUBoYIkR
[O7@SbV6V=e[Pm7=aVPQPhi_LH1PN<NMom[@n>=fmJ\U1Lc2ggh]=\6TKUb6Wc6>
plSRJco_4C=37F>7AQ?IWn1B_j6MjS_`6D<1?[oJen6jHMGXLL<P\_YkWLUb\@B\
2lIIF]`CI7=MGm<B6a@WB4=D59>OP0h?\b<jl`8BkoneE?T?i_F8^E7XFQ:Hh<Bh
Kl_3W\`3f7=GBm<B62QMSG9p<^I@Ne>3ndS2H1iOB3DDBFd?i;k\U1X2N5U6NL`1
CJ^BiIZc5@90?moo;]b9916G<>UjC0[d5<Moc<DjEo>MHEQh9l?_2b?cl59Z;j1k
L_3HlAm8PibGWj2Wd0:5[1TG<l1]E0RC5<JEc<Dj=Uh6@iqKWCQ^;_ESFZ5Pl@oM
CfG4>O@\XMeN2P>ZNg]8=:Hi7RSBF=Kdi?D35OO]`07NPPUcgGU[@n5V@9hPY\8d
Z@>WZ_obECE6giiDk:E<8:L7[OQ>M^bU9L?MY@_YmXZ\<:NYgma[O2<B@chPYk^d
Z@>FTg5\PplajfLDSTQ2Nb=QWUS2BQ3^Fh6hUk7`<T3iUJ8niEl5fTXAAKGT9FL]
\^1?EcNE87J4OR>B:OEOS=c65T@nOng1KkJNkXSV54nOgBj8i[5e_9GHn74WIMIQ
n_QP`2Y@]Mo4=[>dRfWOI3c6QD@nOnm5OL87qVY[7lmIZ0Xkc2PJ6S;>3Ac_p:bf
aT07Ab\MB;H<Pc55EUHje`l<C5lZ26JbhQnJJMfi030PNV^0jAlfH^g@NMMYJ=<H
?WnB8]P@LBO6SYWOl>L;]1@<_BGDHF]VhTF6QP4NMlmBNSN<e4<<SL50:b\3QH<L
:WddHgPI0BO^DYWOlEh6odnp?VgZO\:3=;I>Oah74Gk]kNFSLNNK2^>Z:SEXREDM
429\c\d6YIUY@L@2YkPR4k8=FTTWSRbAR5_=:oQOBA48W^X[^5cb8hc8J82;XoFj
^Fe1SVFOPL@U\9?Am[5NDPa0FTioSH<@E5@h:oUOBA48LkfAdlq0abCh9mZP8[kB
^04O^dFLN[m:EF4N8=OQmLiPM:C7\U=nZ0<E5U7o7J\0>6fNYNDWiKI6HaYAXl<i
fj79mWWZV0^[lHZ:0dKBB[UR2m1^l9hkm8dfaOA5fI^MC`Q`kFmfi\[6d^c8XdWi
f<U9mWWniHXJ6q<aA0N[Bk^bDJ7IdlBMW5XIYpd`\ehgmMGacg60^l_KjmEVWWc1
><=U4e]bJW:D:FB537:TM]=2IfUUCCkfi`=h5]H<P6D\NPhRDXBgEP3iX?:jBmRD
qI=NKVBTQG4=eaLY[I]Xb70@blC9R>5cX8\17fe<P=LPXE[^a2?PbGcJ^8JgZEA7
^;k^n17aHJ[WB9GKMZBN9a4N<m]Pa08T5:jR2ncaTW]_`2U=[<V6FQh7Vhm40Y4=
Y@k]l1W1Fo[@S93h]ZBN9j`IA9Bq0E>83jV_X8R[mL0IX39\Ek13QAg14@SLTXNk
2FaJ:J_MGOKDGY8P`]\>oGn8hnR8ZPSkgh`@5TkJd]9QWCPT5=7@SJL?TeDebBn;
<aa1>dFQ^fO]eBn?M<XK3U8nHd8e3P9Ig9b\\T;\d]PlWCPTKOiJi9pc?m3cTXoj
Wo[Z;6AK@F=lTULc7EZkSBZRAOXi^ng[FQ9oUV8bjg=CglC^42iBmY0ca6WXLYA4
0]ZNJ^1]WT\j=1mW=V7VkkQbA`\Z[`_lLZFZOccTB_mdailBH:ZnmmNc5NUALd>4
IlNNJ^1G6\QH<qbToL4C]_f[C<DfZP<=T<1fG8>1LKM2[GkWlLoXO[f\>VoKYgi5
1m<G4kRL;momeFY<;Do]H`;k8i5l3RE]`W?;WY<X_<Wd9gD7kMkH3Vk[6H`g;mG1
U\REG;C2K`Rf;1b<6<o0hlQk]55an:E]`WWYjQoRpjdM8g5><h6ia4FMo28_jXHH
W9g]0^DcBb@gZflA:bNSOan8LkRAFk>3FObP^0R?SWGae:7SYa;AUE4=_\[a<J<U
i?__`nA^A?nJjADA:XC=5L6P599\mUFn;ZTnlE<6]JG3T:i4[B;52EUbN\[a<0\E
51lp7HliSblYZ_kdOeEQc_4>h2IlI<P^4Xi]Ao`H6CWaa@=e@kKFiCUPg>H<8C9N
j@9chfW=h0ZLGa``F42Xj8T<Bheel9Tfh[1DWN[0g<3;^`\SfS57fJK=RFS>LXbS
B^H2dfk3hPL=<aZXF>eDj8T<C2\J??qOUUY7489Abd[9gId<Q2n^6d58O9MMX4hE
aE1B_1?a3<6:=N@G0?lodTTD_[FA5C<hnf;BJ2KcK0nXGF^>EIan;GLT0BaZ@NTZ
CdfWZMGO]PTV=0B_SV:TfoTkF<6HBoDonEcBUaDdKfnXe0V>EIaROQ^9Cp1RBoMm
i1b]NZf1O\RXXOoLAK2>Wl;l\iqkO^SiBR:FOE9j0Y2617OQ[6aOXc1Ij90T;SW^
A@Xei6dD5WM2E4k;_\31WF`k;Q<n5?i@hUW`LVM:VL<7VTEmT2QDOmNibT7IK7DX
ROAb?;<Q5X\A=S7T<m64bPAHT:NV5>M@kRUHLjJ:b\I7VTEFF4]W<qNM`b8J25bo
`aPKSaDGkd7Z`4H`iBncQKe\lf19RddHOoWn`kR8jn;30g=T_f\<H6C2kdd_gn:5
b@AYWkLX`E?85K82>9ZC_7W\0AN[518d>UM23;:SmFl=Y?jlkPO0hlJ2b^dkCIa5
GkAVSGLX`E3afPM`p?NgN6Pj4M5UH9^\H3GNAGPQJ3:YJ[0\Om<FLjE`Nc8mFS_n
V_<foT9N:G36XMF1e]7E`Fa>WB=G1neT7EHMXJV\e<^qhK\MZ^p2e^7G2T$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI222HP(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
L0WK7SQd5DT^<WjMd?e2PMiJ6N\^1fbomOHnfP8cqH5WV]c8@YM?FN7<dQQRpOVa
P25d2ba5Xme`Y:ARZ`3ZD9ZOhbA<7?Ug^ebqcAST3?qF:[mKBf^VIeU9\H7h?;Qe
bRC>W^YFTonLGq=cJMlh3BjjVJfZm^\GAPoFH:NT0Y53mg3Sp^EUTZa3`LF9WGZo
9gJFg@O=Gj0kUDm6XJWqjRFFbU18S=ZZhfYDLfIUhn9M5KeJJFVc4HFkAGUqATRY
=WB;4]]TD]e<QZcUJ1P^:QCLRI7D>7Lf[44@CCnbmSC`N6f6NK\Bq]4l>iknq<jJ
BAopYVVdBUGXnTcFP^^:[Y3g1DLlRL5MmjDUQn`DaacJOG2CGe[3XmHfW=Y6In;I
>:1UY1l`f7R1;THe1\LA633aSLY<2h8l3m5aQnDVolCk7H:U;?Ac0ilAGYcOT<cf
b::XYJ8C>7KE;TJ>1\LA]\Hdd`q=;MF72ER8ZkOnRhf3=J]FT9BV[`U]K685CTfT
]>n<`KnjD_mLeBVL:nO_\j0J[UA=Dlg;^@W[ZZB`J_`Tfc9IJ[?3VOJUDYL=C;2M
0RH?[d>c`2VJK\i3<o8AZCdn[>1=Cd65^WY[Z6B`J_`YjLD:VpWJSd4WSD6=526j
e[hk__nObnbYaMn_nJ?On\lG6C`iJmVO7BcN0U<BROa:I_=m3YW]cBa`Cc?=N>Yl
HZM<_:_DL>XAMB=5c<2O9VLP5C9PkJM8iAQM2>gTWnc``:]mGfW0Gdk`7P?=HZYl
HZX\l26Sp5Y<>nMVVRDM5;Wp]Ai`a?NJfbb@FMafP[H?2_i`;H2KHLZMa1>;MgeZ
aTTo84:VWL9OP\T<B=CXf0M5]@mZLJKZCbYi5V1Yn004c9^\:3WiZ5;8l1eFY3FW
^jQXkUoc87ai0FblDhIkc0i8]8RC<J8=Cb`>5V1Y_V:Na7pjO[?mCPH_SOYD;BDG
\C`XW`CgeRjVIP97gk[VY7BLdH4IOlZVK@iWZ3[TBMgQd][jiG[f\l=?SVD;TE=`
S@Wj=Hm7lSdl]b;igA`m3bB;K3n<N[6=Sbh@ZK^5KI0bdZRj\]E]\DY?SE=;TE=C
0hNBCqmX;nG<GdNOWg[FBlEl@0cnU63`1J[9b`:[85<NY:dV<MO3B^g@HSjoLE7m
<VS=fmm2NOJg`CZ;2YOnI4gG5UUo\:Qjmk>?`kN[5SJJUWm3E[V^?c7ghmEnCl4K
aa6=_lmdYeMgSJZ;5POnI48^IF;Dp\3@ELHh\bUdVaKi7K64lLhfimD=d<i>NkgB
8`\86P_T5mT:IHEcjBN86U050?PJh\AXA8Ceh6UJhU0]^bDcHGkU;[Lhj;[m_Pgb
>d?i`lQ2]B]Vj`eG9Em]lDY91gPHn\KGVEC3j6UlhU0]^<J:aLlq7cXB\bRed[QB
[`K27EjbY>R[WkcPoil=5f6b]]=l\daGCNj5lATT=1c<\9YB]:=n7F`gCTOV^[<R
>b1XJ]^l_oUR`91WBk1eef6e@Z?I=<FoW<NWYTKU;DKWd<?WW:iX7n4gMT=l^[jR
>b1XadU>\2p6O\<U7ajjEo5fGRVl>INhM2Id<LSKD;m6Wj02VbJ9IQGP3jiXU^@H
Kf6\PTL4;906K3d:RAj3EmE4WJjHGIfn3AP_YXA_dMCdW]]G@96UmmLUdHNGEYG1
\=caQbV;;`B6]A0RRKj3E6E4WJj=IgLY7pRN5K`^d@3<PdJ:@\`kED56BXF6U[0U
eB[CRhjJmol0Y\Abc>\>[k54k]XFC3HYaVR9Li<4]=^<?SJW0jBDgcG4q@09D6B\
FMLBhBc]Xj?JAC@cAIJG\o3NPP:O[odRD7=`Se6Ga41ag3kY8^]?GI\TM@54Dj9]
lFLe]3N972\N8lTdh]XS5AJmGm:OG\]Cn@l8o9d[T\Cjo;8^E59P:f\g`@mGJE99
nFc303N97QnW?DmqJ>4jNc3B>BQQOB_mQS?>BW7h6F0_[NBiqla2ULO]3`M39CZC
RFNMKLM:YnMJn[m4g9cL::^f0cNn[d4=dW[G:Z`Qol9egIBUClc^R@kQEhMZB@6V
<]T0o?icm`D]_O<QCEch_`PfAG\6=9]m?IMm8G0oH1m_^IBX\l9BKlkVLhV6R@6V
<QBfV4hqGnbG8>j;1dH:ef`o[75TaKk=6`?UA;\FEI31U0^2R:mQemh;RHS`c3B7
>c9c1k=QG]KGmZ[dXdE>=3LX[Mca2akig:o?jhnF9Ij[VDFmOQAZXlZdF`6]?a7P
;b=MZkbKG=hF?Z4<X91\=3LX:AbE6cq`^IfDZXDPg]cJG@^50J?91XAm:kBSnhBO
DQ>0g;I4d3jYdEUfdW7ACDm[b7CfN]6`0GYdNk2kgBbe5[InFQClC84m6PQUoW?o
Dh8IhCE_CY\03JRF@SI6L[F^f`O3N66`5l]MNaWk7U;e5[IQSh4]3piZRh29giOM
F`iEOJ5Snf=Z0f]]SP@hd`H4nAM?1d49IDEW_Dioo3B1>]^I=DDU`giLCe8idcVM
`FVj2anKnkM`@6c]0:o`nQ24KkQ7NaF^DiB=3;n^:1W6ACg59I2Un<iHk^=i0cVV
b:Vj2aVb5G;kq<9F^d[^WQ>I>Kde:^]^>mfYJa7bV:FFKFUq\jPL6@c^2mdND7fR
WJj1jCE@2\;Y3OGeQkbb3ZX\fGX80Gd:T\3G3ob90;2cef6C\3KeNY\T]m1>@\BY
kdW8Gg[W5\Ao8JR_Hk0S\jPHC3]4[7SeIRTHSXdeW[QLafO=\1`lfY07]Id8@\BY
EZ4Ao4pJ2baIn<b[6TiJEUn^8TJ76jfa<B?f5U?fEOj=PB\658_WKgi8V8ORWn\T
UkPULPRJHAIgK2Q96Q_cK7]L@DIoWB61<\;kM^fbEZVaO`XS4>^S^C0_aj;;E[]^
i9OeLhSJVL@WKVg9o;GcK7]\0NkK=pTW74k;Y2SaMl]B;KXeIn2EK32R^T2]N6BY
7kf^FTf\_ebF<K[clDLcabM:L^_F@JPQb6V5O`_]_51oFha_W6@XZLbKDAjQGC`L
fV5@0ho^]6[`ikSWMJ15;M<=3NSK]EIQREVM:E`]\l1m9Na_W6>J?VIBplDNV04W
Bk4hI`O5=2hfZ:7Wd9TOP]J;0SNA@^WPJjK^:;5^H>hC;lVl<X=[5HVIilYc^cb`
`X4aYL8SkBGgN^TWFnOYG5:Wi8NMlC>7QLiH8ZmY0bO;LIG_:C47j=V3FljT`Nb1
1XE1DL8SkMCg`dJq3[k3nn_ISe>FMdf6dHE?OOa<06FO=0om6[aGGP6CCo2=j`DJ
=YkCW@W^RgM[Fj:m3j5AbJT?]edVL2^L7=2@Y=q4n<`eQ^_53lbDdOQU8jf`aROU
Y<9Y6Dk22CU]?TPViR[6\d1Z0XfajgjinafkAf84Sm;A_1^F>[T3kDkJ9AML4@Md
;7h5>49N2Y2oflX?T9S3G7PHR^e4?9@DYj`=A9R48GL9_4^F>G_3kDkbh43H1p\S
[IZ6@PY0dTLQeHeg\h^^B[cCAb<WR2c3lP8O5H;?WXN4gj9`bIf25hGc]OMlZ^\_
7@:`41k=[_]i05ceb<XT]Cha@`]dge73l2CVm@Gl0NZ=1W6WMmZPS;^SAn;lm=\G
GP1`^Lk=[<]i05DlbdcRpj8<ONlTDEZA=9YPLi41QoN[?SKfmaL:]V5>^3V?G^2@
ega5XfWF5UmRP`AGiIa8QjC`UVf[cUOY>69_a@E50G7:7Gdi[<We9Y5lQoifa?BP
>4BRTL^^XeQhmoY?hfaRVj_Rc\ficUO1;69_a>L;RoWpgB5DgA=Ned[V4:HRhPmb
c]HWUdJ7U\nS9ejJGAfMpnVnbfMPckRQ4>8oW9mX6Cg:k@5>JPhI\KEQo\J2N6eZ
gU<AJ_ED[AC7?O[WSA<E6nC<SRXhFRU]C8<g3VB:NcPVdO34P\KWI_ESKPS5mR:f
HZdN9\3P1nemC60O0a<]InOZVYXiiRUiW8<g3d4n45`pje6o7@M0IFTPTbclTAFc
JK]dL_C3ha`IAjooBe4d2c2kgJHMY\gSjaLaXN_[ngIdAWcjhfcSKXK9`kQ4eO\0
UBEVUk8PDkg_2OegWXTS^ZXTOJ\EI[YXS5GOPHRa?KQHJWkEh3QWcX6K`kU4eO\0
8W\B51q5PAfJ5]GniNHWV>[;3@oY;ZD;<k]QVXE6U\>QL@M4J1O^ZZcEB5K8oOW;
ZPG3[TR5^g:EfK>L?XKmHj3jGX?ZUQH<=@Z[Yjk>U\]=m1EFbio`E7>RTIZfa23@
WiVS[lZ5n]m8fREL?nLmHj3FCljGQpgR[li<<a2G:lMXDhdWN1E;9G2EB\_CTH^i
;iS6=YNKd_m^[>>;dj[a:m:AHNOU:^gDcU9Jg=S[Eb2`9B20PfV1ZQnIP63WoSKi
PIF2gReX]n4>EAT9`ccIcM5ElHIUSdge2HDJd0S[bl2`9BH3X?WLqLN>cKIUFQ<Z
PBCfV1eF9J_J37RQAXXcH<<;iP3TPn@0G0F^PcfNnKj7\]YoXnU3kLQ=:AKDMLml
1^99:[:>08JU@j0?RVKPdl<YTo2K;>8?P^L_Cdm0Eml6^:^?2\U]3Lj[>cKQELmN
P^99:nnT;?5pCYRF=Zc3LfG]KdW<V3M`5X>]AC?U\VMfZJacONSdOMkmaLCmeU[e
6G_HSf>JE=D^CUcFgV8b;bAildG@346?e9cUlYYhHLha=Jcc@M=X]eAVZlBf2blJ
>E1nj<\gc=PCC\J;iV09;b;YldG@FGHo^_qm[l@SFdH[nAa8a<SQ_<?>B7MS`B69
SFde[?AU:o>;=_ZWgc9]PHVX?H@GkdM87iTmkGaVB7]mYIGnX43k8WaQeq5GfB0j
1VDX_;YeM]]iSQG?<OE7\[]YjAld^C]GSnG=KYcnb_ET1ajbq>@d=kab<eelURi?
HKBToWXkJ5AcnNC[okX`BLHdf]^<c>78[JEkDC@99bG]S2EQo>I_Z]IM_TekY_O_
D\jGEHokQ0=Df<ckh@XT7RMH:QX5Nb2J<ke0iENoBTUV:NEK0>CLhaIO6TMZT_O_
D8311X6q0nT@;ZHZEYeUNh77i^fXLl^5=Y]QE^29f2N\mE2Ii93BJCKU>V9Qh[<T
Ro@]nbE4`;Koh6iEb5l]F\[o;XcH_e:Wfi?I^kdbgb<ObX2`@C`\9[_Y?[045i[0
K;GhCRnD:;W=hRU6<5ljFVjJ;XcHQc58=1q\VX>HQ4`30M9hkAHLnC25]l1GPE[Y
hSK8X\_CW0P;DJO4[8h?jbX@@`lPZi53WaG<Z8jLO?Sl:VGm2jkVfInZKo;9QD^?
D]cY91NYL0eHmeM:JaV?DM\7I[7EXG?S6l?KZ4:LOiG]:56mN9\VfIn<`BFYkqml
<AAQAZ;;X6BYXOGRMhM3>HLFkI;o1QoFfe8QF\NMaCEWNo79^V0DncQD^2G_KdOR
VL`iV_ncK2boLKDb309fdjf<V41Ui:Y@h^2F88iQh\[73fOnGjm9N4a]=?eX>SoR
FG`fN;hcPRbiYJDb30aSANJ]q9@@@\n=LN<19Ce^h3VdZB0<j8mIJkaX9`LB>E0@
4I2YB;2YTVU@2RBNjaBLR6[_Z9dhId\O?0<>1899OUO:7f2TXT_6:VRLKLLn[[AR
9WL6dN8[mPYmm>^QOGEMkD[Z29`4d\\9@05Ek899Oa65:gopiHI]^=X>Vbo4@?ZW
GX17D5lNPnGDFfG`m3F?H3J4^=Xc^8WOd]6=eB1\GT:8`HhkXh?<mNYZ6B6363kP
fBd5@4be0e>5jg4:>SDA=L1fn4fAQKilCn8m6XVHY22UF:F;]hWMmhXH[BmV6hQJ
fBd52@KeDYqc[a6jgTk4g0iVo6H3OW;l8_8[`3DCX[F=2bF;1mcmKA74om:mlmi2
@Jk[RTH6h?[ck2^P:fB]g;jd8C3GdcQa4c:7`J9=;4>k2TZcc64hKE<bHO2F9=G`
>mQ3D5<\hM^cRVOI:PB]nond8C3b^0fWmpcgKbOh77W04]6NgEF2W4M>`LV]VfdM
hm?MfGh:j224T?pl6Nb:^E<a4:TM\];RGH8bPQ6=iQn>8VgB:Bdn7Gk8[BBH`C3k
7]^DAd;SN6EN>3^l?jD`P9>0QZREa?k^71G4j>1?iO3A2N@2:\l1I;H@mOQY\md7
m125N;@IC;i<>H]l9[>;PU80lBKEa?kLQn3hapI6QWZLUkSHS46J;Wj:BU[CBFKM
AnSOmV2M2L>1W:RL84mYghFf0Gc8Oik]4:2joTI43N]lXdXH5Jlo6gaaaLA;dj@2
PP?cclbMOX0><YYENkS2mO^en]WbLdfbAdmjJJIbF76lZKXkcRlo6gbj0EXIpkGW
@I8GUbGP]6M\hIdEHAfG17Z:KHN8hdDfTJ=5WUA0Xao5=WK5m>h2Qi]NeQimXkFO
@LM=fhGP2_h;Z5URSbSpcoS2I;=h1?<a=T9NLiYW0:i2`]8jeJMLhPSjT^OJjJ\a
XjBn3`<GEIOR_1cd>BAfcOk96NeaUkl>7QDif<8K89X65=XT5;V>QP6jCgShGiQh
Qk5m\afBAJ0hH6\ANBmechCSDNfQUkoZ7QDiMmLFSSpe<PS?<akRGOlN`[Q60F=b
oKX@GQobhHF@Gl8LT1;G6aP]aL1MQ^[A\h[8YP0]Mh=eg=WkFSO8>3:7Q4`OaTbi
glWVGCXKKTX^GE3YlNeafLK>^N_CB:G5oo2nZRJeMD=eKJC?F<I8>[n7Q4`T;C`k
7p^4QOKe<=TkHRY0c56fa7VLefojfi[`8cT9gWaJ_l<cPd_eTa7a?jBhXeaak^Wo
<j^F2a1l9MfT32DLK27`>BSFU[b7LB_6KZ>94H2RhYf<EC7Kd>ITm:Ma4fXeO6Io
GR^F;3nlPmfTeGDLK29dX[InpQ?FJ0=<:?M89GlZ6]DOC@DIggej]KnjhR48\?Sg
Smnfo[`MlmcB9>ck89YDZ[;baQ4]LXPS1ERE0ioAZj2_;bUIH`JNR96mAX4c[_dK
ad5DU_\[6P=M\ZnPWWR@Lk;3WQc5JoPW`ERceioAZBc@WBKq9DjeJD;mGS1[e`o9
ESN9F]AG;`h<P>TkmCQ8h3RFg]ZXlUb2ZI8ZnG;fXaNFhBF4q@[iY[_nAHfhS3gF
\MCC4RAg5U[a_@n6Ff`S0mF4]]lTYOB>8L:8OC=^@]eEXJ8aonJ1[Y5Xlf[S9ekk
?m<hJj^LOCb<mOaQXJ1coNJ4f6@Si6UN[6]Q4[lL5V39eenVNIJk6YITAJ[gSekA
dm<hJ^>ibUIq<JlVXIEhJT8`]5H<3`7PW6c;L_jZM3TdFGX6=JVS91L@Jne=9^MF
_GZS;_d?Uj@=a7>aKR=7fD2g?8lXToSTbgQGi3hMmnN5mYIN^ZV_LEUkOQUkTmQ4
6gUKHTe_TNm==704KO^_]DbE?8XhToSTmOMm;WpEJUjiN\Kc5g9UkHfSmIj4Ok5c
bidAeF27546[6X>fkGOZ>=?SJ3a58m4jF^Ql69_a;On\]ZSfFVI355HdN;cV1in_
YdjE_jjVN[h3f]i;aZNH8NkDQ\Aded4124349F4D;Tn\<cjIFj6351HdN;cRg[UA
hpWgW3L25?Ic_^DEUKmDbaQX0<?DQ^APLP>Jem;=KPo<H7V`ihbIU[fTW41MJm4X
B0liIiWZH@ISKFZ5L3RdYW4@eRF2A9QO]4eUiPY^^6Ul2\hEglj]mM0hYS9dP>SI
[GUi?VWCgUJSBFZ5YaRdYWM1h606q@lN?jIMA;<N[QAk?N0TkCWFE\WSnVjTk;KU
EXWMZ[fCBS8=13jZR=]j\F5Y]kKU25^S4iB4UFQYLW=>fJMh3iWe27Lbi41lhn?k
DW0Sc^;A@k8`_^Z22TU9A7^;SElY8G^=_ijcABQLfW=4fJMh3<V?_<6qYG9EFLFP
<ZQUidj8ieZajSm1T6PQEBRN?DE4[1b4b8NfU`Egm=mQT>XmC6e3Pc0VmoF:A<\4
oP1S^_cWKeSnTaQ`^\q[5XlgW=h4kYWfl7cgLbWe^hE>g[?]g2?ElenneF>F``U=
1U_T[DORQ9hXV3DkEK6Dkn2mo?eBnFmjmiPAmJg^3G^U^7AWEQWGK\3I^7kVdE;E
a=0XT23lTYo_oh5Q4ii0k@XmFdlhnjijdGKAmJgAFNZMSqI?<WgP\C18]Q6FCaIK
;ZFA82;@Cgfh;6IA4cBJ0eO29_^mG4ESS2V^833Xa8j@k`IlOnVn7D@D\PaSGjd1
l[mATXcJji6?IASA7QGVJa9PJAh\kLDU[GCRiY0JW^@@SdIm;01nj2@b_1aSGjUS
ZN?Bq`MS7F1;S[T?KhH>GeYmCbenVQmK\Z3OlSLE4=G?PTZWSM=6^OR49fAh4Q0a
3f:@9`]50=>E\`mB[2bRWZQm`UXS=S3FSoUc3^L=IZ3AP\<lS_V``7hWMZ@SHZ24
Wj:YU`NXc5>CA`I012bRWAAKS?HpJgQ4IK2mj549BmN98n5Q1Jd:V_;C3AZqEoQQ
QL3l;1XoN6jA3gbjhPX8D?k=jIb5k8U7^Y2gS:jj89RP<8HYVdgN5@YN2Ui8QVTF
Q;>ePmH=Y4m6@G?9KW1Xo[@S9GaKZoUC?4Nnm]Pa0mT[:jR2ncaTW]_`2<Sk<V6F
Qh7Vhm40YA=0@G?9XOhj8=qQF7W@Ib^PLXb8Q``NXMN\>IQk0EL;8=Y7Fa\2JJd=
9_AS^CgTnXdI6O[h^`ZZi5<H=l]7AXjYfLVbiYXnCj_Q`THVMnU^JdQ7G>kPnJHj
?2X^^j[5>5A8INag]07Qe5Ja=eT72`fRf3XbGIInCj_;GcYUEqg^3=ieNjK=Y]=1
E2;<6GG[Xgj8kh7`QKoNBc`Z4eBDT8QNUh:Hb0:12mb@g8?n=e\Om1ck_T@Y5Va1
_8HEVFbhI`fOC1jN7MLe=YG;Q7jWogIN6CnP=fYW4R^4H3>DbNEO1GcQ_^iY_6aK
JFHEVFhXP5Z2p`k;hHhEnP9jMoXKHamP:`5=eoS>HVnWWfRSMTFV>0N;ZV[fOSCe
lMIFNTdVqaCQ]<88AOI3@VfSHEX4ODY8S7kfH^ZWk;15Dma9MjWjES3OJ7dL1LVT
]8l5:7LP8K50R9RM;iR96lYE[G_k6BUDnR:aeM[lWEHGf:81ZKhkO\U4;81FC7B0
?3`5Lml[3f59X9ARY2RF\lEQ?G_k6ZV69eMqP^FW^mM=7@][2j8^T<:_1m7PgIlX
nJb48IXl;9EN`M_ekG[kAXl5o07kj9IH<Lo77A_gHS<^9HGF]5Fg9\^A2B9RbU`Z
XKKO?QXe@>T]CmmlPjbLLNR3OJo>8[<a8E9UiAhAH8=LYHYo]c[A9\^Al7T_fdp?
\el1O_`mhMd0hB5_n_Klji@h^OlgHcGPjR:2cNOCCcJ<JaLH@bHPllob6AX1nK[^
boOGSO\>giSb1LMCRL7omBHZNamfbKVDEUE\INLg_^W^JY806[6QgK<bmoi;fo@0
bhJG1hABglIb89[CRL7]e=i[^pd<@57R1Wl?dA@1L;8m`o=o>NXgNQkC:HFLYVl@
JQ[:4E2fEA_V353:CmF56G2FhLMHJb]K8PNJe9K3?ZgT=I;JZ\CnpjUoL6CiYgbk
^WodKIN82Jj>88:?`cF:HQD0DiSmpUEVh?2qZ;mOODK$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI222HS(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
5\ZImSQH5DT^<R21::NWAOQKZnLbS1kR4f08T8o[;UPDNK8`o;>1L6pKD:c>Ila3
0@Y3>Ek\i<;]CW81ZRF8YF]6mo`q=2VmJTP1:0OZ=4JK2Y94ON5A][Xb@^4pGPNo
3?pe<1fG9IeV`N1UQ[aQ9;`Nf0AO7Sc3T0gKGqR8jiAJIg8`28VLJVODQLYcCYG<
oNiDf7>?q@gWPK]bXAD6oAFo3FLQ7_m<N0hFiZ^G61<0_KEZ60l0[QojO43[j@>j
XGi8hjJ52PfQplh9@h>=H;KmN2Sm227CF<nVkJkcl0m[9]gpg1VYjSXBKhlG\3X;
Y83^cERA5jInlCmbICNa5l;qiEc2I3YpeDi:Z6q[LWA9JDBC_TD1k;2B1Jj7]UZc
jkfcb_Eh72?@H<Gm]SFo7IbNoNCGUBRObXAlB]Y[Jf96II;1_ogg^\Jd?Jn19:ZE
>4IFHT0\7?i`ZiX1SO08Ve6CHUZj6Q6d`TS\BVK[```fIK51_fMg^\JjaS0R7pZU
5?THfT1VM^5T;C2[q\fB]IOV5eD@ZoohOiMdn6c489?SBgm>lhg`3gZaA5o2^US8
Q<EFm[O@gK6D_fENM\D:A==NkVDI^EeOD?cmFGX=0@?LU3d\R9g8J^PUIl<TmdW@
enj\KWQcoQVBA\E6@\47MM=;GVD\mEeODWnm[HeqYHK2QKFNXgK`adf:fZNTAZ7f
_So:S`2EKcaGMd^NdVDD1kfD<29[>d]o[I6kPJ:`YkH:F=1KUgRFo6=3o;N6gdEe
kAO^MP9Djc0>GJW1QQFkD]klnBd75LiYLCX\IJ0OY]>XI=GXUg1no6=3U]OEGkp\
gE<mL?1ia5YnI`]K?:j\6JA`@Snbc0KBQ7;B1>ZbA@d?U`66\6EEiE^QJo0cS[I\
RbSh9i_GaD@iL_Pm_SV4G9mdW=3bNAHGQdcRC2BmYOO4_5hfR;UQ_`L4?3NQS6B\
TcR:9Q_GaediL_PbHVNK8pkBf3]bjhGkR6khh2_=i^5UY>B;mZ8XS=^[WSY]h>HY
B\HJP\cMNAON\:=LI]8Hd1kbIoKkjZFkYnKb>9dSj@i<l8I6DmnV4F7[Ub;F\;O0
_l]ZcQ?IR6jF8aC;i5?Hi]ko^2jk]ZFk1OKb>9J8FniXp4jRWl:?ALhm9>h`9Fl<
oWA5R_[N4NA_SJlR0GoSm1jcV1`BVfoIao^o<iV]:?R1K4f\7dH[6NCPl\3m`2D1
_?eYnjU1N3[W]\l=nRScO89LE73RBoU2ci`P?N7L>5Rc>43ek=HiZNC=V\3m`Rhd
X9CpeLH0Ec_E7@cCIFD>SDBFc?[K`oMaSN;06^gf6PA@=MI\eBij\l4Ri8ISK[Ha
[iUfe1_Df1DA=@6gD1>n3EYZ`UU7Im5ck<85[^kHWan0YO?70HWeMYlo>6ZE;GWn
Vi\aeM02E1eD=@`AD1>n2nZUf9qkPV<kB`l_OljWUYV:25L\KUBNS06eEC<3DBQN
MlVCdY@3Hjk=iihl81U<A8<9LJWkWoTmWi1VO]W37=FPf7MJ;bM\SLVbZ2WNDLUe
J`glMMaIEjLjUAOOURAEBf;CL@VkBanhW8DVOJ^37=FT\?o@?q8]0CEIWdZ>AR@W
^6H91kkFV8X[h[f[LTH\J0EfgkNSO2bU0ZeblL=UO^k9FT=EWH8Tb@?WNaO>YS^E
mU><1nF1f?<X_UaXdc[\c32DhHSiG>M^ZH:VNX_g;YJchVAE2>8nVNKWi5O>ml^E
mU7>2k^1pje5l06?[oBa65]j2kYhV]kg\ljl?\98bTMiaH=IZe6Q;I<Sc:P1nCV7
[``1iSX7I;3N7GHq=]_iU6^MJmKQNNW_l;DE=VG1_Y8dR7Mj=V>^R>M8cc2l2d95
U_^KAC`PT_BXo2i?=k[idWoeEm4SBknGacRiSdpKJac1JZlTNhaNU=JFL>4>kSZK
S4_]hNHFWA[aY8aJ7n7geg54glHD`9I<:=iK3@BKEiW0@j20N<W3g3lLN<5PZbTU
SVQUIUdnW5eU`75i6ZO2cQY^PJUTiaEaD>\@3RXKnAf:@VG0J8D3g3l?FQ\Ceq`]
^4UW8?6>Y]ef<NFjWPOnaf?>b^Dfm]eaBQgE=_<jU1_2@WmP5^9oHo_j]3::6I`W
J`;BCAY>8nbI9cY<PaWUSfb>K7Q9:Ria1TQcVD7L4lI=k=bg@8<A@6GhnbZ:7``5
H7JBh<Y1ZkbI9cUk<\?apmh8Di^IR@do2G3UO_U:QPTKPB;Q^Q@[3il8E9d@k63R
jW4UKLO7n8W\SQJ@Hc@f6mj9KC:eiUd1PnU`ZhEoAJ^k7A;<^I;93Xl3HK3gZ`=m
8Qn@>H4`3^Y[\9i?Y[@H;m;OYA:iEU?l:nU`Zj_Fc4SqQ9joOam<`TAILB=i7C5o
<Al@:3XXhP`SD^W]Z4@O[n?16[H_Q;\cNCF=ao0V[g8dQQdWKG?HTTKeWS[2g203
m7a042<gj7AZ^^j?1janBYY0[TDd:mQ:N3C0:ARIYgHdQOm@\G]<TMYZWS[20FNW
HgqiejHmJ_?oU`MWKmHP3dKSk3[LiZe[ae1Z637XA84L9fPb>WRLiaM@H6Ala4B5
Wl?iSG0L8j0MU0iUPGnF[:k>=5EJTL8dPQ?=6c5:2DL]L>@3;?2MXifNg]Q^UR:i
WTbij?6]8E8Md`YUPGnGlZ6dkq1@8l<cTZY6CPIoGkEkbciXMcY_fhiPnR6\jWCk
WP?XKQ@RnWa[7:SX44W6i14EJ_1YWlFY^YB6W\[QXk\T;S\d\<TC]AVh`de\chZX
7HOQegQ`;MYj52P=9G3BQH?EDj1P_FoY[YBBI\[QXkSl@IXap8<Ro>P0n@\YB>aC
J[6PISaVmNKgkSXB:L0S3bP3Y?KmN@dWZK5Ni:fZHhTll0Dgd8NU_HSgbd\:TS=m
;LH8XXJVX:gKWi^];>0G0EEidLLlkIPNKH:a?@=I5_0ODkDYe8:Ko^SGKdF45S=m
;Gik8JBqYKBYbTO69=lj_cKJ=9VdeUO<KKTdeOX]p_IhWBVC8aAF^fk>Oc0gNEoV
L^DLDGcW<>P9@FM9[bmZIXP:\GR7V38G6U0<X?GZe6Be?1ZdA`i:Ve96m]X6Ma[R
3;]Y]R=CS70=XEoS`<G;W]_R3R5G2ojEHCVSn1gX:QBZ11`=TLiD0eEB`]X6MeZ?
POAp226YIiH?V1W]C]3AIhjC1D0f]jRQZ`4>McVUZ2T<]^8nL52`Vo:Vg0[nXLb8
_JoQ2iZ1@XVQ?1JUGfO1@;QknGD]?j`c4h1mLc@UPd0jViVU4X^9\Rf2cS[M^i_4
OJil2b2PiXf_?YOmGfO1ZHa^Gmqld1cfFUlmFPg>GIigLo@WNT:JGSG3c\5R2G`Y
HS0RD\K7IWLYP=;P5CJ1KXIZdoWljILL>DnDF>7FU=Ph[m4P<p;F3f;Q1DJ^S^Cl
?^N;nI=E2MOGa[V0NE`bh^Jdd109fTnaDg^Hm?OT4_SG51ZL@b;BSnonm33TDJ5H
STIcbO3IR9LGZKjb\a;b?8bmAhSjZ9j_I_OIICmgdkRHiXWLDj;29ANn>33THb5H
ST]l]g0>qB>3F40kP;KWcc0RlFOH22\DO[\PF:4cfE0][a09_3WjSPgF[SH0<8FG
2keO\o5bRC?jHZTm@MU<WLSEaMS``9?8`ni<S8S^;=^MhkDYk@all[TFW]Ka]N1n
Ih0NKH^f8U?HmZi13UUo1LS>iMS``XnjIa>q[8LfYhGmGch^7Cm@8<<DFb:ACZb?
[a76T3Qn2_d_N04k<MmlVoV[X`7oi\BY=DR@7J@e1C@S7NS6[`\DPKG57g3U1]DU
42Z]2;k5_`d@k=`[GfnFBh\^lKnJmM_^:TliMJ]Q1m2>VN3Y[`lQPKG5LLb2fAqD
TZ0I[n00Y;`@cC8^>D3D7?2oFZe2k>0EP8TCRP775PXT=Y]Y0C]L7>KHEMHm^BUD
E?\l>bnX]T8fldIX^5X\?5[:`V4C1Yj>PGTlU23QTW:PSZ]9^D3`mBimd@9Z^1cD
L_T7>P1X]91fldI>YP@QTp[>0S@1]B6GXT^bK0Kd@aQJdBBb9KWB]I6HIf70[Jfb
h@J3?hef8QJ29`5>LHEYFI36VELHh2e;iEja02O`C43cU5N92VD=fERIf?nYj<i\
VJ[eaa44KOP>leQ@PW1Il7l6AYL^XV\;JhjaBbO`C4=63gf?q5El70l:a3];X[Bp
JYfJ1[iDcQJ7Y:UlQ:[jQ8?`6PYnf4h0<>9]\ZhMPULI8T33Co:9NB@fX`4hOaid
J3EiAGQ<9:HXEiT60;DoHh3GW69[PZP;S>_\?^J@3LZc_UC[NS9MfBXCGHiSBaHk
Jdm37Gnn9:PGEiT69L2DfmqBcC6^EWhWMGK=jHXXDfDmI_oNI6MO5WZGMLYOP]4A
<If`DRe;VfOV;m<U470?hLOB1EmBj>FMV=RJCDBF5F6SMYQ33eTcm\[kM\[87QiR
Vn8BA81m312:?BE==gbGhXWBC3^fj3RMVXfJCDB9G9XaAq4TX\>7>VYSeJLjSdoK
R7^hLkf`F0HL1Ad]MWV6lBGFU7\[F>Im]:CT<HGWA6Eack44:j2AG0[nd8\lmD@b
hkGWJZmFJZJGY3c]6OM56\>D1UXe6PUYcGd4QK>P9GCadQ4jm2]AZO[ne7\lmDCM
EY0lqM\^eEUHSE2IT<[Z5NCh8nPbNo=SCh3R5;?dH\26_b\^DNYmVXM>LL1JU5@P
kWj;FM;Q<J`_?IRdhVLoGC3d4nm?HkEfJR7A6R?dTeANDmG1[b?PD=HnbghljBkY
]BjVcM<]4f`cAIRSAVLoGTo2H`^pT@dh\@j\1OfD^Z<G3=7d]6:BRj6N9VF_Pe4j
YP5CCbnFEg=R0Hgc?bQmC<ec^O;^T4RTPFLOce2mJKT_S]K[R^pA5lo7JgCMVgEW
GibQ^jZT5OFL;V80n^LHA3Y7AcZak<TS_hT:n1=m?67\3PVW9>ZANgDjDdjoV2jf
2ldZ;eiVj16]Hh^99NO[AKl:MY:5eP;NQXeToV9fg5A2<_;g9TgA3iiWDn0oDjHf
2ld5YYmVnq=\<KFW:\`E3UPGc2S;cG_@3bdE=Ec_@@Y:``Ql=b>:93adI:mdEE[V
?TAWj?HV[[nbKkC\XVb^ldBNR`]VJIINO;\;7DKon1801L35=[7Ui<A;:GXO<E^f
1nYm0F3mbaRbEhC4;;D^OHBUnK]VJIT7GBhkpGEY5AZiPThBlLCCmaZ3>W:`WT0P
oG9nA6ZT0RPdmi[LR[7>bgS=AMU?m]l]ES6BGWECGMa8b0<jCoV9M`fF;RVb7^oi
TEeUl7co<k9ehPOW6TWU3id>A4:O3<^BT^GZYRE4kMjijf<Z_ojVH`fF;nW\QABp
N]KmL:miUL7jEQ>d4HF:D1X2nkZFC1gfLXNci:U>[T6NYL`PS1pd\XH:8bA=TK?g
D<o^=Xd1:Eh[_2AHeQldM8kDT0hbeg?WCmPk:7PBBbO7h]K2@7mo1f\G96SkdYn8
]BG3^_lh52FJgOIhYh<F[_U9hVZ7nhHmFIE1\?[Z`Vl4APkYb16J15fGmId\dWT8
db03^_l_jSeOhpJ6_?fTmWSHjn@^MIIJn<cA]P;ES=ZXZQ;jn;2f54FAZdS1LH7P
@;2DcY9Mdj]iEkM1djkJYgL:i2A[nNoPJ?9V8@JBJO8FY?AlWK<`dK2J_oc1LJ>i
;]j89`kDCA;IU901:4k6mjO:oTAAg9oPJ?CY@ZJBpPK\_=Fe6U\med0GSZYWPZM5
0ViBX9=oVRiRX[=P=aPD1KDF:\3EHif?e\[[_4=fMQDShlAS`VDUcD0WD6K>hU:O
IgNh=C8RO0nS]R9`O\7Fo:c`fVXlDG^[9QR44]cJK4D6Ll_S0GDdWD7_k6K>hVP:
\Y6qJgbi<h=4m]o<]4HmW6TXYcijmJ2140XGoCAR564=f0bda^9KiJXM5F:907hB
g=QPJ_aGdPMO=PFYSjPHX3_=[;j3MRfmcgUZ^CkUJWDDiWg_L8aDM=Ff?blAkQgo
A=SPJSn7<P`3=B]:SjPH;P:__0pj1m<6[Ini2On05FNeX19eCLfJ@;=1ZKXoiElc
]3RgnFbAm2pUOeGRN6kAQ5mnTI]Q?aWd`b28JWSh9\Xa@9JC8`VLZh6@9n\QLXRn
X3=c8R4NJVJUP?8NIF^3K@?BblWDFPj2XOG75[8LO[R[@nZcY\d=TK4^m^OKC\fh
QYOVLTCoJUnUP5khIS73CcoBblWWjGZdCq^6?LBn9A]U1bHQ^h9_eOA`gmh?h4;2
oSD?^0Q;F_TKUSHGmELdIa6a3NQIcOcJKUV7^E<gLMl:SMABacYVj\hA_MPmRhFL
QM9CRGN_FlJBP135NGHoaV_6<njT;3X;F]]7XI<Pjh6:[IA]:cYVj\CLZ[HQq=J<
\e]o\BWZ_`7]d4B:HF^7_^9UYhC1E34md6C=naOi1g5T@Cg7Fadj><Qj^c0F_Q^K
hQ77F@bVIh0>af3oB10298aq;h^WGBnR?G2VF>Gnf[W]BFJ:Dd4;AE=PeKFcADmQ
T];QKfo9j=D?26OgYJ@KXD<F;W;[01jSkX;fLjL=H^NlEeDF<dnR=B3R8K`PFl5X
<jdO5JaOcX7Q?iH4jMmlDD>G;QgHj1`AkXCfLjL=mLPd3<pHZdS[RV1E:fXoB^gf
:S:MX<>Una]HmAiaZheKeVf7JX0iE[nUJW[^4Nh\BgnSa4iH=2m7h<UoDN_:O9hG
_\ML8YE2NZTCgJ\SZE0:cg@oT\IhMnY9]>QMX[@[hi`gaZOHl<]Sh7GoDlS:O9hD
EE`E7q<JlVXbE\JT8`]5693`7PW6c;]_j5M3TdFGL66JR35<X5mnoOKM:@]2N;e0
`V3L5V<EVG5\e53V=;h46]bHRM]O4:3fJVWAcbIGDlka0FUBFG>5k9LNM>i3mJH;
`XkLE5<c2IO\Em3VG;h46]Y\bWI<p09lMlSMiF2Ujci8=DfQBA;5LI]DMgQ3=Fca
6YHQ^_EE:2>CTUcWdiYqo2@]ERPiQCEQXAk^CSA39<llQ_6k=?bGbG[UB[\1ZiN_
E7m5HGgJFMS_@b8bDKN@o;M]HAo9amJo?c;TXP@fl28J>0YiU[o>GGn>APBeaYkW
Xf^fSF1LfB3>Oja5@K28oI?ZUA5Xam:X?c;TGg:m>7qXRN@@eekT;WYZ1g`o2Rkn
9TX2X4odWJ73kYAgK1NKZN1cbL[GkV^fKn;k2Uc7ESeLE=0<B87a=hf?3dD[IeHk
eZRmG_ZZ6jV63KR9H11ImO0@M8GYbBGNoiS@:eCmGnYEElY<I;QF=`o?3No[IeHX
\>^XGq\YJL<OEVNIgEBdQTm<ffecGTK2O\NC`9Pbn91;k3CnWGdK0CZ_FMgeTAbF
><KIPT2e2SkLSLnhP?[Z8_R>M]S;a1\`M>]Y;8f;1lN;BGV[ZhZHb7gn>fJ?HEdS
ZCR`F59eVCkmi@jh?a[ZS@R>M]jeE08AqZVAJYM`0SI;mS4l>EEYi8afCa4H]PPK
F<mY:]<XVCJMZ2fKX8k26hk<F19XWlK;WONf<a5W>eAfW]O\?5<?5in525eUbbN^
;@\oa6V\@F6bmX0U1a4lSU`EQm3e4`Y1_8ND;a7Wm_AcO]Oe?5<?59\1]UlpYiVb
;WWPF@ITXF>^MoL9f=o;GSoe9C9ATU@Y>WJ]9oo]_Y8NiG^IEGHnX@lP`_BGfOWR
H4:CfH020n2=Kk9]_AFgI1RF]R:XHI21NogP_<?l`YdJS[<5aCQWa_c<Q[f_2OeC
H<0\mHnn0n\LKk9]ZYOJAep5k3TH><?[OooP?0j>]1K4^6W1aMU1c;;F]9;OVcHa
jamTkQ42PPag?XcafAga4FR^d<nX8;Q:b\`><eOAEO[TYCdD6dN4YSU]aUMj96of
`VF62W<iP]65eeE_3i_a;]_nd2mXH<O5b>m><VOAEO[^FZUheqoS13`VQZ14[4[l
<C1hJ6gC@5IbFQ:[1V4F9DTQ>ElfO]__32_H5KhkO75XJX=HB\o2i?=k[idWoeEm
]CBknGac9TSEpSIGBYZ=R[fKa8TloGVi09<lNlH43]Ee`R17b:EiAXd75jMEn0CF
8oen;ShegR4P3n=NPa\^fKlGUdeE<BPYd7oLo:jHT_UaBl5C=bJ0;NNZYeMamB_k
J6a9bUa2CCI:a6=ONa<ONRlmod?h;BPYdJ>kJ=2qcV_gkKfE37MPhfJIB`^IF;UY
6[TQcT2ko4o[aJaB?0I;Yn[L;1k@jXC;KIoL`RRU0@;_Fh8GNg\8PCEPoj2U[ob4
2_D^Y>:fh>4HIXaoi;XT9QGg`KV?;DI_Rg]RH@YI1@N5FjQTmgoaPo;6oj2UObm0
lBqLEL^XkH<ThoYdAUi=m8kRWIgg:]>S6Z3l6<p]7d2_A`h0C\1PS<UQVUbMj`i5
l6VEH3]a=J`f<`DG4fH9admPMVZS6OUY6`1P2dD]mYT6@f1EL1:VmhmcEaZn0Qk=
6k8L5iI2=:eO\Cf[kl@akj\\I=0CGm4Z]_bI2f<]?[=J@MmE?llVmhmc_ZcY:qQh
OineoGomYlFj<>6;iFCjE3I>XeSONI9dL6`S[]@6F\^\BC^0kA`UdblTWC;3[9:S
PFbE3UUkAknmgV6faRbT;oN40DK0A[d97D^:Vg\EbZMi>P^T3dI<d]Gf1A_G3NPS
1\bYmM_k]Qnfh^6faRN?^:GKq8I1ET4k1BS=gmWPlKZ6Xj@VP7H:Wl_J?:@Ga9n`
IR4DbL]Vk9k3ja[>9PNm3SEH3Zi0C:GW0>GNhESX0a;?ZU^U?j04QDi;=W`3WkZ`
6dojF2]<LD7`6dOHn=o=2^;`YkiQC:bnkjGa3E4LBa;?ZPZi`U6qWV:G4:g_c@;3
N=N5?Wbi\nERBbKAfbZJH0F@Km7JJnS3nFlMbVbbT9WPV=kVMhB63TUjnRMC?o:I
jS8QIfl]>o9LFSRQYhS_JXb36U]cn0HF4Fl[e\]mFRFaR[IbD7j2_T`Nn\877oU2
jkiZIfl]GnEV;Wp=9Ah44IYVjCIE_T\=iM@2FNNAg4mIlk]XbkE:]6hHEg4_o@mo
_DYI3EgC62\HWMYJc?oLQjH9`M\DH4A^80X>j0=0GKoJ?N9ddGebJgM4AQ<aIPLX
ne\Pf[<:B@IQIjoDcl2Laj3H`=lD8VA^80XY0`]RhqlREA1DoFPX`ATY;1;EEPBL
1e6ZCfNkg:>9QX^o[^Io:G630DBldmR]Zfj@oiKW3hXY5T9JbU_hZkFD3J0GWo8D
e;LTkgJo1aS_nP\Mmf5;F_Bm>0EWZd70PVh:g2WFWK7YYT9ToVhhO=FT:I0GWofj
3]>Bpl`aceJ:=oaOYXKih5CD:Q:YUeHQ17bI^jCf6@FPcB>g?G9PQbjAKi@dMOU0
R6WogE@FhdZ]FB[J;ACZ:WfR0oe1CaZl_Qi\ZTF=7n]S33i][G9:`hm@86QNaEZ?
DVTADX@96df7Mo[W9Ah^FWfR0TlEIAnpceN^hVibYI7ld_KD5A<<:C@`oc;ZGNXU
051GkmLaRUnZA8pZ[I?U_b;<DKPV\WW[9o^eh19F2RA<@eTI=Hd2GkOjngQ>i6d5
`26mkkCP\b@KUPDBaS\6aobc_f_@_<jo_Q?Xd]0mApSNdEKQq[Z3d86=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI22H(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
bNcd]SQV5DT^<N]l2KfH9P`77ZmHMHNiBeUiU?=87TDmUL;g3g;7;OO6UmOkJKWG
2>Gp5k13gOiK9VY;?b2p;iWc2M9;ZBF9IK3opJlVgZ0qTOW`i8QKI512]bbdEHXo
o>@E7=8`Kfm]37qGh_hS>MNeWYZ<5@88<4QPWaWX<><8ROH2Bp[nd`T7a@9IPIbJ
U;QSWYBlHgj4]:]?jQpHV>BYWjq3UGj;1pJ9n^k`24`3YTegaIEIfLYKSAMBp]e`
jmUo]EHbAdgcHIY]bbC\D?F5A@F]EZO>DN;lUj0FN9hV3N=KgL]f3]7\562o@]Qe
g^cYDjHX?;m@A584NMNO9VT8WUe?GmO[`EYKnkAGR6AJU>oS>oQpXY2eUfnXbn42
VQhN2<`[eWeG7_WDQ=DP1Y<eUnP@HJeR7MRJ=eHR6KU>CY;n]?ZKXLFVCOXP9nbP
XHRREK`T3BoSa4Doc;:AcYJVmNLTC12Vb1l@86^O05q^oHo3UlIh1e5^M6RSi7o0
]3>_W8;jQ]6=23`aMK]W7;RnlJC?IWV:[oHF=4AW>NG^]2l4oBn?1c9mWTW]BNJG
`3210k=k>bkX2Zh>@0kiT6EA68H=5E?iSpAMSU[4UiRkl[G0dYLTTZiBoIe[FWlC
h<fE9``bOLQ4C@kD@8llqj@76YL1mTYDjjP`@89LHbX[9JYh1nCWN\PT;_fGd0XN
I>VB4b8`LX^\`cd9R@G3<j=oDPFQd[Yg\Df^F[mSS3cq1D^QIh>j_JL<Mjj:da7d
8N5CbU;ARD];><lT6kChVk28@k;V5C:SFo^2KZ7P8G1F1H@S\3d:cJ8e:R?4fS^W
mNWdo_n6jIWS7<T:_Qj_J?h_@Sfk?b6;6kpPe=FW0TW7jedhmaHKFQFAJ^N`1eZd
a@5>UgUUIZoaUK8Ei@<:B<_n808c>SWNZQEP6U0R^=NfjYLiIAGRf`QNZcTZm]8D
A:g@Ulo`;nQIn?YI`BlNfPJ<Sp0OiQjOKPU?W;_=@iY?oJQ4eI4MIhNMfJ?lLjN\
`_CPg\1\>om^e@O5OfFK7DD=UT09O\hl0Zl?eAJDh^k:N?boICHkOnWc`RHl^9NU
[^nnPfN?Gh?cTBVDqgiX\U7E6<NKZQ^AK]Jh`cXT8fkYT^MEhSOEe?gD0<HNaS2n
G7ARjnSE7IcNQbfWbgTD<al798NCSYP0G=_aBH7q\oi8o5lBQ1=[7:CCdjh:e36e
Z?@hfIN2_iRd0UR3RZc3feJBB=Wi7oC[B3jWK?^O\8oXmKjo;d15PCZ0<7No\D5_
B?a4SEJfdicC>3n@Q6QeD`]Y6kTneXqdCl^oamO>b\1XFGhnHR]@\\6?=k6FF5<3
ARFBk=ibCAao\65:[N1]>\nbH[D4H4DCoqU\4JE@W=PHBM[Zag:VE3ZM;FYjA93N
1^eDdT0X^K6gPRejXlLC^QdY^HA4iUT8SNU?NE7fk\fTMf>?M96a^1n]`A8LgKU;
Ia6DRI9AdXbD86PVVC_odP\2phTS?^jl;19a<[J<Yf@OJhJLQoD]DhTU83i=DK82
YINE:2K16LX<U=@DWUIE=4UiWh^HVMj[b3JnGZ=fLahGeVo<k`GOhAHfJ7ib>jVH
H`8GQiDS8OI:HU2qiAk?^>j[^:ElB_`?DPiGBl5GOgBFZfW7JIdAOlHbH7VIlRb4
]cmFLTJIanK1fBZdi2fB\N??jN_@bZ?gKZ[8P4pTUI8dLDS:aGbJ]I61:<gUP=Bk
MR?CKH2@^MPb3RFU8IkjT==6=MC^1;2I?4cWDagT<Z[X=?S0k]29iiHIgLVFcm0P
<NnE?Sh5^;TfdHmg>:Kk^cL2d803Oq:oW886X>^>gF`=M5GCS?fQQhejdj0ja>eF
Gdbg;=KJAL0RP=P5ldW^^Fmfj=onRk::JWfofl8>^7491S7V3:3FLmFWLl?_3k_F
ADni_:VkOn4iK\1SZY^Iq6o@o[7PSP4YLk<Sa;X`ADX67E:W9G_Wd>T[V4SV^KJh
]dMKagoiJ=EDIInJoBU9H6>Xg>Hia444jS:dh_:_=0d;ANa;COl<cAT8kkcCZ`5N
n_dWLa5@c[XqKZ?e2fIKE@7QnD`S47ZJYD8TOHKJ8E?]07m[l\oNL6XaBnkdTXB6
k7FGJ?K5SgY:KL2XBBj8f@IVA0Y6cAJ=7KqoiC;FKqO:[>7bS$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI22HP(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
;aKlLSQd5DT^<h=`7m7V^npn\\M4A:X\CHAEKCKg]\:WTN9_ohgYWU37J2GB5\eS
]D\^6Z6\KZZJGMeL^\ohIQ<>Zeq_d<So5dWmU=XcdDVkF1YL@ci^kYNGkbK3d0a<
S9J?;LT=eaqmMN4B1qn6iGE2U;1=]j2LPn<6nlA5^@?=E3^<@HaQpMR?Sh@cSV`@
j3NSN]Q=@k;`^[]IK8bQ4j=pc<X4l75f?S4TIR64?3DaCS=`6FdZVj@7pT`aL1Eb
3bMcdW6L2A[?eSbG>jPiKoWSO=N4:Ya;]pEV0gBJYqk\Ohj3qJgPmJ@V6cFUQo5A
kckD@H`k5IGIP`b;I^PaeM?2DP2L2[Bk@_PmN3gJDN2eo]nUKJhC8:811QFjkPJ<
<<<kgI>7J8426W0R[PP[Mo`CUJKUFNZGT[Sb5^TqSP[M@>6bVgSR^oj7BlG9S3_Y
0iXJ0TYB@_a8ZJ\NF_2c6ZoHDUmOn6PbomYlQ]C3SR7Mm?3d\g88m6N7XdG<<Nmb
@g>EBD_bB_84YED[dmYmnN4h1SS84>q68LRN2GYQ?bT_AdBl?F]CKK>>`ME<dkYe
5AWG0:WL0ai>h]A0Va>_b9jVBfLXAX26JjNnUmj`?YLPSPYnd<ALHOj64[J;eXJk
5=eVSfChm>46>8Ya^0CA6pSD5Y>e3RKAD@c^@K\7d6;2jT:U<B\17[F``9dPK4fO
I4Rh95R^WibLcRB0_EAO@iS3CU88fSmAXNOc2KZmO]3QpG\GTl6=T4I`4XWlCO_e
6o=V:S7^^567]=d;m:IL8S1<WnhMhO7ah^;B60YIk@mF5GOAhWDV_JNNLAAG_?3e
3P8USE23[dY0BDdAJd:fSc>gMR^1Z9=0ji0pP`AFUAjiC1TDnNC2lcQ?boeAQ<R4
hh1@4goP_KJVHlflP2eSa>]j9?4_XWk49e<ZPV9_B=JkaQ8f0TnQPE6haI:FEaO[
X[_15glEkY5<aKQQ:PEGb0GV^1pG5\=Fc4UD_l>gAf1Hl`Yh74X<[h[\I;h:?Chh
3fGDP8YP@fGUCRY_od1i<bZi4k7GI59akDfd_b]5L?<]Z1?LNFen3G=HK?PB?<GC
Jn3co\deWDEDT8@E9q\k<jh118Z0@KRhS>ShqD7QCOU0FLLJFml7a>DM0aohA46X
F;>fdF]C4XO9iFPK`C\DN3LHJaa9gIVS<XJZ?DRdjfNo6;LI:aVQF?3be^7qMC=m
D0HL3iBHbcB4B7OJ=D4j2=VEJYmLN8^5e5IMPdUXf=6L>;I\U?Ym1oTKCmJ7M?9J
8S13H`kR>nL]30]SSM2jM2;ToLfV38X]8X1RA`cAHD7n7BPJHiqN6\La^XQMRcR?
Qcn<ILSDR;AnEJ4m]P[kilEmPAUY57X0]:mcmCR0=IWY]=JkV?lNTBMPo]1nM_ND
3a9;_kLX73oXJ^?KZhJRi_5G`QXD4Ffi^dHCX6b?1qbC?<XcW<7Rnaa>iG;kDkAZ
J1d@m2m9lj2hZ@=31bI6O[`K`\7B]Kif_RlljYSfFobeKUn^?^LXjmTmmjHgQMTG
h^PE6ML?I5^h7AX>W;8SGL?V]B0bmMQRq66dZ]lLVT^da8nTo]n:=DNn=?AQcU6K
Y\1I8i7o^9cUiRdE>YZY<8egE^f3;7?<T6@;URKWkJSLBIV8N^]mCS3pSdQ4jZj^
Z8Q_:HBkI44\=e]9SZIG`4\<379:Y4eK>F6^mM2MAb3a>^j[RMC8VDcHSc;LM^<l
:]?kNbaYE<gRXEM:8:D6?WR5O775YRf2ef5Q0:bkc>No7=pYK45SU4@7>`0J8ihW
N;6C0=kQXKT3E0NH>b\[[AnBFJ:IU4OMEGlcFeP[Wg8ReWEYMe2dk0GL>EQh5dAe
jc8;Q;;JfUe[nCA`>=CjLD7g^;DlCogoB615KpC_DYmPHlJF42HkbaC]:?4aQH8a
l[JBHKU]XmT>S]G_;HHKHm]IjXhVEbT^PN9nUjCQ?ClKf8AF;bTDE7B]I9IFhFRm
^O1]<9W]6Y6?_;NRFn?3ZicaLNXapH@H[BLjY^_eK^N[=q=O27FC6;JCEN=0aV2V
T^hf\1Ld>^<X[c`A56LZfD3U9]c@^UNF_=M`V09fL=foH8=:<74oZI0C^G2Ifnn1
6aI]q^CX3\ipn@>@OSc$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI22HT(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
AGmABSQ:5DT^<_PlU`WANn?6j?gRAh0^E77qShi5LnROOVaXGHY<qBfDVAk:\2DM
hl[SWpldVS_6pdJ4XX2;0LZgYO8kR:8hSlXVXXVSAZKT06Vq;h<f5oO3YJSo9Z`9
5k4V9UE][G;HLHkgLmpf2jJNF@2E>c0IhBPZ`5KkD2fY:=[n>TbpbIh3j`WqnIEm
HS=MmR=6IHpDl;RfGpdEWUVeTeaO]^<;TjZdLia4i0OcE8UFN[@OfZ74UYe1H8ZA
d0Gc[3S]L7c2J4<IbIdng^cE^_3O8=N5[UEYNOS5@jlB6L876XaOCGa1N\IO^85E
JE>^hC3jqMC3A2N1X^Pb3C\IDd[P8Lh1GaI\DL6>foLTMnGn`UU7nfgmXB[79K5?
M?:n@fifMMmb70jAikP\FA3g?4^P5If1Fg_=>?<a<lLTL[4l@[b=[SFd_nGjYiCq
j?dTPog>9o0LKH3>Vk\\9R;C\`fe6JaPCV:[_Yf6b_bAQL]FoQU2[kL2G0f_Ziob
jVQJOH3^koGZMIX3aiY;NXZBTE;oe;k0kV<[@<bGDIFZRC`QV@>3[epbX_V25O\b
X;Ahfc^TM[N>V0qcDcIFO=KP;V4T1=5P1EV66kVoDLDMWdU^S1F:NDI^SCR^mWML
L;LjA>8ShDRc[e>cW6dN[IZI;X38[lCThJ]oKqmM=n2jIe?IWb6=MLoC:dXnOUJd
k`RQUG1^DKgRnZjCR8lPofPK344Wl_bAT?g38omgS>:2KGj301M1Le_c:LQmoQ4b
5=c7FAA^bKm9EdK4ZlDdlAIbBDZRpAMB]^Ui1nkDU]iUTVPXDY57XFo:?UmJXIaU
Z7DOR@51CUZ;FUdV:inWX=l71kjO9AUJ`<6@nRhVn_cDm3C5bNa`\[3D<gXPZHaI
:J>5QP>UdlJFXOo;@Glp<5D5FPR:@AjnNMM1n1DGd;56gadKV@]KIE0?_Q?=Yk[6
W6oo]\KF><Jaa1JWmgY8<1DMd=S45AfOf9Un2YlXMmXdb`:D;Zl3`E_=3d`MI^Mj
GI^ESmVgWopI5127c@QNbCC79h4Wj<C75oT_EeS\]3EYU?g^Nf26XfXO47I\0YUm
c[5Kf<j7?hGI<:kKK]kdbP]l0O7N=j@Yhq?U7;Y`UK2BZaoD6g;moC\?lKEnEi<D
147c37?=l2CW4cELRON;37m@\[NhgYV_:i?92J34EgQKUHOE719P]55oGYLecT6g
J\BcT>jEH;d]CbJBg58UF3RhpYDUcWDhUCHS49R;nl`2H>H<H9^88L81UoKDj?>H
GYW;Y[POZ:0PXlC^6\@M[E`3nY=MLkI[amLk;mANF01KTHYV6J3b[@PHHIKDj?A0
XO]3PKAUoGo8m^ep;R[h0fH;of[Hi`GlQ_RkS9iKPa?CSU]9RW4\8_McB6fGGB6M
`Gmd:G^IY<Bm8AZ>;3id?=`9KE>9Z]Q`WE8CSL2Shfm@N>=kiW_4TmQJMC;]N\c[
4bi_GKqf2hVIN`jShfFDb:Dfd6Y3=Gi:Rg89Jn3\;H4U0fk_=9TEjaY2co@E^nK8
c`HY8XIfVGkCN7k9Ah_VR6iUhcnG6qOnR;VOiLj>WcDF<X6`4lfVQ3=MRn[?PP8o
4]8g@q1<h>o6n@AX8<Ahd[XVH=DAhDIdUIHZcN7FF\^7gLfBU5AlL2@C87@P56S`
IOaoam1fd]fj825WbLVo5cJ;1DBK?bK4DMQ>ficFG6T^a^M6YGXF:f>7^K?0p[YA
541V=^3A;h41lb\]6779YV[hmMd[4emP<`HcAUP0:4?ee\k?I^N0nUabkU?@I[Be
U<CB<d3AVd5j5gbc;M[LkF5cUUgaMZmmdo`Q7ekoA9;oI]6_GaQq^DIIHBn9ldg_
@g<^HE]GMkmJiEJ6`S`jCO0\Zj_9eZ;gON=LmgMnN:TG`nRMln6<^4W\cjo[6d?6
1b=1YkWYnLh^boZGl@a]^OaEAPR]E2987cW6Z_@lCWqV5FiVk7Vg_Y5B;@cAl1=O
T:m\Q0L9PS1DkKdU<pd5RUnNbBDS9h=nabmEKhbY1;]B5_Oi10[F\R`OjfCG@k`I
Y`N7S>XO;cFJnL:TCUdU80K^o8mSQ1:`?YKgB>]SpfPOa:bpn6k1cDH$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module AOI22S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
RPMaiSQd5DT^<;MK@9n>h04G6T:YFg2Ic4Gl<f@EX\i??KM6p0E=1m=C3IA@;ceJ
R62@1ekQCJd=0qGmSYHQHD\;[I:EKIeQ1goXB\IRikp46m^\0qXAbVR\:2>9=a`l
6U?J<aQPbHoF3F8jbPlXqW0c=XiB8mAc0ma4fHZVfXIl0O5ZPKoXCZ?p:`1OVQ[B
XTF3ZU]D=^X\ISUF7CYoFQYL4BLRiGd35>d2Y8GQ1lB=[CBXqJ1iO2V<F>>e>\fH
DYNiO=I?McoToeC_?qV=o=SAaqQV9jASqU[8cjLEm4DeBm82EG9MbX4FJ]C>NWh>
`1M\::e]IA>S73=oEl35<:k=lL9b?`fE@UjEhV2llBD]Ja`J[5XW9`H8jb?<<Q0e
NgM=7N`6oJg:kKkUJDKmKV6qCmO:@I@H6H_7MM<eXoD81XO[Vkk;Rf9W;Wko\J@L
hZi]HS]Hn_AfR7F6h_FXf=ohCZg5Z6]F:HE1mkloMADlXTILG9^@1Sm^PWa8N^GH
mF@Y75T30T9i85q]:]_;PeTMEKF3g]I;_`K7J`HkQ@nUHfj2bI?PX1BH3YhMS\<o
M\GBmD4>I=3Yh3b][:jk_EghEZ8LV0MPDf[OjcDSBFE>hC27b@B??h?hOJ3BmW0T
C]E`2pBM9@:?2;j7?kUfMDo]N<M>XK<];<JKUKN7`9pmPHkM3nfPMHL<Ibe`RjUV
fEoO8TI37?7O[VcQGUBoif?fRSbUA895j;KAZP;J\9SmmY>^@MP7MJMUGa6=Z]lS
=qP2BKa:OMmc33QB;nD1TefU8`64\bOX4XM5VWW9W4CD[AQOn<U\hSEndD0BHeZE
O2P?mDS3CIjcb[DHH^Q^;>A]_D_O7^<3UE15E?HAEYWfIAP3CWV0>hZcp;bIhjL4
`VYJ3VWC39H5DGRMoC5W814W[X>5cRHkIAIeFSaDL9Hl@L^TjcX]e8NNE;I3N]L8
;4YEdPIH>S`VQI>cHT9:k@go5[>Hf]OTo55:Sbj5C]3nS1@qRR>S9Vl[V?4_;FLk
9jAh>3>[YO:cn5V\g6N081F:N4\U0^0e]0Edc@62kS[@J>T<RLNeLj@nF?e@meZ<
UYUm5EV_WO>PgNJHF6D0kYA_kZ=XmoZFg^[13OpG=JHPc`IT318T97iaj1^F6377
@Y?HlEMC@V;1M]S5i?NmBb;D5B:Ti;?eL0[`VNVG>U\Z=:_63Z8kL5l7EoQ8Cp_7
OBla8S3hX]@95UU6hV0XUcV3abb<Df`l02nREn<IZ5Y?S5g@Alai>R;I:TC7@S_X
Be6JQZnUA\DeP;;7j2W?Y8DL:[ncBAml]_aHZd@gA^gjQU\o4]Veq7K`dg_3Rj63
3:i3HW[E5G?>2Co;7=^o5GJ5DC[9_XHf1Z?kI3Ci=_F_3HVGmNh\m7Q2aT??khOJ
3BmW0m2`C<mM6EIn1<h[b]JGNF_bUhEZ8LV0M1<VnWBp^oTaA>GI9?n^>THN_J6E
SSE=SPW8kHmlFEX0VDlB^inaO;f5][>0=>9Od71O9faN^^_8ClA<23O86jdB\1?9
2_Y\DC?;gCj8=E<>BRYG8ENOXoEVc]L6QRqok5I:EOglJQIHF?ob?\;i6J_RmgAN
lFHTadNj6VhYJT97jYK[j6[CQ?_X5Qa]1VFooPLi[0AEf7F;6loZc[j03qXG1fh:
5]3WTh8D<RqalDdjmMeF0a]1;nR55Co]^nkf6Y2B4`aFk99N=Q_Z9`_E7dWmE;\Y
41PVj61]UT^a=KDek7MAKY1FQGN@1f_SCK2W;RGTKJhGkL0dLHn51h7jm2gF7jQ=
hp6lY?g<bD[:4^1FmKfC\AnG7AcL7BXHmYcEbmdB6<i[KGn3M88KU]_T37nB==AI
gZ6UCdCle=KUS74@nH7h]Li[:[HD5ia?BD=EkHT2E>[>]_\@jQnTLAF7qV2oBgbF
?3`ZIDk1@PAYB6I7f5`<Q15g8_T@>`1eUg^J?l[5c>X1dbcfI@FeDihWjVEDo1PX
0Q`hYREa:;1\153UA1Y^d:6eRMTE`6V=jJVERDOJHVZ[UVXqFUlE;fgB@4e?TU>A
0E@7Sj>fS8`IWmOjQQO7cV^ejgIG`6T@k2a71M1JQ904e6L2F=oeh^:K64nfNfdO
Z9EAnoqJ`h8RVe1g6N<GSdKK=^k3@GPZ3oPJDZ?c8coN8H]eIQ]:<A^>NPEcXqWg
cC^Tpm5o>_eG$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BHD1(H);
  inout H;

//Function Block
`protected
LA6NhSQd5DT^<SEh=VYYfMgVY3fgVfi8fR:n9KZC]?VcRGPXo22NfjoQGBWbKoqQ
Hk2b;_ji8anB9KOo]EY=IX<kdYmf]Do0hkn@nNVm3`YN=faCS[>mel>kL[2Y^ED4
<pj`J99@Doi9I1V5`;8bR69?7^ogBp77k>j`p9dL4lcM9W[61anHZW_cplCKAjEe
XKGXPbKET>K`A7=^P?AI6pnHmg92LqPSQgA9fQf:QLXTa?k1mVXI8O>RMoI84pPK
2022T$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF1(O, I);
   output O;
   input I;

//Function Block
`protected
7\jW_SQd5DT^<5YH4okLm0h\Y8CEF;@a<GD?an`QZTnYW0QjFd`b>5DR3=ARgXcR
aF2jV7=Wc]Wqjl_e1Y<3Zo=JIa<]IWY9>ENlG2pjXJ7`Bf5G^b=eojR76BD^hR@m
Se=GUZpe@XHUjpn=oKFIk?lXXki1iN5SBE]O@5qF`;f`\PpDmFA8Lq\XLh_ei1=Z
J5o02dk?lM4k;Bo:3NMCb`94PYRoLJl9lWlOC1G_>L2]dG5?<8_H:o\c\=XCo2Y6
GeDNee]^pFQ8FF?S$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF12CK(O, I);
   output O;
   input I;

//Function Block
`protected
R6cYhSQd5DT^<F<M5hEah7daB5gg5=qQ:@0\26XL]VJW62cnlf0?6Ve1g2cHVT@]
]P1nCcUVJ3T7Kbd758p0nl[VTUf^_8;6Lb2H_;kQZ;d5[V=PfWa;:IkqUffkEnqc
;lV5[V90D7OcMc??Ne>mB`7qE\;:MF<qh\P28LqVIoD8]<M?]_mUTjPIB59iZUa\
hIdB7529hVCco?R9jI2h1Wk9iYm?hQH3f\AEFjYVaKDE2S4bQHA][K`B^q0X:L26
o$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF1CK(O, I);
   output O;
   input I;

//Function Block
`protected
eEk9fSQH5DT^<4majTW;4@X>^0mFG`9Y]AJNIdP5H[JpHldQ\Sfj9b6^0n`N8T@=
68?Gb=p>@nUTa8TB`?X[1]mn@SF3L41j>2`aBMTW=;Kf94ib_BcF:ME^GpBoQ@?6
po:A<7Q7dL[gFE5[=TN]CJFgcpU1JAWFDpJF_FFLq>^iLS^>ooXg35VeB=aRNb<;
Q0^d[ea5\=<BIFWQ_\[OndS4h7e1nlndJQGcJ_o0j>WHWY?2KU<IUV8SadHqeJPm
`A3$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF1S(O, I);
   output O;
   input I;

//Function Block
`protected
VGmlLSQ:5DT^<3RD[1?lN?4?AH2Hf7]o^cff04KGldE<Q5m[We<f4SiZp6[4AP^1
NbE_0^=pXgHgh1[BFj2<@]eJ89n@a0EQF00`XB7>6VqiU7k60qlVj>RW4N48c7Ih
JVYSL_I@OTq>9Elgh;p:?kFg<cJDG2gjM45CGYp^\65Hmpd:8]OLTAk?:^Yaj@VB
d<gU:K^3ToFMCIMSj4X^j?T`afEbPCBW8<`f97[cN^c_Wmd0R>`GaQMh3ZXY^m:m
p`JSLg]7$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF2(O, I);
   output O;
   input I;

//Function Block
`protected
F4SIOSQV5DT^<5fYGXj>_VmHWgViUAOeH1?lVoG;g_6cCIML>5hPYP_EWlJG7<En
^a:I[Aq=TUc;BMoW0dA5F\FT:h1`nb=Hk[M?FX64SSRlBoikh_Y]DPpO58<B>OR<
TO:j5Kk7eG\i93cJAL5binAk[R[76DHS6QPWTAI<5^Ek[EmQ>hG3PU\Bg\XpWWgZ
B`qf9j\XE@^;`VVfVYK4B1K]]=JqXBAV0KHqOVbCcGpBfJC2mIWhX6ggP@hkM3O[
4h:YKnge^AA\:no3fCkA:G\ob_AbKIa8Z^FgaGbT>^JBA;F0NV[OeX1=g;g_0qGa
l_OSP$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF2CK(O, I);
   output O;
   input I;

//Function Block
`protected
P[khRSQ:5DT^<?7`L^OdY>SgqDFk2NO;4ABDhP74U6hc1_g4f\XR=a4W;lX1dSW6
c`YXp0?icJ1LKEXnh9c1EO_gFoHIffTZEM\Xq4Tk<nJqA:?mg=_e3;>kEa1R4g>e
Od2JpgGbKH0Xqne>iNcpbiH_bN?FdJY09f6?6D<fHme_Jd;;Z5TcVN2:a0iU69PL
T<Y0ThKTc7:I`ZkRX0lLbPVd0K^gmo91JWM_ALp8WIQk?[Y>[T\]bjK^:oCa6feX
W7Dqd\;GZ]\$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF3(O, I);
   output O;
   input I;

//Function Block
`protected
h7aUMSQd5DT^<ZT]4MFe>7`V5?4Q<Vj[3FQDGPpITi]>hgDcEGFGBKe_Q0B3YRMS
iOJ0Bd>>U7_fmYFVXBg`=ReOl@OR=7V\0ph7adoNiQ1N1;f:gB@8a_W>Rjb?SqHV
De?6q?b6AJ:6FmoOSW=Yjmb1GiHTDq=AHc6h<qekgl9LpP0KD=5HbFjR]eW3Z@:?
g9aY3dFVgbKUEl4WWJl6;X3T`_TlZFV`_[EG7Q\E0n;CeP@VcjFT`O8];G=kn_Gp
hiCDILS$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF3CK(O, I);
   output O;
   input I;

//Function Block
`protected
>@DZOSQd5DT^<2j1clOV\K>TRQFd1h9Q>kU9h@L:3]BZ>YV;^\6pRcMWH]U>A;oQ
VZ6Yj5AnMbe?T`<BZF@d88`q@GTT3Q8d19?e=B<H5U`RH19Ii`WK7]U]D7[KdfJF
9GPlC>>FC89g^X3pXco1ZmqjjT?7QQ8TV7B5ll4Mecdf0=Fp;?R4V@Zq?018n>pl
QZ:b2UYi4_A=;iSl_FB4J:YkDRFOM6d@WR1>23aa7TSWTZ6Sh:f;m;nHkD[0XAYl
7jn_FP@B8iXRm\:L1qG]4_Rmk$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF4(O, I);
   output O;
   input I;

//Function Block
`protected
Sh`[YSQ:5DT^<KSKe6N;kYORKm@O?SX9ocmc;Y87W`^Woi1BRoND_=V2RbMB7PWa
pQEgD[Z60:ZQh[D2knNSY2d1=Ja`16ATWfD9D6GXKq3?mS;dWmlIU7WP<Q>2382M
OPM\ZhOU81lJG`LQXl9bJUA=gHKFjRCJ0=WMG5IXqgRU]Lmq^B?_5XZb8I`8;0h_
3mjiQ>;bpFeH3fgYqZ0LfB`p>jAJG]UK0de4ChMH@29O]K80Ie6LK?`ZaOdfod]0
KKnlVj6n65[0LALn:P]6kSfD>DLefefjS4a4NCkaF1pS1N8c6<$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF4CK(O, I);
   output O;
   input I;

//Function Block
`protected
IGW\7SQ:5DT^<kobBn26GCeH2hRBA54I\8NeJFZNOO``Eo@ZPMfIcEJj67FlNR6C
[6_Z9jF8B;\kmiXq82Jn7cAEBDL0Bd3g73M^4QEa6Am?l0^9\j@dfPKR[Fl:8[=f
Imi_34qo@DBZH?>EbY2h>QED>1cYK<qY1VEgTqD]g_<=\GFWPmkSIDkVl@\1G@pn
cfe2Y`p^5U;:7q7=o[6B\KRN1[<kjMmD1<@7X1>I_jqYMK1[9SKF@6CUBk[:b9ki
K9JF4Gmo]J1?X4ja0gW8Fka7JYRiNePH>5[lKXRHJB7YZZnoh@]^4DA\\\_iTpR7
^lYX:$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF6(O, I);
   output O;
   input I;

//Function Block
`protected
NljFgSQd5DT^<P2iDld[[gPH>UlQR^=gp>98IGocfi?fS2;al<CG7f;BGQ@CA4CN
hkTGV2O[=R4aLeIkM9SDXg4_6GhKXO]3XHoTR9nm]pioIhQMoB1:mK2HIC681f0Y
422MPqom09iSqcgQKJ3mi7BNd?[JYMHo0;CHYpaKECRYhpX?bN[^loCVAb<Pi1UD
a1C;Xd1@nMnO6N6Wh95E=:dJ2FcFalJ[hlF\WoKA4q]eWV;1q7M4X^Ne<9MGL[MK
omfaCHf@:QIH>VW7nS?6@1Q2mC?;jbOiBdQfnA`Aj=fgJRD4[7n:OVAUSh0lh7hA
F;<p5Ef1`JY$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF6CK(O, I);
   output O;
   input I;

//Function Block
`protected
5cXN2SQd5DT^<PIlc9E1i_:Z\6F51\8P2M@;dC\ETSGl;Iq=h9c1;A3R;2^MkNHY
U^?nBB[YBE2UejpbG:Uo6h6fFdjFB^>[\ccXmVJOko0f:bp547AngpR;`VKciF3m
6H`Qhn<_Cn9ljJqY2l58b>q58gMKbqoi9>Qn6G9e[U3gVXCoPM00F<S2ol^\KiF0
6M;>J9h_HRBZH=i:fIh240B[Ogg27_oNEL5_Y8X74jFMG`5HqJHRCCLg$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF8(O, I);
   output O;
   input I;

//Function Block
`protected
X76`_SQH5DT^<0YY;RROkn:oSHSRm5KV;L<Vhd[9jDooD@R]>1f\CZJ9VI=p]jSj
@fl[L7E\P;RWPk_AVYe[S]OAdQ7Nq<S\OH=04MQM1ERAR`M79g^NmFdU5dY8WORG
YY]RY9DlM?ZMCK2ATIejeA`p\7U?h`q@ooZh[OM38APh\^ReUWdij:=q52AlUU4p
YfU<>7pflH32h]`ZLdVaOgZT@nFaYoWlO0g:3C?NFgJ80L<;Ogj`2`DK5e1if?mY
0JeBR;UfIfc7K_FIMII@aIjS?qa`^m@WV6mPL6g8NW<Gg@b6qoT7GYAR$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUF8CK(O, I);
   output O;
   input I;

//Function Block
`protected
nd8n]SQ:5DT^<7o1JVJ@]SbT\Fjh\0]>4InFc7\W]mcN:0bmIf@hKPYQBKm\@Zf9
I9hXmMnkp^e8;kd\ZL2\8@9SGHK_6goDiF=<C@Rj<3J`gJYm>>O6`dUUZR76DU>?
<9?qoCV4moSo_`eKDPOE;kl1EAWJ_8CQKY7e@W^223o1hSnAqcln=CHpZm7NjF\m
SZZ1hcJF=AQR4^=Op5^cf:^4p4Imaa1qC[2JPH`Q>jjNdaDIo6ZB0=3Cod1E0<je
:C2oH<^ZJPg`8d:5Y\F`bdeOH\beh`VZC]0JBk[S^mFW>b?\<=qL92[aAR$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUFB1(O, I, EB);
   output O;
   input I, EB;

//Function Block
`protected
:BnH^SQV5DT^<`YMPV3?glT:19aqTX3D[5HgI8[mGXldTIH85j1;E2R60cka\I[?
lhj0<mI5>3e5SMXRb2A<Cg0niVUAl@p`<X1QMICnB@H2ATXRl@V<1Y>gF><jHqO1
aGamqKIT1QPXYBjH?8E>SNk:nWCiji]HY8ePq_KgAX:8qKW0R^Hp8Bk`FNg2KOBN
\g=NX=4:95:4d7lSL8?W\U5Q`7:8;MfeFKij7J`6QbiOfQA3HU`d8_nNW1@\;:kK
Bib:f@q0HW0`g97[cN^AD60:V]63ec2@LOjJbdn0lX3i1bg[n^6P3E0EX\T5V4_M
hUZn=ae@B6kJnC>VbY?SmbVFfZLOCJ@2BJQmCSIC]6GHYD04lY7jlc^O5j3lR6T=
k0iRGFUJZZ8;k[^YY1\^4JMHZla2<cfjIOXcbXE5FOL17H]J504@dm`l;BaPn9n7
^JB`mjGIX72jll[qn]O4<lQl>2gPQb>LPCL;dD9g_DZjde@dfSk1;JoN@:E]f7jE
_EoUaQ:7?Bj03ISFKg:qm=QH8>4$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUFB2(O, I, EB);
   output O;
   input I, EB;

//Function Block
`protected
PC:H3SQV5DT^<HO18N8@1I4:63KEmn8=mOHnfj3eq4ZXB\bBGE5o\B_FSkF=lMCE
4iXeSP^Y^MQ8eUl41@bq3RAK[5gIkDQ^N0enB1]jXJO[5IZIf7VN5RqCc;Ti2pc_
O2Q4mI3KhjX?nOEa[n_9gPbJf?2TVphUk]FFjp06YHaB6j09;W0jZ8MMGnKf@fjh
fP5<Q4;WoZ5WX^BmRRDSX3=RONORRXL`N1qDC=XY?pXnbHLQ_4l393SoWGh[;mQd
]DDhAk<J1;CU@oUQ5k=5l=;k4ladD9Xa1KG]H74\=`XDj^7WBFiQFDbQM6mkq>GU
0leI2XVCe00cIWa3M7We0AJdTFd?d\o>PFc907i[YI7VAJMY2c:VgOc>4a5W1>^8
n5jOXbl38:cO;:9X]UOSYTYR[fKSMHSfi:;aAXJLmCUBkE^CRAMOX04XB59[8[hY
hdafncX6@XN8WGbaEOC?V6P:_[a6l2bM?mMUUUF=Q=`Nim`TOcG7PP37W7mI7T6L
fgC\1b607q5Zd6jl>$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUFB3(O, I, EB);
   output O;
   input I, EB;

//Function Block
`protected
mn9a2SQ:5DT^<4dbnB><:YN67ec1bj\AV7ZYA8mbKdK?<K8`o;V[L6q;45mAbn`f
h:SUZJYODp=mRP=6dSBV?IBF]dcI^<N4a3R@af8`lK;E4Hal\ApkKcPkRpfLFWmV
l^FH6g@I>MFI[@g6gT>KE;C=Dp5WDo4Ufq?7UXUjqE;RQYT=;K5]F5^SRGl2eIVJ
4mg92:d<QEiCA7oG<gfTSBY04AoQjGbH`>9ilWXU^Eih:h;mF:`dXQIH:R:qL`JN
el@;[]3WIC55=6RcOU?dEoPi<S71K7R=FU;2IH8PUOT`gO2^J>YeV_RCKk=[LC<a
mlFX2bRMdc5Y:PAN1em4EeXRHQ?>_EA@8R`YaMglJWi\2Qa;9ZUP>`;aZg>cG@`D
d0@PI<iHJMk:olFn0li4Cg>8g<=H9?M0gjiS`j5ieTeYbol9JHb^;JWEf_T0_:Xe
J[j<63>Gpa35L;D`$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUFT1(O, I, E);
   output O;
   input I, E;

//Function Block
`protected
_7b4YSQ:5DT^<[I`ESXG<b5hLgJ@=L`UbKcWI@<7j3O@YIL8]W;YhbRUjNOAJKWG
JGGqN`enZM`ceGmDK9nnMF==YLXlNdAfM33`=<6^fM9S2ONESa0Q2@l@O2Gh4LDZ
DEoEC<piB4ONIeGMQl\=len]^C3i6]QG7\d7EJSefhAEKhPZfmc06Vh[U:OqeLWm
mGp8c[]jNZ=HOjgMoc8\C7V@F\DB@U\KXp\?dI63Pq16]=ZQqP23\kZFUHICDhnH
V@GDkA5YY6P>o831@9E?;8=8j]a8Seek`4<3KLA?<W_gDS6_DPYD@3_6KRQ0]5i8
JnWp8UnAVEMDgFl@Dc>@VEO38Oi9Z2L2jMVEa3kKAYYI1>5mog<dGDcVN?UU4KPe
8W<gZaB]iD[0SNk@a?\GGNM7X_7@j1jYe]PiXU[GafND;N0FnK4IVD@:^NOHJBO<
k0a3inEE]J^fhZi_o54T4k39FIil_MLOEM:00;6:hOPEoE^7:435L?GDb2nc?GA]
WKbJ08JnOi=qnHjU7ni$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUFT2(O, I, E);
   output O;
   input I, E;

//Function Block
`protected
N>EYbSQV5DT^<h=`7m8VinqSV<YSSkN[l1^6oLd4AZ=kUo@cokcV\k_XbQj=OH>:
TA2LmfV5E7l0a=>_YDLChMUeTRqFo_A<?P1[Z92`TRYS9KVkPiL[T[a>\4kNL1Ac
=QI<g67>XCUHNCqS2VIXjpfn8>`RcQ2DGPo>L;oFo0D2k]4iQa91p>GO5B__qd_8
RkJ:@LE<QR88dZc;lY^1eYd;5]e6L@:K@L6i@O]Tk4m38S27[H[bq9lBhL0p9InT
T4AG8;HNATHEbZhaQ77TcGBTjPkaRXhCS[S`P7JLSa_J=YX>R?>?nLGH=LgZ98f9
D[d?@882`JL8?Bq@6Q?a99TOFoR9Ed^;:_QiJT11HjGGh3>miXeo@kQ;A3iU\aP:
Q`SZ[`i0ZBUPld=@T;9VI@]lP1nDV`=de8]coNCCPfII:KMdHXK5oe<dnYM62BiN
am2Qd^S06Pe:2:Peg?XZDOA=VM7jedVU`0lU>6?II3U:W:bcOD<C@>hAD9h_DWbU
W8JZNk]:n48gVKJ4AEDK0>3SE3qX2o[YH0$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUFT3(O, I, E);
   output O;
   input I, E;

//Function Block
`protected
Nimo0SQV5DT^<;EMKDK`:85_foggAh0^D7hpJ?n6U46\iO\]8=7_Ie_]<H;lD@ME
el3eD\Rk3]?dp0EK5a9od[TDBAhoJ_X:CD[T3MM`O229_TDicO@Hel^fI^Gq?P7B
O6qlQKN9Mj0L]SU:n@0N_5Unce::83I=Opb^3h_@KpE1?Mn>poE2JVQ8ZVN_a2=I
jnOGPEd6LB<iF]_6bNa?cg4MW75UUcVgm=W;mDL1SZK07OCOko781E\I=QlfR1e9
dI1qNRdobZW=>@\nIWZ4RGnalkh_a\\kFeh3^Qg^6A>een^5`gfkOPO^SjmoTH?f
\kj0NC;AkZ6IWTS=>5Z[fE[nU@DWab6OlGQIJG:W]?\aPk2WTS:[R6?@ffMg4XlC
JM4Y<e[fJ2hdAoT`<W1ZKPSS3[mXS=^2FKP<DhIf7E^Lk\@Q`IWmd]Z3:]6=CO6\
E3\`QS8J^C397M>_knYqLVdGlj7$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module BUFT4(O, I, E);
   output O;
   input I, E;

//Function Block
`protected
T:e>TSQV5DT^<`bYMi[YL28i6QX:X?hAc1jhI0?QX\i??c4IpG:JEaHLAYa:9WQ@
fF5o0imQ0>^AKkb`7PKk:\FoQJ1oIiAIU^[=TJf>F@;I?p94hP7]6U6FcC:74UVB
j=o1`iq\Ag9d6qEUK=QB1b4PG:D5bh6RDRo5EcN00lH1qX^?55C2qE4fcJ:q2B=\
jJ>>:SjcZP7GMX<2Cg;\_^M@`HdM]31<f1G[<XWck;T1=jAgS3Ti_n9W?6\j2`9Z
`A`:`O_55^Q[ClqXF:1gK@KiOXfEW`j_fJ8S`Zgca9ai:l?W3oTH?B[@?_Y@M^gS
3B1k0:K4l?T2W7?X=UhO62Og2j\NPTICAiFWVHmoH?VbF1bcYbg?<[imb<dcmeWW
X;>7Ah7^AfH>S\]>enTUL:b4bS^S8Z^@M55kL76m?n0XDd]T;FlHH=WE7T[?Kg0L
T5]]PhGHk>5cbG0C370Fl_b19R1l<4pn;:W7YVjV8402^P?PS\<m7YA]8Ylpda1@
_Z]$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module CMPE4(OEQ, A0, B0, A1, B1, A2, B2, A3, B3);
   input A0, B0, A1, B1, A2, B2, A3, B3;
   output OEQ;

//Function Block
`protected
1A_^]SQV5DT^<HZh`e=XANbjXWY5lD0KS@EbBKEAVR_mNGJ6[NnKhjo4GBVYKopg
BL9IFYb`ie]SZJSjTfqA\lk:l:_]S9HC2qKeAg\0pDX0aGB^[:ca_G14S]IQYXZl
h<b@SN81D`Xp6VKmVf4@ZXHJ@Kk7nKLkNVB;ZI_P_7bRE?p<W@eYiWeD\ME96m5e
BF_nY:0TjcgER7>\WqOoUYHT=7K2\IYSqXRYc77Qo45V[^;V?b`Ml_ZS4PiAMl4K
jI1p<Z@?P\TAcj?j_[RGO[T2\l11Da0X:D0>f:9KHPd2gdLbN^X`pnV<T6D`pg2E
PP1p4jRWl:H=LAiiGLHF\478KmQf@NUBY5nciki6]DVoaXW94mhjBF0c2XQfgHTI
X=VIihP@iHTUN;0AmjaT5nnN=lM46HY]5Jdb\oilD[7c8ZV<KG@lole<RcSdNRch
DI5P4728KFZJN^F:@;_E5=nN]lMIjjgW5Jdb\oild[7Z8ZV<K3@lole<6cSdNRch
Dg5<4728[FZ998CGlRcdp3L_0P[5PjkWm8=\;2GRUa_LaW8Rbh>Pd=Ji:[IJC?ei
k@E3cI2d;B0hRHSZoO7]@[B<FS6On]^gaLAl51>2UgiK<VkE130>hG=i0[CR;>dc
Ke>K\@bb3?nYTZYdc261R3Qh7B163]\1hdK;21A2BYiKSa^TE30>hG=i0OCRo>dc
KeoKL@bb30nYDZYdc2e1d3Qh7\16^I>bfE=Y?q;B5APn3QmX[0fLoY:YW:4_=kQ;
Ra;?12I9PmJ9\G`Kbcb[2N;>Y;6NBD[\ADcmJ:mEIh]V\`]DUMf<V15UiR:Lc1i_
A]?HR^koPkP0NSRKMA^`Sf?bFiVVTKR6boQ?iM;WkAUEjL]^1\g`^b5XiOQLc1:;
<3?ZR^koPk60NjRKMA^LSf?bFigVTIR6boQIiD;WkABEjVEJ^=hPicp;hF4bUM[Y
DBFbf6CNWXQmI;hmELW[Sk<YmHoJL7VQE4BLRf@;aVDD5B4B40:nYUeqMaOeH45D
?eG5?ZKgLVZQON7l`84\XRD<nR]UheLK31ST_cbR]^]ld1_C@Ghlm7oh7EINckS0
f?`SU5Oh2e`E7=5UTK:AofjeR[]I8c;j6VF_[KUV=akTVeiF_LHKP:?5Mo8>@0>h
fmMEU12X2g`S]=5f6U>noYj?R[]IOc;n6VF_[PU0=akT6eiF_LHKPN?5Mo8>A0>A
ccICoAncqhbUNR9c799AW=`i4^R3XC7XAPD@=CAbg^WK8=fl8\HJDYMY5S:SK:Yn
bPGGh8j4Z`lM3A?_kYl[7MQN10_A`h0egY9269>=im7KP12O8O60h:W8OR>>M8;U
hBMS\U;gBhMgY\mY<Y^_<LFRi0[A`M0e0]eCo9d=1m7KPM2O2O60h:W8OR>>MW;U
CBMS\U;gBhMgYjmY<oFEm3hgRq@ikR_k[CBdof=BdK`f<_ETK`:N`@EoYT4o;Ibm
5f?SAH5Ehl<5D`2W==c[A`ZkYj2Ud4hkn^]W6TL56`3FYElKafR4Pg>R3CLk;jY8
jJ@P[@=BGbc[nUOGbh^8S247OP@FeO>=f\]BhG5W;W3@YEWKaOA3`Z>R3CLk;j58
j?@P[@=BGbc[nU5Gbn^8S247OP@FeO_=f\gmY9E`NMp9de?;[V]FKE@amPhf\BKB
mj1@]IZk0>66=IM[51\[5VfE78Q:^H4a428XAiZf@Qf;8<RCmcGWHM=XhmHDBdaN
ICI\\VdV3ReXnI<OM5IaZe3fb27<mhPc]N6^]?_eIaU9ZT?Q;iMWgV6lCQaDEdb3
ICPT[45V3ReXnI<AM58aZe3fb27<mhPT]N[^]?_eIaU9ZT?=;iPa2SZ26=lp1@FJ
V>Yi0d5KC7;WnEkE;b\64dNn?2@@d6469LTMSQGn0X32KS7JnBKG^ASXh_ElmlNM
Aj;H@Ek`PJ:7kgWm`6K]QnYZf=:aJm4ffZFMYcOlC?``]YY7Eo@UJ_N:aiDh1JO6
d<@o@be8g0dCkJWmD6K5^YP3fN:lJm4fXZFnYcOlC?``]YY7ko@LJ_N:aiDh1JO6
O<@oW\4??b^Mq=WK7LK\gWm0KFj=0]hIn\cjFh1QTFOG3W]ob3E:K331jJQ4`m43
i2XR>8:lj8C\IN=bgi5Ml`S1TdW5bE2TcOhD3309OEY;en\oAVmBgYfD?All1KO_
kYU?BV9W6Ffm^=G3aV:k2`@cO22[]ElTcUhDhnHX9EV;en\oAemBJYfD?All1KO_
kGU?mV9W6Ffm^=G3aL:k2bH3EIM9Np5ZPVIha6QBVSlCfgZQ3fKjQXmSl0nm]oE9
e\C6bX^Wj?W<=oT0a3SYk\G1`<aR8?ekc>d\]Sl@^n[eA_NDF8Sek00J2`<83le:
eiSjlKPV54o7i^o62cYf62?ij\fj<]5@J`E[n[lL5ng]??N\FG7ekk6mGC<83le:
ei3jl6PV54o7i^o62cif6Z?ij\fj<]5@J`X[nCYFJoUa>^p7XbeOP5e4gH60B`7d
IXGM7MR1X=5d4PR8I<3AhAY?cJ0O]PZ;2WTd7O37O<J]PgnY2e]:TTN12[f<TCYP
^9CZGI@QR^BgUW9In<U;jbFEGWQ>\i>SUe;_>HD5\e^T[i^7lNmL`m_1`?j<JP`P
A9daGIa[G7lgUW9In<UdjbEEGWQ>\i>SUe;Z>HD5\e^T[i^7lNmn`mIKZmKc@3Np
djidjWSH`FH>_DfX5SRcH<R\:K`fgE38IlURTP:lpDdUCnTC;b5f:F8JIb_e`6:J
VgV5MF=9CZZ[kX9SeA72bbm^bfE@^kIf7QD:DERnI2Xf=RLci33:\X246^C_1WBB
M=d84k4aCFR[>Jl^CbD`6F:07YP_20FZ2Dig8g?ooD_2C693f3UIA@TK3^e_1>BB
[`YQPkdagFR[>Tl^mbD`6F:07YP_2GFZ5Dig8g?ooD_2C`93<TKJ5_BC;qQLm@gY
4kAfPHLl4O[BgQbWM60hB5gn_bH@X[Q;WE0ac2DYfhXiaRe_FXEAjH7GFdQZCBmm
E3;bAJfGhAGW8IdU`39n5]PG@IdOXWI7DQf[cEW6RN\j36_N7Z^FUVm@JNQ08IKI
[g;GBeTGeRG58c^U`3beZmPR@IdOXWZ7Dbf[cEW`R4\j368N7V^FUVmYJNQ08IGI
[S19f4?E^Kp^W9_Gh5G3MMb`DG6\MYF;`fV2KJO?fCAW@RfK1amJj`emJ6T3AB`_
:I`g\bOf8Vb6^L1Y5no?J_TGN3a^E1P]Sad[\BnaKNaK5R;ld_i]EOfeX<9?CX:2
7_6]l5F>b46^FaG74ne?EcRkRJF^91`bSaXGc;Ga`N7K5R;hd_R]EOfe9<Q?CX:b
7_6]l5F>a4B^FaGO4n1>Z:IaZ>npNl;d@I;K9?\ZH4B;TMIL\hW_PBS7Qh3FPL24
Q`D2n;[H4c[@RfGe7`lX=KMVif<57YI6nAJ>K`5IFCQWS<Ji9i9^f]\4FiYngo25
b=i<d`RdQTbl?6=G>fj2oPQ_GZhZN>3dCf\3K[AXcSL6S2J_ai9a7PZNFiYngo25
4=i7d`RdQjbc?6=GofjnoPQ_G6hjN>3dNf\G^WCgc_TSpgZTNTPfF;ee4Z8CmZbi
:ii[2]ROED=9VY[:X1m_AAd=GA4=qFdPZgBoMUS3WOc`l`623`hfjRXkkP8?WW[1
DlXONoGf]34a1`kY1dIFLhcTJnk0MZIj^C]:b1Wd<OIcSn:=FFlJ=0:\fcDEkdb1
DfP59miI0_OCO>j8ZXc?MIK_R4f7RFJC`=AfF1X:KN9Q\na=FZlJ`Bb8PcDEkdb1
DBP5JmiI0_QCO>j8ZJc?[IK_R487RFJC`mAfFDd\?jd8XpY]FD=MP7mIImQN38?9
5R\n[:^O8Xm^RCJA0AfTi7nWY:WSf9aI62;e9aXHN4NVOj:3bdmPfdoOUa2>KnlK
hj@KBP2PiVDdi_pDjRdKHIQAfTWAR1Z2jY`2@5jG5ehjG:3EnUCC?ffN`UlG2\2m
gDSle2aJK]do_C2jJS1LOIgWi2c8\@QOS]`NjU_\XDl_NE^?UU_hgRChNK`nffK`
[lmQ][Z:YT7=Z0AD2`2cN4jW\Nn^^M\OM]i<MUlSDh>_>E^?UU_;7R0hNK`n6fK`
[lmi][]:YT7=B0AD2`2WN4jJW[cGkSVp_9Ei2n:A`R4OPJBWK]8cFT\]mN0F7A?1
1eL@`g;_nUUkdb=l_RCBXZUh[LL;oH58JUk4YeKQAd10C4bV6Fc@`Qm@>AKJd>_Z
d6LND0^5Xnd^\K@DmoUWhDi_\D1bN8fI_?ii[JUZAYLn`d626Nc@RDm;jVM]di_1
d6LNB=^AXnd^\S@2moUWVDiD\D1bNVfR_?ii<JUZRJFM8JPKp86]>jE>i3J5G^bY
>23hONY`EaO[_EVEPjlXJMVLW3n::?P8B^jB1D]qbBFZcUNGkg99ERJQg_c9>965
n1i4RN0nZ:@>cV770SHl8I[dMAASWfSUdheQho_HJ=gbP`g17[_XeXihHLaKH:9T
K0CZXe]l:i@Z2\\;:QF=TOUgTa=`m>beMBR?6nMCb<14O;CM7;L[MLB?Heai3e9>
BPUlXe]l:i@ZhH\K:QF=TWUjTa=`E>bCMBR?6IMCb<14`;C61DZaT7inqnf8;VFM
ZBSl3gg?1I5ni[hdMmkEN7gi>MS`L1H:?:dYN2L@c5]:3g1@;O_;;n?FP@kVX`39
J5\;7Pe1[HF]W6GHKV\9n=K_TMB`A9:SO@Ia:aZaFlMQ@]]2]5KH3>VmFnH0_h=K
35JlcPcIWHa]GB_HV<[Nb=K_TMB`AeJSO@Ia:a4aFlMQ@[]2Z5KH3>DmFnH0_7=K
jILZI2VhJqkH1kjo27>0o[H;bff9?^kEXO8J32IKMD^1GJ_:aAR1M8ZiNTP[55hO
iMo<L3nhT@7SWa=^I]iZGi8=8U:XXl;Fd_3oTcV<W[iKGO_YBV;4hlBdV`2Qde:Z
Ph]IXNk\VSkGS^[;OgidJi<kl;:TXlf0dSUfYLV<W[iKGO`[Bd;4hlB@V>2QdeSZ
P`]IXNkJVckGS^?;Oga^96@^M9qdP\be<0N\3^f6:Pn3_DCDe9k4DfOlT>a889li
T`en4M0a48^4U;IAZ>TE;hfc=he4_EWcFjdlDiJXdN:Z^5Ll_1MAn]P2fRjgP9Q`
aQD1OJ[2;iice^K<BU572O78llSd`g9<c^4lY2QAndQZi5i4A1ImHMB2fRjgP9Q_
iQ51OJ[28iDce^KCBUf72O78Gl3d`g98c^MH8mnkn[RqVQZ2V3JaOn40G]MQ>^^1
k^983AbidHVm0BfnEE\0PX]a79^\c@m;123Rc@Rl>PFYG>EUB]k\o^AaB0_>a=fa
`U5IOVEih?o@ekfAFaJAAaDI[@On];JeHE:YiAlR9d8DVCgVQ:@:oeRV=4:ca:fH
[F5OJ2n`hQo5ekfARmJ5AaDI[COP];JegE:UiAlR9W8TVCgVH:@4BE?9mHlnp]K]
M]e`PX>cSfR94iI]k6\?MgN>47fcTQ6T3FG4kW?D@cIZl@@4<2HmTWQ8V?mFPl=E
RMH:b@bSB\QB?I8bRGJbG4_Ch4E45mGTBk5iU@dEHNho^0\^VoBU<RGeOb:8E]9d
L6O@@@mPCo`7UIKbR::bGlDT14N45mGTBcMij@dEHNXo@0\^VEBUVRGeOb38E]9d
LJO@BIlUnV1V6qIM4Xf[T05RfReLFUge0]2Icc]=R=8Ian>USEk`WC_mnSd9[=M9
o\P`K9PBeJCElmVjQ<6g]_cW6Zh:lQFQ[_SGSnC:?PKW<WJ3S_TBIn7UVW_E`^GV
1;n?aOMPLMEBb2I@j]=O`YcJ557boNF0[<nASDc\1CK0<WJ3S_=_In7UVW_E`^GV
1;2?a6MPLMEBb2I@j]?O`61dh>^0Beql596BJE`G9Uf9nPA[g=:T^E:OmI\50;]K
7e@SRD75XCA8X9?6Y]f39h2Uh3O06]d=\P\i@cfQSLloT;^97jLC?9PVB1:6>HoP
BelhUO^YMA2KWBVgIhK=JVU39P`WT^1l2AHi`HEQCHIhVW\9^j6jL9<[3[26>HoP
BelRNOaYMA2KWBVgIhKlJVQ39P`WT^1l2AHe`HOI;KXF_Z@qW2b>B6[NU[IN0_?_
_:A3ASeY`WU<J0g4LJqoO_eU7UePmV4WU2Taae4\VIQo]iOGPoH<O2d5af35l`:4
h7]M]jjMhYNlG9fZ597kf]C9YPK;Sl@8f5_<fhfWak4e`]VeOMe842cCIKc<Y04A
8@7\W]EY9_V[d?P\A0koKYhJ;6a;_:`?XM^<Khf4Yk;bfndeOMe842cJMKJ<Y04A
8@7\W]E99_Y[d?P\A0koKYhU;6a@kEOOD@mqf825dBD11m@6V9[_U<ASIS2S<Yn2
JElL2U?8X=iAOc`6_[jEFdTIc?3_b>0RHO_Ubi28=e48:?GZChR8[<<9@J^>Gkd2
9QKS:n?5N\mEk;SGSV^FS;kEMebXU<6Da?82foN<T>[l:]ZZ_Vg?[><f>M^?hfo4
9SKS:n?5CPmLk;SGSV^FS;kEGebhU<6Da?82foN<G>[O_A>9L5ONq`TGOUW^Qo=Q
AVh:93Lc[^4hL>D;C[e[Kenl=b?S4GP5g]6jK_mgWGGmgEghTW5]DC@Ho0;nQ@ZG
ZGIdj09bRN2i>gMMQ^:l=\1lX85Yj_FCMPJ_NX2oQnWCeU@@N[e?:`Ph[0Qjl@B6
ZH:;e0>beL2iYBkcM^@l=\1lXBdY`_FCMPJ_NX2oQPWCfU@@N[e?:`Ph[iQjl8jb
AKn1Fp`DGYHLXlClA9J0G48`ddDVPCE564[]:mFmWq<BWhg@fhIhEEWZIc@fWmZF
\DFS3eUk6e48TFV][ePJSjCJGh5feO5U\Zcg;0c[U=<I]]MiAIDehXK\W_c_KJ\9
9<eRoh6^FH6RT5\F8:6=Sb5J]>VAP0;6lYHk4hJ<E4<iXC<8oLD`U3=cSkc7KT8a
9YlZ186^FH6RT5fQ8F6=Sb5J]>VAP0S6liHk4hJ<E4<iXC[8oTeCCQnW1KqdRna1
eCGDYCa2RNnDE=<975hLRD55hn2hgm=IB6^LC;UUnFFa@P=?DIYhPeS=Z\7X]R7f
>3DNAZh;m>=?\_Sl:d`B5T0aj17DJm[T=E>4ji;eY:2Ff3MoP:im]Z=4RNHdXT5?
Mi<N86TaNNb?8_S6=d=H7\_aj17DJm[=ZEj4ji;eY:2Ff3MIP:1m]Z=4RNHdXT5T
Mi7=N460mQ1p:7cXj_<`10Me;lQ@Nne[RkaMdRdl@I4oe6YZKZ`P?l_=G5MTn@3>
[4kJGW=PGY5Q9FmHIbP3bUJQCh\gHa1E\0`T[Gg7`n6n\;YoFRc`_6E9fQ6^fcn[
4f:nYYiU1B@e:oBi7AIXbDFSjdQMH51fDB`79o\W`46n\;YoGNc<_6E9fQ6^fcn[
bf:2YYiU1B@e:oBi]AImo`C?KGX]pdT3lJ3_]3GX_Il?<SKM^[58iQeHDVO9^X^]
>o9b6VNLYWf_?o4N20;4V?GPDo<7M[CbHm^1Lc`IAV2A@CCJ^jdd;nogGJjanpf2
jJHH;aQPcKiV`:eQ6n8P_gY1K^BIP=2=FZ7J<1n1iafal>m6O25IS]mVOi6m;>RB
4mgY1gE262:haM`<Jmd53_V:R<@Qm0b6FDQGJ9kHa5PSD=\2IGkUB>Gg@2S:bXfd
QVNk@7E=BVaLe1`VJMD53_ofnC@Jm@b6FDYNJYkHa5PVDW\2IGkoB\Gg@2S:bXfd
QVAk@:<mfZ8GYWpcg^g?][4clFokVUP8`K3cZ4WjcngJQHY36?7m44XJXQLWmAd9
RodVTokSlE<0\cbR8mdL<JeXimNAG`e_l4_05c^=I<iURFna_?PFi[L:DTTPdGAl
O8Ko7j?a3Kjcb8Cc4RmgljKXi:9J]Vh_W4_o5c9nacBURFna_?PDX[J:DTTPaGZl
O8K]kj1a3Kjcb8Cc4Rm[lj`C9MDF@9cqO<eQ?6mm=@]SF@9l^Ci[6UGaT:mEj<E9
:b^^eH7H`l6o_\V;J>goOA?YYI9jk<HLd@Tc]Y]Gng@7<c?Mg?;4eXf[hT^V[TcE
fk^mWR6YlMjLPCoQIgS_>QT6807?Q7:NOa8k2o3Ln[GUPcaggG;d6XfFYASg[jcE
fk^mS@6[lMjLPMo:IgS_eJT0807?QN:NOa8kUo3Ef8`@8LPkq2fU29DoC<DDPmNF
LV]>dNMk0FebbhBVQ:L=T8CoImEI7m==HYI3EGXbS2M1kTeaTX_cK8]?l4aEC\mf
E_BInQC`bHQ7eHoR=l@=5iZ4f:20[V]4=1MmScUm9[4Ja\OV12>`IC:HQ4^7aT<G
=_EInNC`gG8NnHoR=l@=56o4b:20[VK4H1MmSD6mX[4Ja\aVE2>`IK:HVK1_meX3
2qRU2_P@LnU9C_V8cNMOjqNF_>;D[1J2h\DFl1mEHDA3h@3KcGa\\BFa3jR`dKIF
cbkXL]YY59IVmbc@h^O4_XL6HeKN4h?eM_g2ePDn9T25U:i8\<nGERJG3<O3;BTi
g21E4bFZenmZIZ_AB\]f?eN[kXLRBT?T0lfP5HD59;X5U9o54?nGERJG3<In;ZTi
g21\4XFZenVoIA_AB\]5??N[kX7RBX56[KPDRlqK_YVPn]he1ZLGajo57]^7fCbO
lWUS>nV\JJMk4R_MmY]m61a@[hjE78fNlX:3S7TY18TX:@ZYZEagna1m]K=Dd?Dj
4Lb;Ji^jGJ@@:gR78KKY765SN2=C>:`8VLcn^4;Kkl@cK6]YmUF>?MBmGK=^d?Y4
;Uj;hi^jGJ@;LgM78KKYJ65SN2=C;:=8VLcn:4;Kkl@2K6Pe1Q=`3`Up?Hb9AO7U
a\Zf`0PZC]:bD2mC74Gm60:HF70Ll4URMLZkGRP^[lB4P7bmGKG`aGnL<DDn\`R8
iknJkHTnFf`f>k;n@jK0lW[EYW0nPWH97o;;cZeE_SH?<>GTY2CQnK]2?4NKk@2c
i_`ABPlWF_`CDk;mPD]jlW[EYW0nIYHi7o;;c7eC_SH?FJG5Y2CQnK]2?4NK5@2h
Ob[Hm3>;qf6L6j`W=@eIO<JZ04?l9<G5^\n4]7[0cLGhGk1o[[J1MGmCK0M0Ih9l
LDc^jERGQ>Kc`Q^b0_JPLSPVdCH1Uj^I^7fJR@TlfL^h7;5@;@mK`YJ?k<P`]maO
\I@EKQk`Af<GLZD9a_mIeSIG7Cf1:<^I^U]l8@blfL^h7h6@;@mK`Y]?k<P`]>aO
TI@EKQk`Af<GLKD9cZ\D0>hD9pH\DViG`IX4DD8c1SWl1Y7S7kRG04Jg4^G0LQdU
nn=6nWhdMbl:]T9=06F;51YF;m5XKQIh[L<N\oa22SP`j@J>6n^[\Bm[cdAlL8T5
9[3MPLO[OOS`5:a52oN:\W`e<\HN6J5Xa4<<JnEElfP:jMX>6NX_nRmJckAlL8Jj
9_3MPLO[OOS`5:6?2QN:\W`Q<\HN6JCXah_][9=S`=pIOaY3EQe?2CJX12bOFFD5
e72`?la;R0@Y9I;L`l887RL<>Q:W9Re0<PF7^ee^\bi0UYU7>[?FHH9fm\cg_=GV
a9jm`mhP3:ookIFHa]:NMLk2?kNAoSo3m`I6A@HKN[HINcH@MWHFj6@5aaYg3=UE
a9X<QQgP3:ookIFmN]<NMLk2?kNAoSoLl`I6A@HKN[HINcHXMW_;V@_YYA6po`J8
@1C3ah<CCm9;Xg89]fn1c\nc>0kE>RNmJKe2\b:_9`M<Fa0d@7aObbMScR1C;2<G
<oo5fnImnHP@]@:Sc39f4mCNkNaH80Nd6hVjX52]GlQFDgfnmjRgIoN<:WP[o5S8
nY0cfaHmVf[G]C:MO39JTZ?JkNaH80Nd67VmX52]GlQFDgfnmKR?IoN<:TP4o5S8
7Y0ofHZl4SK5q_0fd[BZ>2^RoSoCb:hlP9V[I[9J>3Gdk=5@dl:j_8ej3Q<FlC6o
AbX1TbF2Q5@Cm32^H?27e?6_EfKFL1:Z0>Q2mI\jU4^RjZ[@\kBEV\\M^8IHHjBN
eY_oUfXUaQEB@_:blV_nh?g?faRH:1@Z09Q2IE:`64YRDZ[@\H<Ef\\M^8IHHjBN
e04oEfXUaQEB@_:bli_nh7;LlTU3>p]O@2\_JPl_8IO=<f5ASOO?H1E[T8`hphlh
[^nSS4?[\Y4H<Xl_THcC=]llaK4RWCCm8O=NdF4iZj6jP:jMRihZTk<nV<NGN;=N
iB;2?b`mZ>N3=ekPghn=8VfY^>HEZd=mTdcX0c[@;Co4YPZ\5TK9_>I5?AdF?hY@
]AWj4bGFf?WY0eNPFln=Bd7]2>ZEZd=mT[MX=c[@;Co4YPZ\5[398>I5?AdF?hY@
]cWj4o^2MgeTMqQ2S=K1blJNRR;@j^aheW8G6^?>\;YL5<beCQ2CA`E<5ADB:K;U
BIoUKB:Ijaei7NgdOe3b7G2P;Go2`8JW]J9LNIP<mQOCUS\JCklWhMBBdV[F9jbl
Z2YXK>X2BZK^0lQ1;`O2T^2QHZ:X\@JY]b8LNQP^B:OCUS\JCkd[hPBBdV[F9jbl
Z2?XK`X2BZKj0;Q1;`G2T\jgC;7>l5qED4JmY]7;AMRgiQE2JJ]J4[FUEQ6YYak1
:cgg1[Be;an=?cQUC7^n=<ZN@T@_]Ig0lY092dd@=PMkX;SK;>j9d^5Da;WnST3]
]c@Rdk8iO=RPhCPBEGZ@nH>36\fjmHOEW@CV9f?@=EZ3LaGK5>jJd^RiRC7nST3]
]c@=nkSiO=RPhCPBEGZI\H@36\fjmHOEW@CF9fXI6H5ARHSq?jjAcN@]9h7PM\R>
6oa5iXnTii@_6iR8Gk]\1fBGFkVahHSL\T=Cja`oH:7MgfEWl61S_P;iW[]SSQlJ
mT]PInMFdoW_JTOE_b][?ZENX`Z8D`;IjcPlLFoEhC;Eb@Ii?hPClJIDWjfi2`ZQ
mM][inMih[09JGO2_b][EUElX`Z8D`;IjcPlSeojhC;Eb=I9?hPCEJI1mWbkCbH=
p[HS^2nC`9RanM;]imAjDBkM]N:MnRd0M@j3F6fI:IJk`D7@XGR5c8m_MF1f_nI>
k:[cae@AK>@b;Y?YZ@:YXOib1h8\1FWU\q=7ccbMQ7KGb<in:dl0f8[NMm?X7L2j
^YjE=jUJhc:QBT8L2]9oN^L<jdF`KAInUA3gQ_>719ARnG6Z3NmDlmhg>_SS9Noj
ij50=_<i1Z1m5_Hfgo`kR>d9f<TLPj38hf=@?K5]@`Ao5g\Y<>m9lZeG>O]\2ZoV
ia50=_jf1m1m5_HVgm`kR>nkfATLPj38hf=@?KjD@E^2^RCg3EpH;o]X2UGJgARW
2oQY2D_3VaI<kg^^\nfk?:jfW<7UaQ3jem4=M\=aD]q^CbVEg6E2NU=D?n6h2kf9
IO<ga?I6T2UCdE:ZCFF>^4PDUioWOP0iC3hKY6YI]FnmQZ9\n:9<o_1GL_0[6hD7
@i=^lWN@0df6<EBX_5OI\OAEdm`KUW8bm3j09FhaiHQ^m6Q:?NW<ifbaj^J[Ph2B
4i=EbES@0df6<EB8S5NI\OAE]mWKUW88c3?09FhaiHQ^m6QKTNQVWma1eM`q37n8
hh7G^nnO_IQ?h033AFTUJf9@oH=:YMLG0dQ0`l]\IcgaUaJ^mU@e2iPLQ\c;;FT?
I]X9leg`TIoj:VhG]H1n=I<\MMiXc\L<HaEBk5E>EE3mTH;9LgbPN=HX?35T3[I2
lOB^l2BJK>>0:nhG^U1od5X_MMifc\L<@1Emk5E>E\3ATH;9EWbGN=HX?\5A3[I2
XhB9\\Co]k5[pF@Jl9kaE<L@Z8EH8QkB_EkIn2\NfhJbhX=8cH6UfZDhE@MW6N_^
??1JbDX[mChJ@4;M\n6:DE]YHX[VllL83^@P<QbPDVlJB_]8dW_T>d2X`Gnh=kPW
VY]RJUXmFEiZ5FZfl>_WdE4R^`JFJlS8hQmP_DjXiVlJB_]8dE2T3d2X`G^hkkPW
VhTRgUXmFEmZQFZfl:EWk;dogHcHFp?F98=3W6I3h`4mV@FMPcYeQoib_<7F0OaG
?lDJ6BoJ[RO;W1Le[i7B=_VeAoF4C=@G9cThS>BR^DjL9L==Un7KJ0F48JRNKkWB
?IUMChCZ;<R6G7SgKKdHmH?ZHVLUb9?<=;V>XcBIE4eRg\=OU0FLJg8@n`RNKkWB
?I05CDCZ;<RaG5SgKK]gmg?ZHVL4bW?<=;onXh>oRhab`5pcR[@U5Vd7:eih5AEK
Cd7DLB7XaUkU_2AE\=bjD0am:3K=BXQg8bI=R1iV_i;PYWk:XOF5^EEMh>EBMiKL
BZ=:aG2HMW=l3_VUF=V]`N61oH[;SJNi80U_8]:L16LB8A2c6dXFL5BMl8C<P9[L
gZciEGWdTm7li_[UF=VU3NT1oH[;=JNi80U1M]4L16LBYA;c6dX``5gEPO7]HhKp
Se47<V3;`4BNF6Q2l_J]A\fEmJY3_41`moMhDQ6Kp@>0;hh<I^EL7Nd9C[?ZJBaU
L0Mh7gdm:[K:V8bgoGb=iO?eEWf:]QH:HS8SSZKESehaF6hi]bB^ah2iFjd>;fLo
J<LX@jlbePB:FYQSJU`Oe:>eJF>4S0WMM^];4DLB2@Pc;hgT;bJH<@_BHjY>2G;o
>3GhNjlbePB:FPfSOU`Oe:meJF>4S6dMF^];4DLB2@Pc;jgT\?A6PH?hTqL^XYM;
[Uh\T@BP_gaI9GP\5mEmTc`hRP]Jh4<K4gD]b>nAIWC^CFVYJi<ZIHFXfclO]hl2
HLU>jj?EO\gd1YWh>FJRW[d<Q;5OhMg\X\GO\46<C`MlI4cW9WmFjniP1WLgN5H[
@=UMQfPo03g41=fN>>1>M8d\QJ5OhMURX3GO\463CTMlI4kk9PmFjniP1WLgN5Jd
@QiZlnYQKLpF>Xh5Hd3[HlX4j0SSOigO3ciQIi50TeI\_LT^T4^T9k=QAI[`_oe<
C5IV[QJ0QQNfWG:g^3GgO`G=Y9_<YQ@Ya7PFHd]o=dgNYL]m0mkAdSolS7k66@a^
:6\I1cn3E`WFV6@kW\bgZ=\9e?n<UQBNM7]o>IJoddgNYL]<Im3AdSolS7k66@a0
G6XI1cn3Q`WFV6@ho\;C4X3><AFpn^3lEMk1=K4>ScUEJ5M8G1U@<6?mf2@hVThl
kGgGAJCHh8JTafil[L8n:e0nfGeFhJZMoD;m27UEfg[L2>WBD`GTSbmBJ:A_R0hg
5^@SRm4]DEFj8NB>335PDO2d1>FDnooOI\9:2LI\@=Dg2RWB?4G`TT:`J:A_R0hg
lP@oRm4]DEFj8NB>UT5EDO2d1>FDnooOX`9b6K\Uk>LBpdRoQRnY;_0;hUgcfgCV
nB@o7GJ=MUYoV0afZ`=\2I;FePWf4\]YckkAfbfB]jkX3mh^D;kcjfZkLb]TlE;3
j3LG\E6fIJ;H>bWfVmKWZMjIW^GiPO\2aog]V=iDhJco_dA8h\JGaf^b>DTQ`Eh3
j5?G043S2J;H>bWfV3fW[MjIW^GiPO\2a;c]1=iDhJko<dA8hS@G<cH^Ph`eBq30
ahE7SF8F6AQP;7IecVpARPZ>cY3c;[HFj;hif`CLBVS1H\3Od8oaeSkgX=cK42H8
I0ZGGI>lZZ<99;Flj8fnLA^6]RVL@B?0`j7@H[dZT]PWVSFX3XO^3Sl_gWX@UeJ_
U3`]ch\67683[Y1;23TA]`BPTj^Le;4\2QB@K[@5k]Tc1nIX2XX^3SlGTWo@UeJ_
U3`]ch\X>6Y3[Y1;23TA]`B?Mjf7`PG7[UmpXM8Gg<Ya=_ec9Gi6\3^0I`Sa\V2l
@UhX6:FA=A1BJjkATZa1lo>jh=m920KGVeW23Je@bi[XlmTUmUjPDokDHQe?<=G>
0glem7Fh_>^3:NXV`;DKk7RGED?C`i=5oLgAXB0K>Ke]lUM[iHinD9kDm0eFQ\VU
0Sldm7FhnY^3:NXV`;DKk7RG`J?M`i=5oLgAXB0Kk8eF^6@gLM^_q706`X;=e7hl
K85D9bZ`S@Q^mE<LCOY7SmZ0MC2e5W\eD^oio6R=HGR0JOSMA6oRS>dle>\moSJQ
4lOHbc87@G87]^mfX08Q_h70>C3<ennP1Y]aAACCYHcmD4DP41?hB7GM59gedS:9
lKI7hc<7nZm7V6U0U08Q_h70>WX<SnnP1Y]aAACCY7Xm04DP41ZhB7GM5Y?e9kI?
^lEanq6nUhgT5enH144i9YGaH]^[FLOGBS1=`jRRob^i>A^OT^Zf;cj`]Lc4oeCc
]Tol<oJb>_i81_mfC5blZ8b]inDS;4m\eWh]:T]ioR=Xh<NCZWT\f[EO>gIT_k__
c1DE_@6CC?ch`2miAC[;:Wb;i2gJ;Fg>=Oh]:T]ioRcDh<NCZWT\f[EO>gFa_l__
c1DE_@6CC?f8`cBPkA9jb7pGH6@Bg2]ZG^IiJ3fVPU3CXj3^Mgaddn?f0@G[[Hh2
cHe9OYGo51QM>OPb0FMG;9nPNl>7[g=eIj?mIogGDG>^0\c4KoWna^Ine@^n^4f=
DZ4iF=K9o3_8P9l3:]>ZjXUGW1g?4lKeBaBaB_LGBG`@L\IGe><n<^7ne@^lo4H=
DZ4iF=K9o3_Z^9W3:]>ZIXTGW1g>Vl@d?K<DR6nqC0@^ajckd<=71b\LkBX]\J:H
GH;eIZNfMh6U?Q8a^^V4R156G;8RSF?aj@7XBVUXUEKT2jG7o?OV9XmACYFdT8^H
cf5PY=;Ip[m3Kh6;^O8DOKaQ`gU00iUVLXn8GTZGa:OR<Dl`BgFK`amUAM\K1kV8
E>^7KZfLnHY5gDK1H0gggknDDfD`mfRUDb:M0Ne]Q;jRU3AbBA]UBQ<i^OgaMk@[
fb<S6UZ1>[RMKMKEG083PeiaffV`OceUPWlQQNT]o;jRU36bNA]UBQTiYOgaMjA[
hb<S6UZ1>[RMKFbE7?HeBkZeBpFMf]A0<_G[ZSJSDV?OcYFnE9WVjXGSiM2;8RCf
VHS2a[UioB=[PI^l57^@ZmNB=N?]QO]dk_?_=M_5T=]U^<P[JK:3<FNGh[EZ8[nZ
aMT[X\LV5[S60__>VRU1Nd]AQlFKa22Lj;?HOKKQ<C][^aFTJc@J1`NhheEZ8[Xj
aJT[X\LV5[S60_JWVAU1Nd]AQlFKa2O6jQMa=ZN5Xjp7hRWHkJn9J9L[QHepN8kP
ED12g`RoTMmZ\I<STCJM<2CUA87flh\na<T1:\7o7;9FCH;TgWGD7S4T]?E`VZ7_
XDOi=M<9:4dLH;XS>V?T;XRjSmYQ6U\TQf70I8mg5X;a6?OD>1FW>lLbI6LhN3\_
Oh0i=ZEf<AaSHcXS]C?bofC6SmYQ6U\ThY7iI8mg5X;D6?ODCVF<>lLbI6LhN3\_
=d0TRb\2SRMmqm;dFdmhOE]TS7;i9AfF`nJfK8]^U6V?>8PP39c7oA>61^>XFeHk
CHW4cnN=:0?Rga=jL_`c5hIS3n6KK@dOhDkF?DedQUf\`KSPEQZJkB\8=7LG]f>e
JHRm5ef_TRfJ]m5a<0WfYh\k=`F6;@LOhn1FgRPbGUf\`KSPEZ_JNB\8=7\G>f>e
Jlimbef_TRQJ:m5a<<Lf=4XQ0O0jXqn1k846SP^a4IAoH@BgFg4KTGWZD2J^T8=j
I;l[<Wk<Y[8f6CI6g]Iona9gECX43LG=J\`k\4MW[LHMc5Vo8jH2K2NHI1`ad\R8
ISKn`=cIJ2@:m6?Z`Jj=7OP;0Xf[eHnUS[iUDOMKSSciFkVa8>5DKk3T31`ad\R8
IS2_`XcIJ2@gm6?Z`JYf7^P;0XfceHnUS[8IDjbmB5:hJ1pFSF6ZDYWfX_b3M>JS
L9Jdg\dcVEK_CR?nYWYLUe:BIlQZ@0FTR2a@D_a2<JaEBHalhc2ISAO79@^h]?DV
>Y9l7K6AQ@=7OB<@EWVZ^9ZU96D:am0MU[5__WC3MKUMgh2FDkG^OJ`7U0l6OfiV
hY9dRKh798=7OB<@EWVXi9YU96D:UmiMU[51<Wj3MKUMgh2FDkG7YJ6DGTVmKQ0p
Rl]Dg1QRcI^UP=6b9JFcN4an?8>M@J?CF`NUlTV2<]6R0HhRWQKKFQ9q3n`FQHTa
0h:fVXVR8DOVG7OKK8<lLZ]CNMEdZC`5KP_788<D7@GLLIfO5aS_Y>lan2=4]Y_Q
`@TK>[OoQ@_K=[2l7l2dGbiLU6E]j;R3an8LXZTGS^U>Xa2PMmI^738c3_>8F9cR
`4a]QJHAQB_kK<2?RjHIGViWU6E]^KR>an8LXZTGS^U>db2MMmI^738c3_>8kncF
?8WIm05gqI8`30b53><\1LAnQEZB561VRd[EDDQ`@TC;MFJeQOOF_B[e7g?CmoP2
g=4f>5WhgIoKaZP8gL:hkOg^1S`A9cghjDCPBhN8g2g;0SkaM_VFRmN4HMk=_9l>
\BCP7Ji^LI6R9BV75LhaL:`D4S1A56mh=C4Deh78a2g;0RLaB_VFRm64`Mk=__V>
GBCP7Ji^LI6R9417FW\id?o]cp8@SSOSj=nRQK<O[bj^MBXgmD?H9K9l_K>5cP8G
MJV9C37O4N]7g5E27ifZ4^7_mYbN@6YRl2X?L[UnJY8jg:dUKZn9cG^DnHWGcG7]
`Xm201:YMNfUXi<aDiR>JYH^aG8EF^9VnAXNn3H33h8Ng:43KSXmX2^DnHWGcGJh
`Nm201:YMNfUXiD?DER>JYHUa88EF^4Bn]9nMe6W=2pU\b_iUH38LfQVE>@QheOi
5[aogNi85\bfDY\LXH[G38lhJMKbU3:lTh@<>1Jj?b;YiG<M1W?hKE8YiLCKmGO`
b4APc:Ce=Qie\YV3:oOhN>VIVWQ>fc5;O@1GBaP7BJ[UBSnYinXhRjLJo5HKMG;`
<4_I?IAeYQie\YVd[oMhN>VIVWQ>fc5=Z@XGBaP7?JSUBSne\nXiD5>M_GCq\H>F
;DZ7?IKS9I73[0J2^Ni0Y\9FkP7IH_b4YA1O]Ja`EIJ:=m<1dJY51^eoCcQUK8b=
V<\`AJNJ9JdT;WPSgmOTX@]0`@C=>1bY0j_F2J2=PToAVE`o3:WbA;GMJ=;7\nnF
fSRNA[I@c:Fb;BPd^hOOU\ZI`AC=>1bY4j_X2J2=PCoAVE`o=AWmA;GMJL;X\nnF
B4R^MG>0P67ZpTI2A6RgT7o6e12?EKF41cIj>od3ILn9BUea:96<X_BIDN5S<7L4
DRM3WYUHom6oJ6@XY:K73nS5<_bdC`;92IbFG8gHkaZGAY^aLf?EXco_=j;7[ngc
hW1l::Gce\VL<TjNC5]S<nAFC\OXH`e92dBFh5I6eaZGAY^aL^FE?co_=j;7[ngc
hnelI:Gce\VL<TjNCFUSiX<fhXJISpkTFog9NNfAO1=a7m3oXRH3j2Y]C;dRAHkQ
fPW>U:;5=KRA=KbEUZc17\ND`jh1:YFoDj]:eEp6;?iOCihN[cjiDQR3bjFG0<^g
KcdfK`R`W^TQSFQK6i:7MKT=obQ:;i>0dekSE`i@iK2X_@4@Ki4DW[PcW6_GFmcg
;Rh1o[d;W^<T<?T>YC^_W`QMNWn;74XJd8AE=M@66;N?@il@neolZM3cc6_Glm1O
U`21o[d;W^<De?l>YC^_W`QMNWn`l41Jd8AE=M@66;N=<iQc@^3<4:^qXAg?fZ_;
>8QGlk3DQX:7VTFXE>;lj^NG5NMHSf?aONm;a:?FcZ=:elbMWaKkQCbZF5_XKo3_
:SDnU44>ON>9oiABI@[gDlUOZ7M:^QQ6ZBXcbjjn:bEaC^1;6FXc8E1QX]d?BL21
:dY3JIQ\O0>9Q3Ad]QdSD7UOZ7M:FQQVZBXcbBjA:bEa4A1B6FXc8=1QX]d?WK2h
a0BdADk5p9G@HOI[6C?WZ]A53VmhlLT@KN@HFP=7aM;e9c1V2m@;>iX<U=gDJUnY
8iiJ0Fk3H?1X2DQ7:jG^MdCb7PJQKD_RiQHh>gSBkiHeC=O[Z:eSmd5Fg9YY@4A?
]19=F<ILB9]_VCfE2j0fjKmd9PFQkLXR6UhUcgQBIiHeCf\[W:eSmd5Fg9YY@b5?
;19=F<@LB9]_Vc;EW91C[OTQ1qR?d9UQZ33fOLSdc_[=31]\2Q>NC6@>HC=W_;QJ
7Dad28IQoI>];?`o@1hUULnU=`;WEfg?ZNK:fi<EJZBK8Y^V4hV3BJhYIGeH_`GV
3^mTaFdf=Oh;kQ5WKa@FO^AJK^RgbBDFfSKoPEHdc`Bi8=]<4QfEeahYIGeH_`Oo
3=mTaFdf=Oh;kQ9KKT@FO^ADK5RgbB@=fA@<[NZkYFqUBXmBb4?`35HYnkGC60N<
:7RNOf<59L?=hlCBge`l40Ad0k7mj>8ka8Z;PSV?kTjldj:g\e`i^n>_Zn46J9Bn
;dA8mI]gG4^qi=US@igJ:4XgI5liOFmWbfL\:YA=fV^@@JJ4bW\mLPCeX^=jNF1a
=0Y7Ee:MKlKpcLH2LRKi]LO4LONDV12>DR8OGle4ODbBD@6oaA7kG3^Uj?a=L]W0
@WBaI8e:`_0LLBNZBJ420@GLgUc3X1_D72mkK<PTV8;EF<6m08Z]nCjP[`Jag9dR
J:RPX:Xf[J@Dc;m=D?Kh0O\c=RQ@XQ_i42mXJ=AFV8;EF<6mb8Z]nCjP[OJ0g9dR
6_RUX:Xf[V@Dc;m=GRKT[;=aQeeJqj6kFW]YVf=?RJW<JT3Jch?@J?8bAUghna;C
[MhT7R[0<=K10[[;DZ[aIgn^CEXgC?;JKAXEg=CC3ZnbOUS>QBQ`9JY7=[Q[AoeC
X=]>P>F?6C3@>i_GkhS9;5\mSFT>7jZ>`C5gD=a0<19LcUS>L3Q`9A]PY[Q[AoeC
XK]>m>F?6C9@>i_Gkm79`5\mSFT>7jZ>`?eg<o4H=39c[pUg`Fa=UL^2fFT7<ToH
aJlN2:99S>CU;:O@ahC14MI:^64dKSQcahGY88c?PObYBV3K^2SnOOjdUERn=D63
@gc41b3>BmC0?BdOahhGTY^@T::Xe_KZ_1bIRog]606hC5U:X?Kl?Dj<cB[A4m6X
@gA41be2HnCf?NdOah?GTY^@T::Xe_KZ_1W7RYg]606hC5U:X?8f?mM_anM<Q5q_
E][Vj8QDAdfC@\5ZdmcQ]=V=8\fEgU`7YMp4oXj`Pc`m;_bDX67glWn;W<SDTjkG
SYEbG?m1f<@CHd1RbaXmY\c<MXcJMVPfS0Od2YTHj]U3V`F2g;VNFLIZc0RkoDF4
2]]`S?7gj>Ueil0=VG1\:FQ;bZl6c3N[Xd:4SJoKAoE3@P\AB9oN;LKGc0CA<ll4
i]d`S?78j>Reil0=XG]\:FQ\6Z@6c3N[Xd:4SJo=SoGLeNBmgTlpZ0=WX58aSPeP
90>ZGEgGU\ZYeF:kKCjVfb7IMJ\k:iJ3EZU?0@NL73DL6^88]GiSi:c[@IL48NVP
VA^NcI^<0RYkl:53SbmZPR7HGR7<^<V9G7R[0DRf9f:jlNXLP:LRZFFT\`\h8:nQ
@Q?Rcf^<oRYcKgoTSbmZPR7H=R7H^<V9G7R[0DRf?b:XlNXLP6LmZFFTbl\`n\2K
lBEhpFSSQQk>kS^_VV>Qc<<AncjHTk7AdCRH;NO;hlcK@eN><4jJmhdK5K35f<>=
>6ohGSVR=5cN23bnini25JW<ZSV:<=eWG6;QPL0;7mLSflHg18DK<?Qk>Wm6WlcJ
McJ9JF5BolDYc3=N7Wi]bJ^<P^V:CPR9462QPL0;7iLSelHg18DK<?Qk>j66WlcJ
Mc=9VF5Bo]2YeKFQ3a955p3\LED15;UKSD]WM`KULJI9;jfLQ1bL43W@PgEBPHl6
D5UWl0YE`CDVkR1Emf]Uf`CWK=C7:eTNh3^M8m[N^2UGUU;jBAji]3O5P[SDkHj8
O7@4R=dQOb65A:4?`MPMeX3aaFEb>CT0g4YjUS[9^2jGUUk9Y<jj]3O5P[lDk:j8
O7@SRVdQObm@A`4?`MP7e43aaFDW>>iA[V`:m?qP2af:3BYgK4L8>A=;KmcO>TiU
PRN>g]>91Y4Hf7<2=3WWX0:4M4JW]=IEGlk[Wd`LD4LFTVI]nk4Y;WMmQS5UM\oA
KP9BFR]\nY`Uj915oD:];8E@Q?dSkHlFk=gHibjPVDjmGI7]@;RA@`QmUS5dM\o@
FXIBFR]\nY`Zj9<5oD:];8E@Q?dQ`HEFk=gHibjPVDjDIIT]1M@`jGdqE4b=7]Ri
HYiDiG8J9Kn57AD1[MRZZ6LjOAXKkofVd8lDW4@>_TTYdcJE3Of[Zg[3B1:?k3Q<
<28FEhj37Rdm<2nT@[b1Do8fK\X<g\DKL@SDgX\VelWWMJ0I5gYUlkb@E=lWD[i9
<McXX]cZ7ld7_2nM;LCDDo8fK\X<^\DHL@SDgX\VelWW6=025gYUlkb@E=lWl<iB
f20mQjZEq_Y]22B3EF=EAA@cCCbJK?YHV6WUIL0geMRnmeM67RkIaKFchE1MEROR
LB[4P6SdAQfD]Z2Z_>CI<`c3;;A>DQN>mnca?Dc1]g]n83Y3j@N7>jQJDgoATeEQ
_hma5objQ_DjW>3kk>4@cXaeU;X>DDN>5KVB;DI1Qg]n8RY3?@N7>jUJIgoATE;Q
Uhma5o2ji_DjWH6kbRLI0SV?XqANoai0O0Z;;alCqKDEbmH27`^3:?bTUN@3QQM[
dQMTo\KT=[Ddm6P2AQ2c\E7\m8QgHHNYmB4>eQ]863fL?n\T>L5FEPb<XTTE=Ecm
AJ>c<B2]Ao?dGA9M0PPZ[H>L>2<ELo>^igQV3daKDK0ATU6o]LBZb37V0TeE=Ucm
22;HOB2]9o?dGQ9M0PPZ[H>L>2<EL7c^TgQV3dNK:K0ATdZo>=lO?>gPSpAY0lWg
[@;CRJlKZb9lY^XVZbJm?9FMUM?LJOZH8]_KP3WcL;>6@C4cU7omLNg>oBS1lQb=
ZcFV\^BbBP=[7J^2V9b4WnE^GA>?JSm\nh[1K5BoJNMM<`W@j=26h]@n[UAeABc7
U[FR9J5MHa=97Ji2VG4<WGE^GA>?JS;\ne[1K5BoJNMM<`LJj126h]@a[UAeABY@
UhQT_c<K41q\ZefF[`fIgSLg5FS2W95MZ\NB>EcIa\PiXgfKCiY[NXfLfMW8eRKk
<g<aY_BHg?LXm@cF`<9M9Y2FP<5j=fQe<_jn=i>M=OT55g`9UBZAR=B?F_O8;m;D
@>[cCm]0[MQ\ZZl^\UWM0dVkUoNjXfnj<_?NYAmM8O\55g`lUBZAR=B?U_D8;m;c
P>IcCm]0[MQ\ZZljRUW[_kRUUQXpD>8T>daE[iCAP`BmWYpQZ4kf9cb7_NWnLbG2
@IY7c@d@;FD<2Gc]VUfFB2A@iAf:W0nJ]FieUM0`>oBfeHoePgV>:8D5Ec]G[9=V
Sh1FBVCH3C6><96CXUffk?DDi7OWdK<\C;ZkCO11e4n[hSHQj>Mf@7N5^HIgaCmV
Zh_EBVBY`36>`9=CXUf;k?DDi7OWdK<\C;Zg_Od1e4n[hSHQj>M>87bYlhFm6``q
E5\R<j0IUoV`b>[9FEYQK5KgbjI0T;ekd1^Mh^XKIF>?;fGFRT=aUn0SP\ahXHfa
>IoOkPi2AfhI=j_WE6Omnl;AC\1L`67Nn<^fe6O\H^D\cRgm0n>\Ci7Y5l1m?AVQ
E]nMUfDRAHGRNo9AEoOULl;`?A7[`67Nn<^fY6O:H^D\cJgU0n>\R\7J5l1m?AVQ
E]nMY4D=`SO1fFZjq>c4LHJ2AdhcVm72XOWdRTDKQPjcR4FSQUkk8gj<dGKYgPY@
jVj`CGOA[kS2oaRB^KD>BAe:cUl=GFob2>3UA2KNom2XD>HP7[akbKBW`<jCjjff
\mkKgj3D=cCLf]]LU>?WM?=QRU<gQC5nH>2UGDKNS4Ukd>HP7[akb3BW`<jCjj:f
SmkKgT?D=cCLf]WL]>?WM2CQG2DYaR=4mpAEhNl]1L4o<eU=>f;6R\KeAAd70RVG
GCKDiS;8B_ak5FKHQW94]WTJomAIBRG:0I?=:e`SX^Cn4OPTJMK9=19M5@:gDkL?
0epV@ecJLl?M^@LBbDK45B5TJe;BL9M@8IL^Z0W5bO^OLY@IhS1aWIKM=Dnd0XmP
FM^kIfjen>Xmjgi21ePWl5XEA2Y^cbKW0MGiR0k[k^V@knTQh\`lhEk]gM`P1l=C
FaQVQ7EaY^CmSilc<WDWF5\TR2C>J:3W0MGiR0klk^V@knTQh\`lhEkOgMBP1l=C
KajVQ7EnX^4CGN@LKH\qNe@>D>g2m[W_K@cEnXP\V5H_;:8IkEa6lU?oeo5IYDEI
`NVJ>BGTC]D[YDB:iaXQ<L_a=VdU>?aC:P_RK8_Dn;gTFQ[HUZn<g5?>X5gH2ji=
@U=`>5F7lJ^o?PPlE`:aN?YiCAM[>=7Z>;BPKW_5`Lg[=dYPUZn<g5?>T5gQ2ji=
@U=`>5F70J^T?PPlE`:aN?YiU5M1bM79dY1=pUT`cbZH_P<P=HbLhK75_mfX4SjS
VM9:VKW;\=_?oODdk:8TqOl>J@QVl5nYTV4FS`kZFl>f7G;XVa;?PfGQNbX6cVWC
m5N?j[1mIfQWI6iP04:@08Ul\Ila;3U8nHXI@i`]L0eM4=J=HMfaPjUQ=8?3l_N>
Z:eDlcfEShe@g:0PBMjE:OQb8[J6M3B?Ia@8LiJ]El1M7gSH8M1abjUQ=R?3l_N>
Z:lDlcfESMe@g:0PBMjE:OQb8cl606c>92l2<pPA6m9Q^QH7:3^h>[D:K5dGPLFh
m4ILI\FF_L8;C\G2Hn]V9lengF9UP<Y;<LhU3lV<YY8;=:2Rf_U?X;WPiedfVmdH
IOBJ4mZn_4C6<`9K<3n\^`X^F3@>OK`<0AJ4N[PZbfQZOV26IkB7nfWCiXd>VPmX
EVBF4mZn_476<>9K<3n:^iX^F3i>OK`<0AJ4N[PZbfYnOAQ=F9Q=Viq\HVKA4UFO
Kai4<hm@98E3>VSAa1Y`lo?\CDXc9ZeG?LgGh3Q@TJ_]8Tk6eZg7nAmh4\HWeb_6
NFNfke2n]j6nKOFT53_\MNLiEDY2oR8OjneWRin_Y[;bW47RFP>G^Q[\n1n_Ul:6
?L<_4\nnWjBE@OjR<A3\MNLiEDY?oRaOjneWRin_Y[;5W47RFP>G4QY\n1nG8lK?
=TCbC5jpjMUNCPhDYSC6UdK9:l4JoQWMh\9TBb_5E?hA[ZbK8goQT_WZaFf8Llc`
P\fFmZ0]LcK^HAKWWF\c1naWa4<f\_Di6j@]KG=A>`hRmPR5`G_]h;@@Jn2NTdgL
Z]lfUZamj=b5\UdbWS6_hcD5aV<ToTDLU7^6KI=B>`hR`PR5`G_]hR@VJn2N2dgL
Z]lfUea9j=b53Nd9[7UUmlgHpd5A\1hUmOQkI<1[JNnYfN19>PH961k<4BZ??NZ>
YIOkd<U8EfHTIZ6<PQhI=YoXoXj8`BTh7leZgfM_A0Vl`g?^XfkRHbLOZLJ?\gj_
7j7d2ED=E`X;b>FePai7fBodmd?DW:^]Ilh=B3g9O0hl`ND^YgAc9bZO@LJ?\`j_
_j7d2E[=[`X;bEFe^ai7fB4d`d?DWl:]M4BN00CeYp\18fMlfm^7>lJNJFha70;R
eI>knQE\oE\88]i?AUU5>nP3]N<7Jj9c`VJ<om45;b@bn^Z0AAf:RSeJM=C3;7OT
]dJTKRSAe3oH8^=UBieA;UBc?Q^[2>9PND>]M5g;o[\d6\mBJcfe<ZW3ITC1;7G=
]bO4CESAe3oH8^EUBUeA;UBc?Q^[2>VPNF>]M5g;o[\d6\FLJ@UJCNL_4CqcL[fE
>fABjNS7>[Dd5`QkTXA<PjN>ZL^[dB2;<Bi`DFFMi3HFP4h3UUQcSGb?m:FGUWgV
;oL@UYjD?T?P1Hc72aIS`Zi;\NL^HBhb@^]VHoVA^e@DXo1j0m_e2;Qhn1ack0oH
C]3@?G^0R_FPZH\k0ad6UYd;\NL^HBhP@^bVHoVA^e@DXo1F0m]e2;Qhn1ack0o^
<]a7E@6g?l\q7nJVT<=3YC?a35^G_51QNoM7hk^QNn`^fCULolePRV2\[]d<h47A
3ie?8j8\6JAaTR3b[XBVS<`?0hb4L6?U2KnQ`DTSS@\GlDUIn6E=?OS3Po1kY2m5
m^J_:4^c0d\j7a>EQZ<?SU=?Ym^mLM?2FTn9mM1hSR\RlDUI<6EJ?OS3PQ1^Y2m5
;^J_:4^c0j\F7a>Eh[<:nL1G\R<bqoe\4fMW=:`h;OXFnnRoWFl]Ug?S8Wn=RhdI
8MRghZi^ceX]_H]9Fdm]<L@JebU>ok@4iIH=;9_=g5cO<3@40@>ijBdkjgi1V<6I
Nej1C?h<B>PHl^0[6MO1Jk[_`S`Y7oaOgIL?e9WHg:;hF3G4>]>i8n210g21V<6I
N\j1e?h<B>cHg^0[6kO1gk[_`SYY7oaOgGo?eYG;0?0V:qC5Y92k\A6]]hJ>1Gq@
=:Y;5mSCCRi8N>Ll7IFC50N3_4G]I@99QK2BeWfS7QjMLTfi]84`neGbQE4lLMjB
>Z<K?9ZXS\::?DdIBJEDXJPd]O\a6ajBDK\QjPYiPoB8@?YA`Hej7;:RgL;lLEl@
[SmUZdnXIhY[6NbIMJKCmJ_?[?ea6ajBDK\NjP?iPoB8@?YA`He07;:RgL;l3El@
[Smb:dY46dkoO\_pQ3cbVgT2KhQPS^V:Ah^9`jH1We>nhIfViR6o[a<JmT1oYV4B
bij>6<Xk@AefY_HG_jZJR[YG65fFYeg^e\2;Td<akOWl8OPb196VC;8<0ef_IHMR
K6MgFeMXW^_0@12>Q6\]F\OB6jOJXIFke>2ESf<`A:F;8cPA196Vb;870ef_IbM3
K6Mg^eM9W^_0@12>Q6\]2`O<=Y<@l5R4qO?WTBG7gKOZW[aMZ>V9lT\0kk2FOh5F
OLkR15Vbd:677UOfVnOCVkOKmOJdIm>Dmk7nPg6DEa]38XQmkmDYWP2Ade6J468l
BkaRXU<K]=Qdd1\hAk`keC_c>[1O_GK=YOeEL2`@3aEOaWQFQmOYWglA=LlYE6Pl
BkaRXQ<KD=Qdd1mh9k`ke@_cA[1O_GK=YOeELZf@46IGdOclkqnE[@X3hgn^95gC
\UQFbdA5N94V\]4cHI;X4VE9UgTN8^Xa\AQg4<Aede`RAi1<lTHYXKEEf0SAQmYk
Ua;=OkK>]0lFHfhQ>:m=4F_GSAhF`m>NM^F2H;4DW\77DbLfY`nZ]1lFOPS3PSo0
ll;7OIA0]MoLVDhQ>:m=4FZGS;hF`m>NM^F2H;kDW\77DbLfY`nZ]11kO7e6<Md1
;_qCd]j4`C7ki;PKW3@CKB1X=_Ya8^Mk`A\[[1hGfiC;o6R2VP0cPn^E]m3]06b7
OIIa2f2g?fSODn:4gh2\`:K6oV]oH]]ZUROO31QT@8gN=[>I55;:80Z4>bc\DLn>
YP0CFd9kh15OFA1YGAJ\X:;nnV`_JX]ZUROO31Q]@8FN=[>I55;:80ZB>b?\DLn>
oP0CFd9d[1j]kf>mc6=pB[R@HgP;?>mc@_UCjfD?UUf4Q1cj3DHDO7;cNE6dA8`Z
F;2Y>aQV4o\5EnR:nG508>X`1W><jY;DYo<2>bGndoR7LUcX^em>p37;=i5mGNLA
3>9BO5`4T<6IpBfgI;maOHW<?]4>NCMVe3SYMfdo[gK8?BKF7KKBHID`;IM:nQdN
6lPFSa7TS6gZ=IaoN]Q\IZNeQ=JKblI[WLPTLc\ad:DSDjTF??HCXEPh4Zb`@?M5
Q_EH^Ho;A9S;gB^cNeB@SZ?H0aIjZl@[nfPT]BZeI:DSDjTF?UHC8EPh4Zb`@?M5
Q>EHjHo;A9S;gB^cNiB@1DKGcW41`qC]oREN4<e7=D@ZF]TNM5KNDSHRU=LRPco2
;13CMK>OcAYXH=37H`2TL_Qo@B<flYJbNdjLDEhgbJanh16PTh2`??RjT=a\<ZVf
;2gmAhHT>\;Q7iJG_in2YdCQn;7lFjCZCbUSKVh;9OHjcg6kT<Z`?lSMGDa@<ZVf
;2emAhHT>\;]7<JG_ie2YdCQn;7>F;CZCbZSKVE^MZN^m`p8>@GkgJFJ?F;`>FS<
jKR@J_Vf22UVf[Kb<5S;lYB\MU28HkD3gD<KjaG4HT1O<o1f=;_c3EX19dMcRaQI
POh?AC`mG5=e2FL_b5c8TejCT`5Mi^k:lo1h^No=eCeCnfB8lHndf^M12ON=iPCI
0ONIAC`8e>OeCF5_b5cITejCT`5M@^k:lo1T^No=eCeCKfY8lHnif^MSb93aV5[p
UP]\IM=mW=@S\UjKF^2m65598k_@IOkDE>;SIdL7d1U9\Wnb;IdHUU9X]JQiN_0=
]Y8L^la[KD:?]]BY100^ff_WQZ8gJZOKS2;U[70VP3?Kd\1_4lk96mIaXXNa8OXc
UDE5>[:KK65R=8NF1C0F>f_>TIlOJZOKS2;UE70VP3?Kd\1_4lk9RmIeXXNa8gX=
UDE5B[:Hbd2Yfkf@qENBd2oVnkHA0l=C4<W3jcC<fi?E8Jb_R>jiEP1fb^BkOOAN
6`gonRTdQ`b@M0H]5co7aHK1K?[LGlk=T4G;4_0>`mL6^2c`0FiiET@[4?`P5k[[
[RL;8Pd9keSAW96TREoa:]hc1?o6_ghk54@;cT0>FlK1R28`0FiiE0@[f?`P5kC[
=RL;8od9keSAW96TREoa:<hc1K5l@`4o=qDdZ5FTb0UekTfLPnDko[q]^nJ\ZVj5
Nid<^OT>mj9_cWn?YIb\^1YW^D>a5d8@J^:Kifm;]EbE2>9bY:?1=WfKJZ7PlJ>F
>UoFTVb5fW1TfkZ?=U;;l5JUgDn8ZcOK;b_461?W;gTKh>L4nCaMHaK]hJXQg>9F
F3;`D_657WZ]fkgN33C;Y5SUgDn6ZciK;b_4Z1jW;gTAh>m4nCaMHaK]hJXig>hh
2]<]fE<qf22Q=DgUGT4kNO3U>aDTVONY4PL\ZKKOFoC5@<[D;m9JI3OLZmcfW5:B
T:<__bXa7SLgWJ@hRJW;6koNBkM0mhc4E1oIRgdDFgCe_W?]:6i1lO3BhVi;j<XD
g2X;aYD]fheeHZ`MRJ4YH10iBCMbhhcPhkG=RgdDFgCe?W?1:6i1lO3BhVi;Q<X0
g2X;aYD]fheeFZ`MLIG?ElSQq_a^^NH9c4CUnH[lJ<F;C^7]ck;TDT_UV3i_N@mc
LhgK;jCPJZo3?m4l_[31\3Mgk]4ca?H37k4SloT^Vnim8;\k@I9PU6cT?@j_3QTV
IAZ[NM?J?Ua9RREl=j4JcG\:K_X9mBXM?kaG0h=FInem^I\k:hITO6cT?@j_3:TV
fAZ[NM?J?Ua9RSEl=j4JcGY:A_X9m8XM?k`h[fXTQp^=Vf6O2=>DA;B_^C9OacV7
2L;MV22ibb_]h^cgAHJ3IT6hjK9>H8d75_f]G`acaGMDXIhX`_KGjB?MM2B\jN6]
`_21:M;;[>Teh4NFRBg5O8KdoQT]8O5;KDDZ][N2hI^LFJ94=cKbgFPiDEBQj^H]
`_nN1b;;[>Teh4OFREg5O8KdoQT]8O4;KfDZ][NLhI^LFJ84=EY>n1S^gkpCYXN>
QgjK=O`aHQEXL5l;_aIF:Y:@36_I5VA;RmX;nB7T<n`EP4ci<AM5?nVc1DO9K7OX
HRVl4V7\5K>=Ile=H<ia65?f>gUDCVnj8N0Y6mDOThED`WbOB_gAV>CRWbLCjiQU
Y2al6@5ME[_=ClNdH<ZXOPZf>gUDCVnK8N0Y6mDOThED`WbCB_4AV>CRWbLCjiQ^
Y2H8DVCm]eMpS^4f1EPM2VKeXcFWek;`Y3><<7P_^`U7]R:`Z1E9E<YVR:PQ[QhQ
Fb2[9@^Na86^ka?khJhYXCjU`BFiYQ5>7SU82=[ORmbl?X:3d`47=<OU6=8VDjL7
cVLP;MNCAhX]S0SRfbZlX?3k@0H]YO5ZNSU8D]eUR]bP?X:3=`47=<OU6f8VDjL7
PVLC;MNCAhX]S0SR7bZlLE30<9Y2qHP[k\PBL;S=H]Ync@[NAc4VBAN@HeITg`Of
7WW]^fLR=JYT3dW7n123`CMn6P7@LAc;dRS6Y^=]O\WV_[YkYX@?<ingmLA:C5df
2TJ0f;hT;8Ab[M0A45Hk^PgeiN=6PH6l`XQh7^9;jV<El[fk5`@?J^m8LL_:C5df
27J0];hT;8lb_M0A4<Hk\PgeiN=6PH6l`eQhgn8ZWg_FOp3nEU>oeBNcPSIBFa\0
gLgf@\gU2i2Sg7^ZLD=Pf=Pc:2aNEXAQWlVI\VT`=MA7CI^VV4]FR0nnbF@=ZNHY
iY_JXHeM27`G;7CiL6WAFKfNnUl4IYB?oD2Q7Ke?i19bVN3HFDW_:MnO_K:GEPHQ
iYGJXH3?hC`G;7CiL6bAF_fNnUl4IYB?oDKQ7_e?i195VE3HFDI_:hMgnKLig5qW
e88;M?83gCD^FNBHN_Yqe]Gj>h07TQUkNiMc8\e@i]lXX1dLY85ba7`Ol;\bnXQ6
3hJmU:W_Yfm7Ie]9f`kiHHkAfoY2WkYHioJ3FJE0AmOJYPdI_7hhI>`OS@lED2cg
Tdd4?jMbhkGhVCoYgFiVe;`EMm?@W3fT_OWSFXE03mOGD`5=_:h2I>`O1@lED2cg
TPd4?jMb7kG2VCoYgdiVe;`E=m?;Fcd5UloHqZmbRlj]>d[0h4f<CPa8@\j2J^o7
^YG@oGXoTn1jil4M7eUcOURRG;9Pbn9TXGP4:_CW]:3Dj97^lVZ]a@EB<Olh7QPf
niacPmFonWX04<@l73oDh?LdjC]5WBS2ld2ngZCJ4<:>b9ogJ[iR5@4B>2lh^NA`
Kicc\mFonQX0f<@l73BDS?Ldji]52BS2ld`nIZCJ49:>UAgS?DNmFpScjj?a0X=J
K`>[DD@nl1clO31R5[TQGlDD?T4X5h2R6Y_>?n_iZZHd8TU9R8<]_n=1HZa6>glo
ghO=20NOkb66bOgF22TFTM4K?X:Z_bMU]?TE2\COm_MGcCBEP:CbccSLCF@@Eiln
hJa]05NDk\D6bOY8[:TFTM4K?X<Z_]MU]?TE2\COm_HGc;BEP:CbccSLCFW@EA08
mB<D`>pW1l0a14h@RoRWg7bTmacJ=k;6m1AZ`E@T@fd2Rc9I?]L;l?8L^k`goo[l
SGHGj_dfipK^SYch[:S:6R0SY_;kfN<R8ffgV0\4^Ra?jo<66;MHGZgJW;Xn`4lg
ZD\d^1\j:mFSc9]dA<U_RO]FdWgJRDEP18HmG@TJ2RqA>`]mEp`FfhLd4$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module CMPE4S(OEQ, A0, B0, A1, B1, A2, B2, A3, B3);
   input A0, B0, A1, B1, A2, B2, A3, B3;
   output OEQ;

//Function Block
`protected
L?eK\SQH5DT^<J=RODi`@caLG_?0Hi<@SF_91_[A4lO?mL3OT@S7oP`dGk4?1aQ=
:jG9iD0E_B7Lp\4@NFb9VCAWMP5R:2LVDBU=Q5<naiN^B5A16a7o]ROok62;C\<<
154hXL>c61AY?m1LpV_N`Ef@B=S[gP3UHEH?cPl;C;YU8VWG81?MlnDgBBAhK9H\
d\?<^]XNS=;SPUlC479bT8TqK`7mCSp6?1El_5kIN;HJnm2PBLM\j3\i_F`^ZWeo
1qRPY0dmjVL3JjZn9=g_6WePoFUR2NF_l2ICpGBJoD\7A5<f:^HEMBW6P?i\DWlX
BmO4miDpK4\=;;Bm439H:7dg]XBR5cV8>hP4=UDnV:qCSegFmb@i<@SThcB:QFp7
RLIHFQVWSDaL2Ke<Q7@XYhUV`Wc]KI;kBW=J71b:oUCNl;Oq=_F:S`=pl7=:_[q]
YH@QBMETlA@0SXWS[o[gR4JcdWTjm<@_O1gPn_G\SU7?m?[?IWQCUe:m1=XTGO?I
eGSPCkQLV3J:D:2>nYNQ`a:fj7OboWb2H1?9BSKP=fKIdGdfch?K;ehGRDCjMkT]
USjeY?<L2?9jMQJ>JY5F`a;\;?nboWb2H1?dBSKP=fKI^GDfch?9;enGRDCjUke]
USj5Y?_mB>H;Rcjp@KS6^eH?XG\G9YW<X^NalkZHelCd?PJ4BhBh_UV[FO=8U9k_
?I4l>7jooVDCmNdKfLILU@R45>W4^CFVkg?ZFkk97k?SW3ehRTBh6]AV5>NOH\E0
hh4hMon]_=1k[e0Y@i1eij^B5CdVlT\Yk6?Z7kkeLC9fW3ehRTBhE]AV5>NOH7E0
hh4hmonk_=1k[60Y@i1eMj^HSMS\\oBMpn@k21TZF=mSYbiClcY9A`7D\8gJDKQ1
I:GPDDfC6e_`MjnRJKNSmHR3ZIhGXpoSZ=KCA=a?Ih_6jB[a?eQIgBRJ62^4:0BT
iJh@Wo6dV6R<AknDK8Sl3j:ZElj;@[BO5]hmo=kR6h`94_obbX5go@FjUh;3hhbH
ih][gVFMOk`^Q`;UYci?c=2kF<Co_lo]:7XP?lk`PJ]fCKoKbQggo`4^e[;QhhbH
ihE[g@FMOk`@Q1;UYc2?c=2kF<C7_So]:7lP?;<f1];_^ZpRZ@_WiFJAkikEMX`3
GX^5e6I?bIf<W2VSQ`A1?CN_c1FIhi>O79=@gUZQfR5^0ikH=]N<En=T4K9Cb^2m
H0V1E;QC<l2HG_B8N`LGAnQMJ6_OOh2e`NgOGf>HP_M1`fPR@khRK:8TUH0O3`Zm
a0EKE;Pb;i=HJ_Y8N`L[An>MJ6_Ooh2e`NgTGf>HP_M1FfbR@kh3K:aSoCAAM2Iq
ScJEYjVl6c[[DPbZaV;ZiCnRldX_mZ\[Gg9H1:\8]2=@CJLM_cMQBGoH=BdKOg<L
lTK5R47O5=P[AOj87mN60Rm[KZFJ<3PVPA9dZ7I@[G7lgUW9In<UX9bFEGWQ>oi<
SUe;_XHM5\e^Thi^7lNmiRmW1`?j<JP`PA9da7Ia[G7lgUW9In<UO9bEEGWQ>oi<
SUe;ZXHM6]9VLE`?qU56<B=IZ4>QiIXdj1glUd41Bi:=V@FLEUF:Dq4UUR@6m4X9
gBWh49n[Vh06J1k2[eNCQ;]8;@ZIOS13Un]@4JJN<EOISjLnDc3mL3@nIJ124J7`
_[3l9_DW\7Y9Z24n=S0OD60;;XBKghTdVGLY\EZLiC:fX[KX:f55=745oCL2cG7D
2JL4[\D<\e09Z23^VY0OD60;;XGKghTdVGLY\EZLiCjfX:KX:f55=745oCM2cLTi
_=Be:Rq5GIXH5>meQ0UEcZfbkFJaakn]bQMigC5NRRSRCRgdEmEgA^=FiiH@WJ8E
ERal3;Z]Raa15f?\kjK`6=WPk<X9[3cUNOAoJ0]IER;Rfhl@6R;DLF2lE?UT_G[\
o;IHAB85_BT6li>\bGK@_m0P?<XG[3@9kQboJ0]IER;LfhY@6R;DLF2lE?Ue_G:\
o;IHAB85_BT\li>CZ=ZP4X>qbQM:cFE9Vam:nS6=[F=4D9o3agB[DU0dFODg6M`d
`MR2>KPX6L3[VF?h`=XKbRGUV34_R>c7IAD8n;FIVK8ZGlGZ5E[0XLX?L6DgK9QL
H55iF5V5^TG4\Ig1Ym9Qnm2ObmIE:iRlI5\OSeT@V`8ZDlGXi`]dX?X?L6Dg]9QU
H55iF5V5^TG4JIg@Ym9Qnm2ObmIELiRlUO9nU]:]pEHfZ:NjLiRmhoj421GVg]D=
MSAp8ha9HEe]PY1koOP:eiW3e>RWm`i4Z0H7lN=83LcA`WbRN014SbF2hbVbBn9_
GL1nW9`82\Sm;ZII2gkaWWg1aLMISnYQ0lWiRR=D3?AYYGJgZCVUiXHVFLb5Feb^
o5OL8A\D@d82;HO8_1mjWTg[kLMIFE:I0cWiRR=D5?AZYGJgZCVUiXHV=Lb8Feb^
o5OL8A\D;d8^j;JJ2[G:p>]kOL_]jJiHNbWmNM@0564X4W8]<?^WfN\=[P02ej10
3[ZSLD25nUmS?]WM`BULU49;j;jmm]RNNVe@OFB80lT1Xo`NZY0]]H==PKBWD8\Q
7mZ_AM3TPZkV@`?P1l]KC>hC8K;3W]hT40jAmFT8<6T1kkVCfY0]]H==PUBW_8\Q
7mZ_AM3TP9kVO`?P1l]KC>hC8g;3WJK_\Oc2\p=;Ui=57B7<Ta0V;D4k1>mL;1D0
5KGbGAPP^b\cNDR\lJhilVkZ72iML?aikPT0Jol]gP\I[>4G5\IbWAO7QV6fNdMF
1ED53d:U^dLj>d8;W<^K]<`bZYT4OoLgAMD2g1=S;b^hS44EUojdN9OOQIMfNP?]
ZND53d:U^d;j>C8;W<^K]<`bZY?4ORLgAMD2g1=S;b4hSn`H0d87\CpD^iTcmUI4
ciJBUVLY_JY6[R0PW95RNpafKUcj<1aU5<HoTNBUF=ON\NIP=e`8iY59c@Ga`:Gk
imDc`H<nUZPbmIXe=ic??QRg6Z?W9Gc;h;g8j\Xh:AfK`Po2QM\ZhKn>cBJ5leaM
?R;KK<:@TTh@n?lP8ShSVEa\KHhPhfc[R4?gLLXY:9:K`]_g4M\khKn>cBS5leaM
?R;KK<:@TT^@n>lP8ShSVEa\KHlPhTB^<5cIJ8qdomeoaRZ[;?6K2D@QDDHSTU4Y
]9lCRKHao@CJ4PBFoimAVJC`<1m9a9@L]Z\]>n[RKY[]:=n7FI67C^[^We>O_gmA
d9?TN`m`Y@NAPJ[eUIK]365=FO[VmjlYV2B=`mfdO`3MFfg7LUG\_SA^he>S_gmD
mDST9`0`Y@NoPJfeUIK]?6:=FO[Cmj^YV2B=1m<dO`3DFfcXNgGJkYSpoO4?UXJ8
0CXePQ8:obO7Hfn^iRXZi4`_Ph<YS;3:6J;m3dJn4OgTlW9\\:?_a^;QW2nE2n^a
nd^0K@@T`EN:ZN55P]^42Z7o@0<:B6[?]6?5:KYR<mBT=nNR>>Z5EOToo[99o8Pd
n9@YB7]f`3NdHN5T>bmb2K7k@0<:T6[W]6?5:KY3<mBTCnNR>>Z5EKTlo[99P8P0
WT5T]2BYq:RddN`7hW@56UB@PNm<l];I?olT6TX3b^RSJ2nXicom8Eh6bOW=VhOR
ZjiKD@iahVQRP<^1o><W_C5jKmfT`4>`41dg^=dm_VWS?l6bVb\km=QVX6G6:inV
UTY4HKUE9:X9N@@76>0EW2CH0m3TZ]>`GG>fc=dm_VWS?`6b;b\km=7VM6G6:enV
]TY4HKYE=:X9NS@7XE@Nn5J3[q2KA75P5?AOBiFFcZ9OA3Q7lNF=]NC\>cBNNBAY
RKegT;5^QOF<g]P:S`RTY4l;\R;X\hmELoJVX4B_B_lGBn]:JjH9;km5I8?ANL6N
m1bh9i=0PA48caD@YT_;[2A_9j2OeQXVW4JCf;<mj:l2B?Q:JH>`ehm5I8?ANLfN
mDbh9i=@PA48ca:@YH_;[2Al9O2OeQaVWnUW5NYlTdp:RX3E\ADB[5W]_jO3Xb^5
oe6DQV7eCo8J9?S8T_KeGD^C[hE=[B29iZ[l^kV9E8LR_O:XbHAcA0ENWoDeLNPI
_V_ggi@TK35p2^Hf4blSc3Z`cWFof5[Si`lLaG^G@i;A@jS4c1Qf_loS;^@a\o1o
KlHK4UoAAEPmT?kb??REP0\Jl?=<kD`2i[2d^6Z_ZaUkSQS8EdoS8W^SOmZR]7\f
MW_XMX7MkgZX2oZ`;djDPf`KN[5Mkn`G=72H?[NkZRU9SQS8C[o18W^SOIZ6]7\f
mW_7MX7MkMZe2oZ`Cdjam^K;me>]qjE[]VPNhR0>?\daGdYjel3QLbfP>n4lAR>4
nGnfcBjQ6O6b]m_fgTljhY>R[WkcPQ<;X;bH;eL]_Q^T2endOl=3`@DLl6i]eAo4
_GElBJm`S3H>X5o12mjlfVkni0kRYj4lk6E0;efid`<OWeadO<_3;[b;j6K]eAo4
_j@lDJm`S3[>e5o12Cjl]Vkni0[RYj4lkmE0OkZYG=YWPpi=bfb_4B@XW@GRY7jW
a1@`6mQ]lHQ4>FO:QA?jp<Z?5j:VUZ8>4AVebVh6HnLoGU<?kBbGY6B3KO1[YR<7
HOSRS@;FoG7VE3`ACdkOJ`24Z1N:Oj<kB@M8?Q;DmnB@m9ECcjDY>?a3k:K<GX^^
7cN[CkR`W^<ciWAF>Q;kA<hbmU:^jjhY3a?IYQ9DOFe@bA1DUjDY>?a3kd8<JX^^
7c;[CkR`WQ<cmWAF>QHk[<hbmj:^jEOgWTPB;pHTf=JDP:M[MHNV8F5aZZG?>d1Q
7Zaj2Jd11nCmUMVEi^fK13O8SkE5EWiglNkU5JNT>X;QC@<4oMD5ocDUU3GUW:PQ
]5emUHl316VBeZ6KT_X<?R6\SbK`cDViP>LF@NHJ4VlWlh<bX>gATID@U`0VWocF
KbemUHl316>Ge96KT_XJ?Q6\SbK`cVViP>L=@NHJ4VKWl0o:<;ji2;p31POoE@Pe
:=h49h5AF>0Df>D^ie:JgP98ZG78?G=JHnSiD;84C5=EC22CAo2da<GX`Vfh6;d6
@U851mIb:3h4@5@kO9lk<W5GMG4@jN4BQ@>l_X?c_h?Sn?2J4lW6a>239`jW3\I6
018_ghbbd3aQn5>ef[Zk<W5GMG42;NfBQ@>l1XIc_h?@n?oJ4lW6S>T39`jn3\^;
HXF300XpY7CU1oA40X3T7VFLcbaOogG1X_1YUU_]G2gaWL0[Eoljj1op@^9dIAhX
b7UccgYPLAPXa[Q3GCF``4b`XiY4Qm@8M`hhD?bITd2Cl[MQLQMFf:KXQ[DT6FCW
21TmeG@h=SEBRRJhgglNH_HViTYhbBKF?flXX7dL5<e]RWg4FU>45iW6@ljfAdRJ
2Ro4>EOK=:EBYdJXikNGH_HViTYhO`KO?flXXOdL5<e]2WghFU>45:WE@ljfVdRJ
:P4OnIO6pDE_?ndZYXV]F`MCVcbSLY1i9]0KIBf:YXb;3hJNNBOVEaMYZ:B?ULm\
\hcF[T[5Ic9CQf0M5]@IZ93NcCE]VA9EW7VVoBSRZ:g;O_ae[l;mP:8K@^oYO8Sd
h8AMeP[R<DAn4iJ`F]5Qcai6kCI]Vj`E6EoCgBERK:g;OH:eJl;mP:iKZ^oYOISd
?8AMePWR@DAn4GJ`[KeL]ckZ6qJWJ]iSZA93<BQgnSBJ4:Tkk5?>?dj:JEldTRmT
kmJYk4k[R6B[L<i54`Q7OAMYiD;BKRW0KSFTZ`^T_92?K^n\HDfIdFZjbmk5TG0n
Z:jSmb?FWnO8\0b9>KE6^AJUT3J\e6^I_bFB7XO\m`2CK^c<HQ?5ojZgbUk5TG;S
ZWjSmb?nW[O8\0[9>nE6^AJYT@J\e6CI_95ZTIibOWpf9>M[^R3<TXB8`GDb`GXc
`m[STT?5B3albnM^IMJBIK]fd@G\6bNlVPU;oQQF5TPWi3SZK3qXZ:m4FYeOaT;Y
PbDKV=_ol[?WE_AMh]WMnTJC^6A;97ZK4>[GGAYTJ4Zh5@CNMeE8@hIOjl[]UJ_n
Eej[5H`oFQW?F8=@=6<T`TJT]iK2cmXPVZhAWb`P]A9o58@h9DAXRMmd8_5]ce8G
SfC[1HlC;Qd5\Rb@F6<T`TJ2Ui82cmXPVZhAWb`d]A@o58@h9DAXRMm28_BEYeUm
T;Wq[M9o@kN7a;7:l:@HR>UUGnj;82^DhiVj?T8:XZfW8;5bbk0`P@^Ji<PJZAPJ
OZDl:o0^\iR\L3hUc6YMCeRQG]1[V>;<L0X_`M8KACJR\H^1aE[S_][=gJ__4j\E
GK1Y[2Z@=dVSL<2]H7@kCKRe0@1a\9AcL0X_`M8KGHJC\H^1aE[S_][=MJ_;4j\E
GK1Y[2Z@XdVkOK9_g`hVqnR>[k?A_o0VJKNQo<?\23Q=RE[<3TZMHZQ5>bWK`M]j
jSa^@VhI@D16MP5iS6m\F<@6i9>HU3b4lbee7lF;8bCnJ[kb?eaHkIi5KeHP39L:
870^0PjkAFCa30<R]dm8nn??=cCMZ3NRnB?b8l;;8V9n`E;]_eaHkIi5K14Pf9L:
870^0PjkAaCaX0<R]dm8nn??=gCMc:hk_;LgoqFK43OYOjML][9oc`?cC3_nY:a]
3E=>Zb5EgQm:cCTWo2<eBWQ24:]k]02_6lQKDQK3g4oo8;0nj5R^5^@g47_h:mfo
jKZ[LGkRgl1`b?Tj60UE7^>C2en8TOTm:M`AK6F6_FnciB0QCmm_^m@e4WL6:UQb
BlZ7LGkRgl9;bYTj60UE7^>C2eh8T;Tm:M`AK6F6_F`ciBG2ol?aE5pNHS1;mac0
X@29I1>>aZ31mg38mS\DGbQld9A2mIL01:Y0h\WBE@U`WPGMZcnQRem9WS?^^m_S
Y<^Vho13lkccjTaG@c@jEZ;eO9RKNn1:=ScBfDQOo><_4\8LFS<^RRPNDG19m?8S
K=]AjEc3Yk4nSTc5SH^jiZ;eO9RR9n\:=ScBfDQOo><:4\3LFS<^RRPNDG1hm?84
GLiom56pVPR=4f>gY3gPZRdo^Xo9Ai>AKZHjPIf@^PWb5^?5nCQ0BYYDI?_gE:kb
`B\9EVK?iYj:bOXQWN<^>^fBXH08AWDn<gQWYmo4=_WQKOE;80_U4dPNVen\UcTl
iM8CodcZVfWJS6;dWZ>8DjHmXJ0U_SD9lk`FYmo4=_WQRfER80_U4dPNVen\lcTD
iM8CodcZVfWJ<6;fel6DdOBdqidMh1IKC;]RM?c>JP0a2D<W5@TkmbI;MlYPW[SE
dAM5HC@>@<F8jjOhM<gBfcaAVCEU`Eo<k8oaY_5>:k_mB=fCFf\BX0TB;aGPN;BM
@61>nGGQ^YWcdiXn<a@hDQQ?ii7TNR8@78mLD2MjYkfm\7bCLT^P?0TB;aGPNjAM
D61>nGGQ^YWcdOXn:a@hDQQ?ii7TNR8@4a=e7b]RipYbnJeNn9FC@idZ3kI_Gb1Q
l[XDVk]BOm3?V[N_`B\D<JY8IBBXE\a18O??L@WWJS`dRgAnd>UOQF98kDn0MGVj
_]<90F56Io7:VLASeE:@Z;HY<=1:>bUP__Jm4OnMHVYj[M2E]aUN1@KD1QncMX>k
_eCR5a55I;7:VL9heV:@Z;HY<=1:>bLP_VJm4OnMHVYj[MDE]Jm55YEUDJp9B;nM
?6OZWblDH;`JKD3A_8842?J^>[V_c1Kf>WiRhoLfTPj>[`8=Q1lHic?lYXS@iHgZ
;1k=[PAPO\ml0^LU_M;Dh=FDnV>qDP\DPlomYbcXTn]MeDjdRU@;[=_pIbX:77KK
ag7D80EXJI@a>nZ?TJQ>gi2c?]Vnf;F^LOSJJfjh@a=?I_eFUB>hPd[@SQYmNLBi
OCP[k_^<2`_<cMbB>0_\2\QPUAVGBMhhe\7YNYe1Dk;F;FUg@?Kc]decIdoAJ^eo
Oh<VJ?f:2H_<PMbB`VXo2dQdUAVGNFh_e\7YNne5Dk;FUgUg@?Kc]decIdoAH^ek
C6EVdoj9qDZBc_^WNHE8NU9R8KR_OB1HY0YU=HcS5MZJX6UBKBLLgoSIGTFPXQag
D5:WLbmmeNEEDVS`R]oVJ?JOnKE@_MbF?a6IgdQ^i<kJ=M]7Wf>HNcbBRajf1JQP
1gLQ;:m`3DfH^8U1Z]TijSnmRKT@Z6bF5=8?RdQ^i<kJ=<N7Ef>HNc<Biajf1GWP
9gLQ;:m`3DfH^hU1YmDhBB\^;poXkJ@=gFKm:cn2Sa[^JG13b9cUoU]4mL;aZK5k
T`A?`PY<6SBg\7384F=\`Rcm:=ZlOjGR8Q9[JjTU[k0\8_:0j2_3gWXLJRZAZI`;
TZ1:JMjbYGZZN\g[j]SDAkmmRko9oJVVD69\jaEjSf0Y8_70j2_NhIXBJmZAZI;[
Tm1:JMjFYeZZN\1Lj?SDAkmJRNo9oJ`VD62oM1J;Tlp\bZOI]hac83P4nf>l4\j0
e<<dAT0^\BHJemqXUK>i^lD[n0\OCG<ZTie`kHXOE`WC?mW:>6TRRNX\m=4Ii\i`
YDZDP8<GNfhN9aF\_MQnPcL_F5_fc@NB5>8CE0_YS7MP]Sm_L6VR_>B@j19?8@lm
h;[MB>>RU^?Z9`lX?1\XBmL_IIQMTFOBo>8DE09:;;EP]Sm_L6VZJ>9@j19?>@Hm
h;[<;>iRU^?Zm`lX?1\oBmIQ\;IBRWUq?QZV\dPR06Y32MZJcK_oWon@_>c6hc;m
UFN[@OfGP4O1P0BbdO27^B77f1XlnC4Z98I__]N;8HoV=2RhNY[n^^oNQ5=[<4Eg
@RNOoYFb^5ZF7Ol]F7Jb0hiXoRRe5C^V?[kflPnM8`[A8O[^NO[dS^oN;@]@<4Eg
@RNOi<FD^5ZF7HleF7JbXSidoRRe57^2?[kf>PnO9EEo3fU5pL?bOA^BGO\kGY3e
N3U2WRmTG_>kD5f5[;lnS8^<43`]9BU=M36?nnnkW9P[bVR>P=HWnOJTIUK39IQS
Lf^CC;[Ee3QNP<DoTion\X`^dm?Go`g51EQCKh5I_e;]b_RmRL@ih_SG7Ua3^RR^
4fHCLa[Ee[nR;<Wo7ion\6H^km?Go`355EQCK??I5e;]b_7mOL@ihlSGL5hS^RZ4
Jq]_MERG9AR8][H;DN5n0K_i8IHD0aS:5M=B_KCj@m1DoO4bCMBLg78dT_\VL?XH
7IB1EHJnfHo4YK7Y`O<IjEbKH^S[3YL\c=dJ_fdh]6^Pb7oQP[T@N?V5NanV_7:H
:m]Rd]Ke[5o\ke\dZj<Gj6EKH20h6kL\c=dJ_f>F]8^Pb7o>P[T@N?gNNHnV_7:H
:m]Rd]oe[0BlNedKNAp:LTC6:K63A8lX>KN>3cea^1R8Td:_99AM\PSmhAX1QH[h
j1WLT9[Gl2AA`cV2\i^8d7cd1Ce[IfWZ6YT[I1_QX5:[lnhVE4<:jPkMF?RIeDhS
Xd>W?m>JdnH6XVVQ\Fm:>YghR@O[44k4NO7[O1_;X5g8mA@V`4Z:jPk0a??IeDhS
dd]W?m>7SnM6XVVQ\Fm:>YgnR@I229QQACCqGXcil<hlYQHh1?gC[jeVN5^<jHbT
k6d3NEA4_eViaaPVKL?eQQI0I6g<fDgYZ5O>gfVQ?cUaEbUNH8J1hGdaZLGa6EO3
\b4Nb`A[o3i>;^Bdj;MQTO_oaf4`TMh;65fYG]dDShD<ESC:Vif6hkdP0LGa:OgK
\@4ib`A[A=i5;^Bdj;MQTO_oe04]TMh;6gf0G]dD^hDhGP0?PnM\qmOnAeWcjSWn
T9mZ5C;fLjh@?qh1K\jU6b<6YNE;ml99LM;5LTgKaWlblO4;?=cDKf_Ff]4YlLV=
oD<m<jCU=8k1gB2R>J58P>NljHaCAHmjjSAS`XUBiT?^H;YM?kDfgiSMPP^g3H4M
jbf2M6LEPh\1WThK_<L<?LNo0UPjJLm@jgCS`8f^\O?^H;YM?kO:g`SMPP^g3H4M
jbWTMmLEPh\1WThK_<A<?<0N26XAI;qJIiKF1OfFXa8kTFSTi`P8bjn9i\f9FMW0
NbITGLcZe4;kfC<^?8C3\D_mH5]mVCA<2o98@[lBVe\f@YcR2^FC3Z_1Z`jN^JF\
]bWH_PoWGI3QGKif_VIX01;Z@iOWV4oJiL2I_b8B_HB;4GKRX^ST3Z_\KYhN^JF\
]bWm]PaWGI3QGKif_VIWW1UZ@iOWK4iJiL2i_b84D=n7AbKp[hO0m_eOPm5HQ3ED
IE[TW1hXG^NVf\cU<JG3>V>Eia5b;5><W?32Y9[e@cGViAe=>VkNh;7<CM_>_E8=
F\=@femRQCk<no_D7>Gb\=JMmZ]eGe<\XAM[=Um\8NYN^AGm[JWje7_BCYjcRe05
FE=4=emHVQKJn=_o7>GbJdJ0mZ]eGe<\XAM[BFm@8NYN^AGm[JWjn7_oe5nWEARj
pom;^JDiG>LPl<?cBS?;Cn59TQcG6`cW9DQ<ClCddZ1NI<B<7]AWLY3]_03HflcH
BDiU4hnFknh3Ab5Y:`NNP;JmP_]GoTl[O@n<P=\a0]O?gn[HI<cBm:2fj>oZ5acl
mo59?V=Uln\@oMJEj`@NPYJmR>OmbTo[U@n<P9Ya0]O?gn[HI<cBmT]f_>oZ5acl
mo59?j=UIFT4[]4@hqk2CI91lFb7SJ0SCS^W6:4[SA[H4?Rc^DQQjIG;M<qGAVWV
170O3LB?O9SFZU8dk:N<kT4jkID0cW2nBeVS4@UF6VnnN4iefn=P>W74YNkZ\^YL
<Ue5PmIY;SnBT4Cdg<Xm>i\W;RIMHWod4]<4CBXTk:QV?Q]6VcGljB14Y_`G^TLJ
A\i5XlRK^EHBO4Cog<^eebFW;RIMHWoZQ]N4CBXTk:QV?Q]>UcAljB14a_MG^TLc
A\QL=>NYWU`q_m;2NmGLIca?OdVB`M_Le2i5JlAkfH4dSZ>SgnjD=@TQc;iaB:[Z
<kQQUD4SOVNhEBA\f8N@872VVTnAoh?M0H<J3ZP^C:?kbd>M]>WJelKmJk:`Sj5W
;9GmhGoA@VE?_;ThkEhZ8AIX7Nd5o[?m1H<JF>XDC:?kbd>M_fW`elKmJk:`Sj5W
bEGhhGoA@VE?_;Th;EhRK<CSgP2Rq?@@_e^SMgHFmmNOVEGUEJBk_LZTEiX;mP=[
aQlJ1@AE9N\fWag_`Q0cUTE=3f[?GZlT0g=Kg2fNJ<Ql]8eVj`:0Dbg0OTc8EjI[
1doj_9[`jGVW8mJ0^XLaX33RB>[GH?lJibfc\2eWNE>A=8WVSA:0gdbg3T88=jI[
1nfjI9[`jGVW8mJ0^0@a^33RB>fG=?lJiffccE;;>]7h6qT1L<99N\>5i8`gKbhW
JTdP;jZ@R`LKVj_MPkH[2M`h:ln=6n;5UKa8D<I5;HU[oOnj:HT\`9Wm6=Ja:YgX
2i=5DIPafNO?E[pf<8agjf5@I][3^`mVo28__d`V2P4GYo\5FD^Ag8dmJ3:0>lcm
WGmnVg[;g>4NL8N:la[7aLMIjlI0K9R2gCAQWTk1iTU9?R683D=]TB9bfBOckPE3
A7^3k0QSDH568=[fMNC?o7NINnL>3:82cC;AET4DYe]9IR683D=J2BKbfBOcHPE3
A7^fF0^SDH568=[fMNCj\7UY2mATSIUpK@?l6X6=hdR<>ZHdcgP=JY3hY[XSh6B^
`N;j3aQ`\M60e@hMJ]DY6iY3Rb:LYXU^>g7_CD:WX53oe2MB2:3?@YYTS_dP\ini
Q?;V_\Q^cjj6Q9;IWo\d]<A<?JQhiHXBKNS_5TdWXQ\D707C2O3?l<YL9\Gl\ini
Q?;VZCQbcjj6Q9;fWo\dR2A2?JQhiHXBKNS_jRdZfjCm8T07pLXI8UN6M\iV9gbS
n[X>nfZ[o?>=P_>1FU6=HZ@>nK73lZ0EX8`JL6E2hCaUBYTN6Mn9\89PG>>d=O:?
k^\G_f[AI7D@IL_ZK=h=oRDoVdc9>V`^Ge;3^:m1Nn1Gm<0]YL1e0?cSU>;GS@2c
R^KGYmbA;5?nbL4ZR=h=ok2oedc9>V0^ke;3^1\1kn1Gm<P]:L1e0?DSZc\_0]h;
Rpg77=MZ]dmg4IYm6GZ8eZJ^Dk7M?9_9faGTn3ScY`bJ3bYHfRWRkX04SgRgmIF0
Vf6PUdDi>b5H4c8bVo2Gl<Jo@CdjeMkRHcLjn8V@`040]Ya0DccL4Y9`9>9@0EM6
YTg6`ehon[5I=:e7hc2bl<2l@^`71RkRHcLjn8R=`o40]YalDccL4YcW9C9@0EMo
YTg6`eQ?n2_A@bLP]Cp?<>EQ?TJIVo:7\mRIZeHIB[kLfEjZR6T8Oh1DD;Fn:9Mp
SKlPfR1V\_:jXh\ij6IJWaCo26?N2fIJdeE@Idc_O9EkPgHYaGib_Q?I3<];KK[G
l?6]OFP;F=K12KY^nWTU5X:e\X_XgI9O1^EA=lGH05HBijV4CM@faOZ?]G_\<5JP
SEjJQ<=XF7RB6OTCnoTU4[:iKd>\gI9O1^EAKnGE05HBi^VWCM@fmiZG]G_\<KJ^
SEjJ1^=0AR9h:0Xbq62nfaHMTY`SnD`Sf9BNlG^d2IcS`6\SeN7:SPKY4=LC=;Ih
1^DSKn<;fcT10]:1\ALHmV5_^@7g>VR=TPNW1mB>n3;2JlU<ffE:iOA>Eik[9BaY
>E3[k[IKPei873B016d:KS1@f@9I@K[[iP8W=2H>C>_6[l[<0fE:iCc>Aik[9B=Y
>E3[kS8K0ei873V0T6d:Kec@jb:gMFMC]q1<3AQNHPXbTbK1b?XHMn0E68iAhSae
0dbj\bn@QZHTP`_lnAfg>\=E5JWVW?:4BLO1WCH`_ljgA2\llmL3b50AfKGd<CiW
G6>6\:f:Nf\eia0PIGQZ]B1A?;E[GdIdEC1V5B[gGCj2L]>VT]L:bg\GfG=Y\diW
G6>6\:i?NF\eia0MI8QZ]BAn?CE[GdIdEC1V5BU2GJoWe=l76bqJ\]?JO;J>\l[U
N9`aQM<<XRij@c=qjeYaedIcUG=6A`gmhTh8;;@?<?]9Q;0:TK1S2OIl23YjUD`4
?\mU>BAYk8<KJn4Gn;13ol0=DnHLbXGKDPAW;=gS`C8RUefV<W1Mm>WGSU0^SML;
N[K0JmRR^IE1B?B7jRbjgA1ND;jANo7iDoAWoegSBjjUUTfV<W1MU=WcSU0^SjLR
N[K0cKRA^IE1B?B7jRbjE=12;=FVGoGkpaKG\S0e:3KZV=]j\S\Y]<KUiFOY7?N3
JK7aH5Ai8N09kBAHYIKBSThRUi6<;75WC4Fa?W`M:26l8DWd08C9n1<5f5^N4j1_
=6Ja`7]ECk^hQjOWX0f_l0N6USEKWE2>laQMPlk=42g6860VA8j9n]=5X@:4jja_
=6Ja`koE[k^hQjOWX0f_lm>6GSEKWE_>WaQMP?<==6ZPATQ92qgbTKkof]bn]?o]
_Yd0DbQY8c^BD>QaM1f?46Kn;jUk\V``5MNmMf`<HZ@[\\Pa>6NTKLT=HAJ_N6[]
EmTaHF\aaK210DQjeS<44c_G_fU?]GA\g7J15ef3Raa=ECc>F@gH9^WeFOJZRB<9
2`TaHNASaTTjVVQjeS<44cVj_mU?]GA\g7J15e;ORia=ECc>F@gH9^4iFRA7jCdZ
hgpWmW[FAZmfm]W80NDU=G]QY]P4F]@oZcF>f:?P9AWC8WbnePLXoDYW05FN?IHM
EZ4oW;gaPoBYJC`hZK;l3:^n`0CA:938oPUdW:_NeDICG[oX[=XXA8kN7@hS8^gj
m54WH^Ri3boYnfF`ae0ld:^7Z0GcIPj8oPUdW:_^HDRCG[oX[=XXA8kch@kS8^gj
o5kWH^R6?bNlNjPnhH1pJDHLo]D_jKIOP>[S6L:dO=N_`P[1XXKDkfkYa9lG`GSb
4fi1P3Q1VYR_bnYZC`NFgV92P0UTV7L4cM\eJelBOL=8IGTAXIDec]k3iT2C8o]G
;\3Y=1AeX[:2NhV3HjZ^JaTZfMchVeP]CMMGJ9lC<9=`l^A<XADec]k3dM2L8o]G
;\3Y=1Ae7c:ANhV3HjZ^JaTZmFcMk`DTJLecpE28JSA__7IgRfK?EdN`1:G2G@ml
^bllm<JW9E=_aR\4hZInj80Lo=S^R7Lb;3KmTl:_R7NMKWGX^ce@\]d?29[^>6`1
BRM]K2\W0KOONoE\O4^\jlVWEOCo1<<Nl5<U7EOXVlY2cWPU[VGi;]`?ZH5^Og28
kRi]K2\W0H8O6oE\O4^\jlVWE9ZoM<<Nl5<U7EOXViM2BQ?>:7go]qk934K3`L:N
5;b0_XTEHD1Y[iKCIRXa5SKCA8cVAq4iX1YhAd3>T`3ca:53=F\PoJPIgZSFRE>o
4FZK9o>kROZX;]??miUNEMH:U7UKY@ISeb]9hDEb=787YB\GH]\`Rl^5Ko[7<\CP
4\9ijBdaeE:QN][=>:lHGc1AL9Of`54DmVcZnKERcWXCcE\6H>^eR_1Oac[7<\CP
4\Shj6daeE:QN][=>:9<G61AL9Oc`54DmVKFnik^8L^UGgpK_hAL54Koc`W]KHEU
cXm80bH=5kJP79gDnDXOLW=P\NX_]HV>XMmJFUi52hdi90im:\=[1aZ3<a8c200k
1gM8H^<MDfN3i[5<3DPBbOaFZ[iTcoGJdE;O5h;CXaQHaHLK=5WmD8n3?JA?THOk
lgM__^JCUF03i[5<3DP<SOmFZ[iTcoGJdE;oGh:CXaQHaHLK=5WMO8Q?O37VhaZq
aLY4?1_\lD\=k=Qd9YQPbHLPEVNL`L43j6fPHcbXQlB`[A6HN>nFd9]3WJ>1mWdH
9RjS3=J3IjYfB4BH]TBFbe<[b3fl=6dR4Nff22BI2ac@8Cc]g^2B:=ALQRN0<I61
a^QRAR3GI8Zi8cQ>]7BH`d<VZaac=XdR4NffSKBJ2ac@8Cc]g^2Be;AlQRN0<K64
a^QR=J3o3l38=feYq\=A:gWB<XiY_SAa3>=k`KX]EX>WGA53k<9LVDWhWFNj0B`A
<]ln0RG]5]^8nhU2_V<K5cSkh^[1LWf0\2DX1KMY\:QT`oECIp6NI\oQ3M3BS1fn
9ZNnFh3ghDf6RkeVoe1o<?D76ea\;]1k6n6efFolGj^iRXX[^_Pe>NTg^37L^TFf
Ikfk`6K@E7dX9ID?E[6=<SIZO=LZ83R8LJWAW=<F[;eagf]6lH6mZYj?ee72I6<@
9cf:`LWPEa]?GSDNEF6=<S^jOfLZ83RQL`WAW=hc[Geagf]6lH6mZY8[eXh]C_eL
FYqO0g9adgZYij5ESVT9R]:K19XQ97MFbBF[SOG7[]YXgJ_1MUDoXRAcM63:5QWP
B0LfomjZoM13cIDa\je<No50ID5\\5i`HDC<DOTn]fd18d]2llgBX^[bfYn=VEUc
E6VOb<[6jJh3Ll9]a8o<?ohKjDZR@cD`lDC<DOT^=f218d]2llgBX^[^1Y>=VEUc
E6VOb<[j>JOo=gigjC6p>Rj[6;=GcnNfO^p:1[R=o=@9855<Z9X`jPd`_1:I<ZjD
FZFdh@eID=Cm=MYVc?KS1AH^3Bm5^X8MZn=@2gMd0fH_E;ZDiETaH0Uao<W0O[hY
o`TI^@gYHh3VRafBF82R0[bKBi9`hk[g4L7:od1D9R;_Wh;8WL^a:0IIl<`52lIY
o`TI^@g]?h3VRafBJ82R0[bEEih`hk[g4L7:od1V7R]CXo^TFFjpRM2DGbHL_`3J
=8nKRlITlWHGkBa`d1]2J6I>hf9Ym:A@UK]Vlh0A;AKI]:6eG4c??6hnf`_>U\g[
e:R3aF8L8=N1Be251li5M5I57NB03i>8Q`29`naQdLO8QY_K9nakRUHDVJP2U5E`
H3gEaI8Xl@N<S<U>1li5M5I5]QB53i>8Ql29`naQLnO;QY_K97a3RUHD`FPfBb9>
[2nCpl=;P`UTRhAa0EIRc@h317FJ[6`4bR6GVGaS4>R37OGlj;cg1>`1km;J;ZW2
oamgdkZFR0c8HQZoW:KB@UYd67N?2M0CGS?ekoESPe6GM8=>`BQXm:2jkmE[jTO4
^Vh]gl_G2SMFNQg5;4H6bUVd60G?2KJj5S?ekoESP21G]8=>`BKX`:2jkBk[oTO4
^VW]gl_G2D8F1XB:5K69<pcnP`Ej2<G==2_VnpO5Q<cB0\K[5NB<F^lA2dAb<N<a
o`8l6f4heZ;HU6U60RbaJb\TLPdj=>ScLoTaWRTXVoPUc@`408W1o39nNN<6PZ]G
PdmWPe9[eQX3nKe`TGI]8VG2PYMHcdCG^gYl8iOM<@G2h7`_Vck_V29UNNAaPgmS
5hmWPe9[eQSgnGe`TGI;8YG2PYSacfCG^gYl8iOM<@lkhLnO0<bb?ipHhVNDT87P
^f2`iSS`DJTVLo`1dQaflk5o^6PZVo_d\cDNfh?k85Z=ilVR\<;O;34C?:bDLT\Y
mTQRWEa4^GFUFbWV1RA[4@eCD6mNkPf>mOOO72WjGldg]G`oLMgRl??H6>fT8UTY
9?h?ROP4fGFnUbN>GMd[c@[CD6mLhP6>mOOO72WjGld;2GmoLMgRl??H6>fYEUld
HKKNAX?pEjH5O<B:n>T4h?Wk`lk]Hjb<_d5@WSEIHGH5YL3ED>@GidnOC>J6e4Cd
U7V23L_;_BJ\_CBHGKEXaQhmfY2?E;WHH=>gTJaaPOH1TZLkLn_B3fJWX:14SWPS
70^Qb]OdE`j6jVRXGC0Fl;Qmf@2[HWWaeHFjTiaoPOH15dLlLn_B3OJeX:14kDPR
70^Qb]OdE`j6J8Rn;aPPk[?mp8_8_BH0BAa6WdD6RUI`I5hJHOBi8TKYWnB]^c=f
8clVKc@L@Aj^:S8>9S77PQA87B[1BBO4Ni:DTYOOK8>Cc4n2aZ]f[VR^fXG]0F]i
QW4lO@0][Al3me:L@K<TDbj@Y8_<bg0`Ti2od^>Ba88Cl9g2I1jdfVR^fXG]0XRi
QW4lO@0][Al3mEdLEK<TDb[@m8_<bU3`TXha_mJlKpW^_k3TVl>n;XPRaPZ<3Y1G
XZ2`STUDSkBP?b`86VBV8X1nGVNZ6^WZ2hS<oB=SASnbRYC?TMSl0FJfc6IkbNLN
Y\YZ4IM=mMoQ?Hc3ZRW@ClR3PfRcm2c?g8Z5<7^R5_WLhlTmETSR@0]QS@I=b6[h
YPD`CDMlmZoQ?HdHZPW@ClR3PfRcm2d?gWZ5<7^R5WWLhlnMEV2Mc0S8@4pFm^_P
bgW=G6HX`eV`>Fe9=R5QRXK6X6^8XeD97i_U`hK4@1gW43jZ^?7;Bgbmf_WDWcjb
e>f2]_I]WTCn^\jK`V9jdWk6n:b]Pe[kAF>P@668?QRmI0^<Neb43ZXd\e[Fc5NF
[A:2lk:B3hfn]\k97V64KCb61:3]Pe[nJFNP@668IQMmI0^fOeI43ZXdEe[Fc5N]
JAD?9oL[nNZqW\J76JK8;@AO?H]mW7kLEgaRA@eeKe[?[A_<gQ`n?bAhIEOZlQI:
nJ3DE]m\MVELBRSCKSR>Fh`?L>NFJ69U8A5PX_J[1FBEVE_6j_V3S4f8nXRkHOY_
\in]VY:3ZGA[WdbjaanRF=H_e6eXJ:91Vi5Qgm\31FBEVE_6g4VaS4f8nXRkHOY_
J8n6VY:3ZGA[Wdbj:InGXI7VMK7Lpo8c0kWNmYBc78LRT4odhGh?VA<j7=b<j>\d
CH7:BWQN4;<qNIU^Kc0>`5H=LR]RgHgZBQFYC7OZQMgI7_j3l]fG^lmNj8bDmjEI
15J^0W\f\=a^2KJOoU[I7_`[O3XGD8f_P9gHm5gO`L0IOnjkPT7=g\Hk>oiMV[hf
?6OdOTX8S8XBNJ>nNQ<;7SAQ4iN;DFf_B]gWCe8M`L0IOnjkM97Kg\Hk>oiMV[hf
5`OdOTX8S8XBNJ>nH2<Y933\SC]gqb^l=HGMBfD>gWdLSe`\;LOQ_?;m46i1c@2_
YMhN>J0:0=7VgY7RBH]eOPW\a`hcRYfCUSjS88=Egc3n\M566IkK:VjJ@bk@SH7_
6_2MoR[khWHYfTIH_NA^amf0BM05jb5il7H;X8I`4V]g^M]6_YmK5e^Ngb^@SH7_
64?MhR[khWjY>TIH_gT^2mf0BMe51b5iliN;cL]RIlWOhp0S?nB=]I[_b5<IZ5cB
S]Y<W0KIQeJBg4CQ^CFlHPk:Fh0?KJOMd7ACjV0XUcgFaYc7VOP8kfS>5TEahISQ
QR@:NdXMhONZbg3L^I`W:UITE;SUbWJ9PHGR`a`X=U^lV20dDf?YRfSoSjdOOASn
Q5YINI8PJ2NDbg3L^I;N:ZITE;SUbWJ9PH:?`M`X=U^WV20dDf^NRhUHIj@K_<p]
HWCj_T^NmdEjKD<MS<BVlPOUaFODJlVZNAmQdl;j22mVnqLb;@JA[QYYj=KQA1[k
[d2`^<BRCJ^hK0l5aC7<AW<SB:3a]97kHY51ZnA`f@>JLm<:TG:?O]E63jPGgO`=
663U2I8gL;jd_R1Oa>7hlP`TkC_9?<?3[\K`E[8Q7>OVEYLo=Z_`]QEZ0ocSE[`c
6m2e2\E8YJjd_R1Oa>C3l5`TkC_9?<?3[\CEEX8Q7>OmE^Lo=Z7n]J<T^b7Q0IpH
ZJofKS`f@cNk4<QTgjWR`9]H6I]hA7lQAAO_AKb=eOC1MSUV^GiBdK]ANG[^0D<d
QCNdYRSn>J_8?`UPNcL_7T7A42FnT>]ph2ILXcWa6IVDF_IB`H2K5nT3cCA0A<Ei
<E@D6BHn=M9ee0ghga]>71FQ[2U^6kTbLg^2lKM7Z\nVk4^eJX`L6_i=aHS7=iEk
Al@@5lZVoe<2R2JmjV[<kG7H8=kDVO5Th>7374g]ZWbhW4RTJ3`d\_igNR]9=iEk
Al@@alZHoe<2RNJRjV[<LX7B8=kDVJ50h>73m6g;EhEc[\LHqVnSIDO2jOn>A6V\
Fjf9;8dHISWnglRj<S;?cJ>L_LbSg[=NOHY`<VJikIPK>eKGKK[Uaj6[J4JAWUo^
S>@Xf0ijYeM7C^2V5jD?YEgHUn:J>1j[f1O9kli139LAAfDHYVIaWn[024U_VA`Q
m>BXlUij<<G>=^2V5jD?YdgHon:J>1^[f1O9k3C1J9LAAfDHYVIaW;V0knZ?TY4P
7q6:A=iBgjjYaLo0SAW:j^mnPDXLY;]<\DSSm;_oVcm?^m[T^9H<X9=SQec[DXTZ
:P36QLX^8Z?:HngiH]\94S3kU0]UR1\5]J4XmFG_1Wc6F8]g1LNY3DW?fn;3jH75
MO6g_6f9Pn?BldRPYU\j4[PkUCAKU_\<]74XmFB_1Wc6F8]g1LNY3DYafJ;3jH75
MO6g_6?1PfU@Ke5B8VqkFCnGMFNZd78Z0cbg3:=^RKiF;<Gk94:LMVk>Tol^HG0O
2AAhYBRq5BP\><KdI]geDdBg0FnV1H_hZgQ]U`5m^XN0egPo[X27eSA1<Q^mS9Xb
hX>>eD5\I<98W9hdnlg;QEK65`lJJn19BVK:;hJ@<EN`Raf9MD`JQNN0@^aA`e0f
lXQi]<;X5GHX=<fYn90UVAlA5ale4n1XHU]G;iJC<EN`[afZMD`JQ4N0@^aAlG0E
lXQi]<;X5GHXglfh2?mA;;nlp?j;LaEf=ecn5fh^G^BO7?GG8_9OQZZ6dQjDk^U0
R\lBDmZMK[U0Va[2LE8igU6=`?aPo<:L:<Ho:UJK54lRN2\C\aPM?kR2O?ADSZ_G
PRHBoEnISh8N9SjPQm:nCUkU0?m7T[kCH<CXGU[hG4ZRk4\C\8_DEkR2O?ADS?_G
QRHBoEnISh8N9M;PGm:nCU4U0?m7T1hCeRkdkc2@[qhJ4YXZja6ccDa=8^V1`:0K
S`bRC6Vm9F`9Xa?K2=Z2al\hb^Web>6M>`61U`:j?8gTSC2mL^_cdCYV;6<aamaX
_=[GCHfW[mVdXLQ;SVIRdb_UQ]fGOfYT8gUaNB1oRDhV:4lMK0_U2DYKM?<bam:X
_=lQX^fB[<VdXLg;SVIRdb_UQ]fGOfGA8_UaNB1gRXhV:44EK0HJ`\7enWq6Y5mV
<UoSS3_CWFEKWSn04POgK5@FWMZ[fMoYHQ9K]S^nSD=PLa=mPhI:oaAbTe[J?Ng]
oR?khA?dOGI0I_:hN6Kf?7FE2>laQMPfk=42g6860VA8j9nk<5e@:4jja_=6Ja`V
]Eek^hQj1WX0f_lVN6KSEKWE_>WaQMPEk=k2g686DVA8j9n[=56@:4jj1_=6Ja`7
oE[]6Al3T4Np80]?jTW@XS<eL:fQj5Z@@UQHiTSS5h^Q2_`;D<HUaoUgG2FCBA@X
ML8kkFbIXi]?_HE4faSSJk9YkdHe?:BAPVZZN=mRb@5XWm`Yk?l59I0d\nKYJcG4
e3a\Whd[Zao`87AXn[JEJhnWb=P>?]BehVZZTKc8b@5XWm`Yn?l59I0d\nKYJcG4
N2aPWhd[Zao`87AXYnJBF`jI7\=2qT?iGmoL5NOa4RN\4A;<gR;Wn[FYoXl]O4RI
oS8lC[l>`CXEe2KfY`?f]DUREDIT8UC?jU1gMh@@o:4lLMYV8a`1AKX6PdIZUd^I
7BbLATobBLAk]><c?=QaH@00mYJ]PT:L9BSPOhJKQ`Y5TMLVak`1BPaImdIZUd^I
7>bL`TobBLAk]><c?8OaN@00mYJ]PT:L9h>P@S=NGmmb\qD?O7Dd`S\SC?S[;j1V
iOA4gY0=8PA3AA6\HHHGmJG;7T=QWCN9bmO^QFS_Vk>`_P8aG<3UNoY8fJdDhH]5
d7ND:G1^lNbHXCjcHlekKEOjl05[iC^6Anj<bMh8d`Ll1GD8kaMh?BYfonb96Q]8
d7TD:GFnLZbDX;jcHlkkK7Ojl05oia^6An54b3h8d`Lh1gD8kaT0?6PSca4nPkqK
hDNN5Fb:UnLT>6@_j:ROHJTEOMOInG<oHUk<gl`XK==Y`QiHBM1Mkc^MMe;kfKhG
jO6P9<2fJXlOOL_NB@T10OVf;1H2cHYhLUgcX]7H?ja;4mmS\_3WQ<[IPk5Y=F?K
nnRgAOTf3hfIlK]NH@9\0O\aYA52OHPhLUgeX]PH?ja;4mmS\_3Z2<IIPk5Y@FiK
nnRNWO6U[jEYlQjpDH[BRF@\e_lH;7XEX^>7ofGHa30]dJ>j43NQKon9\G\GGXFZ
`Xj@GH;fnFD>U0Jo55<gd\OR?f_00Q47=hOQRD\afmEmc0NX;NNo5\7<SZSR1o<E
Xd37iYFRYa5BU3@CDjef4OkB?g:RHCkk=8OQ_D\aDXLGc0NX;NNo1\7jSZSR1o<E
Xd37:=F@Ya5BUR@gDjef?2k5?G`YZA]mpUO\B1Sg5>DRDPVnDpj34Jk[l:LH67I?
D>HCZT[B9h302YK<<2R=QY\n73W`Zi0VT6k9BA\lE2NaKQ6;oGFP73m\APiLZUVY
6?I0JQECFZbSFR4>LE_YQ]\\SInL]jI^;agn2\_Uad;56RKXRkjNLOVe7;iiANkQ
RTIMJ<4CF:>Foa41L[_YQ]F\SKnL]jI:;7gn2\5maf;56RKXRkjNLOF<7G=4?W8j
EEq:F\:M[OUC@dn>o<5^fnmXiiEG8LRgncHADHZ2o6_LFHMR9m<oe7K89d04@VZ8
C=]RJjNhY0oO1mV][683k?23LI8jbPNS>Z]gVH8lOS`jCQGI0F;_<>NWF><cQEJT
@ol:jPB<jgIO^be@k^O3D?2^LILiJ]LSEZhgVH8ROSajCQGI0F;_<>NGo>_cQEJT
@ol:jPBlPgUBnBQ]?ijq7fMeW@\R:n>aTDAm:^Ini5UWD;M7L_9M`P1Wo4Da2]`O
>?Fd0nZokGMdi]kU8VAGLco:flQW0]^diR1\0?PBnAc8\Nd^X<j@L511I_d0m94>
S;@EmHClg@ZQ:::?Ua777BNB9]g90dGiYBFO0PPBDAcW_7m3X<j@L511]_d0m94>
S[@?mHClXGZ::::?Ua777BNBCHgKEFFhG9jNpj]eDh@2STm@d=_MMnR3X_OdY4fA
9VNQXbhc@enFPccTkjFh<4Z8joBQhn>27o1:FT5oREecBE>7CSEGJ?M5C>EHjd?U
k9S;gB^cNJB@mZ?H0aIjZl@[nAPTLBZeI:DSDjTF?gHCWEPh4Zb`@?M5QZEHjHo;
A9S;gB^cNgB@1Z?H0aljZl@[nL>TeBZeI:fSGjTF?n>Cl1ee6g\LTq:94H80?KX8
Zbc?0JhM>l@0l2NRV>a`QoLFMWf]g4ej8@9P9<DQ4PAMdTmiCIZ7;Vcn5IO=K437
Q=Q^6LAbbdRa9E4d5Y9lXRpLj3@\X:7;]W?mKLNQe6k]jLAhjWg41>SMifRB\F^k
_RH0nmjWmAB\jGO^c^N^2p8Bk`FmQaK=S5T\j4OLDOn4bcJBYMH8X4T\^Y>:d_D8
lk:=`GgiJ7UJd<b=cmiV@LCUQW=1hR;Kj[WdTUeH^[_Mhi\T^]lJC5`o^I3<Ya^M
DR9gdGCUlRMJfYWa:72E_M8[[om4bZ;J^^e>e2ek^[<Phn6<nXlJC5`o^I\<Yd^M
DR9gdGCUlR;Jf[Wa:72__`8[[oO0bb<d2LJ]CDq0nT@;ZSgE[@=BV:HcB918EE?>
K2SiSi^dW3O;Xj]lM@D=0X:4>VD:gH`D9FU6em\2VlUWjdLYc;L7jinf<c2d2Q\8
imR;Al@PO3]l`DjU:ZnJQ7PCTJ3a;K__CiAHbAj0SGh_cDNY]FLgVemf9c2G;Q[@
2J\;Al@PO3]=`DkU:ZnJQ7PCTJ3Q;K:_CiAHbAj0SGhC:D`J5P\F6A@pD7>\Nc<\
SJHRH4eXeX0\1G<9]@BTBLU1c_lAZaZd3VZ`K`iSMi\01TNT:3F4?C@__h_LFf6J
QHeUE_VGO:1UIe\ZIM9DLgaQS;l:D:QWhP=\M<75_^?:;7`@fc[6L6KAD9NA0\3V
Q<kZhHUmOB1Ui]\6]`_jLFaAS;l:^:QfhP=\MP7N_^?:]7`@fc[6L6KAD9NA<o3?
KcESM?UgqEDmE>\V>AT4MOTNU?fRL4h>^Hm`2`S1Y5E?TAH\8kd_DaeTk47WPMIb
`96mNdP8YNYgUk6CgSS1cDMH05_e^]7jH]NbeOCES1N?j]ACAPE9C]7=K[57SPR^
;Il<1G^XQEJWPo8Y9S6e;YNZ[5@e^B6jn76NaO6EN1N?jOACYPE9C]a=N[57SCR^
cIl<1G^XQEJWP12Yd5[1kAYUGqHV9M_[W>Sgg@V:fQkRa^GM;2i1Ih1T^P66[E`X
hk^bQ[8DoRj4kXZcddL9fbVi;GADW2WUU[eiT\@45RUHg9[M\D6CFO1=iN94[EO0
1W@Q\87AKI:H\1RZSeIcm?XjORH]_lUbP6eEYOUHeTUOg9Kl\8VhkW1=iN94[Ee0
1W@Q\87AKI:H\1;ZS5Icm?X]ORH]_la]PHJQU4JAVLqcQZAOIlPP;^Jne\WjbJG7
oMmbj<g8GK]@`e1bN5lCQ<LJTWl_IfYl<Obb8lM?[ga4:TJ[2A8451JF=K_8kfhn
:eIYEjl[:^X;<ea4ljEV]37K>bogank;od27fHiTGeLcD3]QTi64DCbA]<n8KfhL
<eBf0Bj[>^9;<ea@ljhV]37K^bZgankXodQ7fHiT^eXcD3]FSi`QhXbOUngpeN2S
=?MRF>A>Xd<K46V?T_iYZ@Xf<CfZ5c`_LI3H`G\bN?<<4^clFRZ4[FK``=Oc3HM4
@hq`c7^;[^b9DhWG;:6C47jKi664]IO[EThPS6W5RST53niOFkZ963E4fZ>ncK0W
=kmX79KEZ?=h4;Wmgl`2:bB2Za2VTTmEo=6@a6[gI2l_lCHBh0N4mamdgKS\AdBf
:KK`i\WIhJ:hH_D>;4]2kbQU:aao7ekEZ=T@a6[ZI2P_lCHBf0N4mam6gKT\AdBf
aKZ`i\Wb`JkG4c`Te\3pDaZfEgT83;UhJ:n[PeB8n9Yif;JcLk>3<i1f1\SKTAoT
0SDBSd@cS<VfA5:MT\>26WN9`cC7mZ;_Y?0@@FX<cef5Po^la8IiSA1aD]Dk_Y`d
l`3SnNP?Yik8^]bg3IfLDi;[b6mFmKjoeGam@oXYY5fRAFiEa8IiSA1aC]DE_Y`d
l`3SnNP?2ikc^]bg3IfLDi;[;kmDP8\FSlo4q1QkF<IgBH1FVa5;FdkC][mUQ]bJ
Eo4R[XTUc3ib5W80FfJ;KQV4<X^GdYOG`@U\1YYLL\fHf9\^UGgE?jMfj6?b8CoH
acjdGUXUPETckiTeC;[jm:^SUBd2e9DYWnE[S1R=eF=MW9X_UOXK1j2fM3=bGPLQ
kcjdGUXUPeTc`iTeC;[jm:^SUid2U9DYWnE[S1R=emoMJbj>k3YPlpm;\OHRXc0d
R9b?YQJAL8Z3Yd5UY?U78C^ZWV;1\Dga9MjWjESAQ[7dL1LVT]H25:7LP8K50R9R
SK@>]cl^M?9fWi@V1mfmC1M2WknCai:7>QgM:Q\Cd\L9S77^^cZZ1om8lQd9Lh9O
YKe3><lVM;mVWSO@>>fbCVM2WkHCaG:7>QgC:Q\Cd\G9S=7^^cZ21Gm8lQ1gLan:
m3c:3_pcc<PY5DPRCdQBR`h=iT>Wo;NHhSdVE6_@oiOgQHYm]N`V\enCbG80f3<k
47UJ>Q_[>0BOcS299UBoHKo<<SXfMoPVC0GFF@?Qhim=Sl?nGTS9eEk]=V>L>74R
FjMfNEJcPAVoL=f9JNJfjJT<VSlUXoU@hb?F8@eQhim7SlKnGTS9NEk]=V>_>7>R
FjMfNE]cPAVDY=Fb3XJSfPgpk5ZQ1iCK6i;2=W;@K3UJ2Am@g2Zn5Z`h=hHK:MiE
^NI@F6G6Xn=nVV[em<Jm@R9nWVDG@8eLHF2`;@1Z9:`kda8N27iC@P@^>HH44fK7
S0DD[8c:GmeneG;C=\[=>beRk@S\1e4eHg3MnS569\``Jc8BS>Rg@P@^>HH4hfKC
S0DD[8c:GmenGG;7=\[=>neVk@S\ne4?0HnY8hRZq<38@MYXCOngOLn03aFn\G2<
pA<=;hmRM6jR?G72NEd?h6IWT6=^D_C3YIB2jlk6QTDnZ<7GIL8DAH>7LoX2nNBd
OPZ__W6BSRKjB8OjSL6jm:1=_6M7n][QW@O2miS7QJJUQU55K\^6:7cjgdMl<9h`
NAjA@S_a@RenC\CGaLJjm5_=a@_LN]`Q6@O2m`S7YJJUQUf5Z\^6:>cjgdMl<9h`
NAjA@>Ma@g3>Xm;b\p0J<jWdTl59o]?NIdB@0]1\]`NOZY@9;_\`;]FhK7c6:9En
IOlCWnc]j1QP]W7l;Dg[a<^[UEKFST=3BiF^6OZET;]hGn:A\f6Y;l51Zja]DcK:
kLSinU7Na;0oXkS<]F0KSji:iAK<IT;UU7F`6CIhThZn]]:>\X6Y;l51ZBa]DcKb
kdSinURNaj0oXkS<]F0KSjLYi]KTVK4F[MplfoV3M:1I9<H62KM`Y<mnoOfcNMk0
l7MaQgmf^amQ^aRg3GWSAF`^e^35Gkl^J@I^1C5l<lX<gJHmcOIQI=KOVCo0dRoJ
V9DB;g;`\g=Jh6edW5VL[ZcI\k41A\ZEVc;ld4KW@7i<^0_NlPPQg=CdbCfGJGPJ
V9DB;g;W\g=Jh6edW5VL[ZcY\kD1A\ZEVc;ld4KCF7iOT3VZQklpCg4f83`oKQ5A
A>2k5DiBKMiqGDO\@RgdPX^g8_F1RoS4XQM0CI3PNG4e@KSG@UOcCUA>>c85Q?CH
0J5BE:Gdd[>D3Ra6:>KkOn66bdnUKXO1<X\j6<be_UZf41S\>8\P\S4X?@^=b<P5
\e9L3@E`dUWSGThAeN=VO4=0gTl;K0ONNF\A4hc`_UZf41S\^8\m\S4X?@^=b<P5
Fe9=3@E`dRWSGThA?^=FZ:WgZJm1p6e6nGGo`IR8UIPlSFB4T8a@500ZFT4j0f`L
FVVMPC6^:7=Qg]3ISkM02Rc>B[I3WVMkmUWVmYkPFINnOa[hmSdZ^=c54?QPHqnj
9nW]P4=PHYRYal7d<P]Y4^a[?UYA>D7[l:780:5]U1ncl2c0\c^ZQj71WBN?02_5
cSl8Dh<hEN_eMP[RgPKaAKeWYe5lbQ]6l>lSSEm8^4@S8P2KoXP:WM2<MF?dNjn]
F^24OC<NdfZ0Xo[_g0CaAbXfKZ5lbQ]6l>bSSEm8^4@S8P2KoX_:Wg2<MF?dNjn]
F^34OhbB:A=jGkqT67dOh3352Le61e6J:C6^Y;EGR<m9X^WD6m;;ZBlMV;PDj=NQ
17`4B5_JnSmD^Y9l?79[_8cFFGC?1jiKcTZZSV2XM?_23N7KAm7W]UDn`9Mj>C1`
F4KV?R^2eWk91ncTD:IGS_jFH`ECCkSK^TZDSVNaDC:28NeKAm72]Ugn`9MjACi`
F4KN?R;2eWk9ZnETD:IbS_\J:C9O6;4pSCj_lhG94jV9UGE`ME>T0NM_D9=XPYTH
U1^l4^`LXWPnFn:`=X]7^g>V5Q3^Q5YVXHjGFJV?]cYi:G@9a`SS77g93=f1_HoT
ch^[IckngE8UGaF5T5Gb[9Eo84o0EDR^Sm28;?Ud]HTo_1\KaZSSC7ghjQG8_1o6
ch^[`ck4gE8UG9FST5Gb49Em84o0E\RLSm28N?UAUR34E8=BpKnI1bVaEYT9nAlH
h>M<Dc2G_;ZPFgnEYhbBV]5W@;DgZSK2HhbQAmQYUmn8CBEZMF?IZUES<mIjY=le
1KEiNLdcc6HcEKDJD<>B[=j387?Dl;be@M_Y\<7A5D=a;d5]QKkE4KVMbm]BDWSa
DKkiNBdc_]k8QKDJD<>B[oj3=7?Dl;be@M_Y\V7AZD=a;dS]IKkE4iVM=1cL8fhP
3pJ>5:8W=QYGKZ:j;`8;EkVHb[dgWnJYS>UiI]PP;ie:7fJXIP6E0>gObg58;7?X
of[i6fBNP[`YibemD<em4A3gW\jPUZkRZ6eRIJaU>kcl]82KF4>F2Z6hoXO9Jg[3
9kJ^BBjc3:`0A2kNghe74lKgWe3>@Lk<ZSeRIJ;U>kcl]82XF0>F2ZkhojO9Jg[3
9kJ^BBdc3=62mk]K_5qC:RE>lP>IaT0kHe:SA>TZ`dbLkef<WcfcMMK]NFm3PEY[
K]Z1:CKAhRalj?27IB?86qJ\@O4b5l\m8CH6ha<[l==<JAGETo=L^5M1m0Zbn[1g
oa1GRHOhOdo^On<mk^8][_bAB?iS\FdUikg0Q`WXC=:b2iikbPll<kUgm<CHo6Tj
4MBAYng?HW]SE21_TemYDnJ;NgMGLgdB?@mIX_WgCh=b2im3hOlo<BUgm<YHo;Tj
4MBAY;g?HWoSE21_TemYDnJ;Ng4GL@0XJ43ER9pN_;:Hl>I]h<X2;J\C65`ElL_;
<nYl9kZo;=;fE55@Ba<AM4PG:N=laAYN45Go7HEeCCU^]\C1WOnG52bm:U5GSA?@
RUYm=oONH=5E@i\TRiaLo>a_i1oJWn1]db`WLloNR7V92<T1ogA]@oomgUX9SAbG
d?^m=oONH=5Y@iQTRiaLo>a_i1o1WnF]db`WLloNR7Vc2<GeKk9obYBpe6hbA:_^
Li@j44[fe@?l\h61Fl_@@HEX3h;4[55D[45N<FoK`1EhF9aFXLQaCKVbOmOP\BU_
cOFoDe8nNY^lh;k5EI`KX8?DoE;eBJaMQWMedfg8:gP\<d6dO=HV61g2ek^b4QMo
c0[7hTFbNF^KX;k4[l5VX8?DoE;e1JaMQWMedfg8:gP\Md6=O=HV60g:ek^bYQMm
SfNjc6eepL=mi5I5ed><4k]8[JQ1M5[\FcD^h<jVll97QlHcn`lUQHoLCPU^[7VO
LjRiYE<kPL1L>?TSNcEZHg4W9J8@7FNfnN=hbZ31Acj7]VX5TgNUg6I0PiFE^Uij
mFLDof]kELJ;DPHaJc`o[0NbKJS@k;NfV4lQ`Z31Acj7]gX5BgNUg6I0PiFE^Xij
8FLDof2k8LJ;DIHa1WBc9]IUCq`iUoU@j7WhP^\RXF5cEWZ^GnH<jCL8JNQjW:h?
TlY\^?]TbUPdUel\=LaDC0enTV9RO]9a_gI8A:20El@8B2LQEaHVHPKBh]PPWa6J
7@AI9?i5hK>7FMDG0C=Y[UbWL2`gJNmnSPIo\fa[5P@gB2kQE^Ya7bKBh]PPWaZJ
7dAI9?i5hK>7FM4G0C=Y[UbWL2`gJN;nSPcEJa4KEXqbBFZc6;<kj92ERJQa]cYH
96nn1DYXN;KZ:@>cVNmQSHl8I[dMG5IWfSUdheQL[__J=gbP`g17[_XeXihHLaK8
:9cK0CZXe]l:i@Z2\\;:QF=TWUjTa=`=ob4MBR?6IMCb<14OGC`7;L[MLB?Heaik
:9aBPUlX7]f:i@Zh\\I:QF=TOUgTa=`HobhMBR?6IMCb<14`GC11DZaTh5<p\j<f
<dO`>YQ@??k[^hO\XgiHhba[hai`FI1L=]05DAEGRdM@[YVQJDe@X`33o5ge>A6:
I8BUU4GNI@J8lhi;:c1DDl\D5oIYYU1LdN8]ZhSSZG_WHcVXi0QJc4lgm3=b\5md
_2]TUV2bR@LCl]i`dc1:UCZH5<I1YU1L^N8AZhSSZ__lHcVXF0Q8c4lgm3=b\5md
A2]Q<GUMDYI:pMeFKkOm`JY_5GED]eZ8p3AQef^f6KmB:j;=U<Seb@1?Hfo@D?JM
S6]08^jUHDBB:8Qgc]>:`\P6AT@R>bJmi]5a^\N18`BICBkZR]5gkU[o<Dfg@QLO
CK\0IMG>Y@2S9T?CVkJ@i43UBV3A8R_iU3@ge:?4K`SnEe5^P]0gko[oNVG_=QLO
CK\0I=G>X@2S9T?CVkJ@iO3U8V3A8R<i33@geS?4K5=iNG^_XpLn_M?^KY3XmI`^
WYAOgDDFe?dRHVEZmIcROEaodchOMZ5?8e=3kJn:j11_]dSf@EE:3LLF3gnHS1WR
6U?W>R^=9R2IZia@KQ_@OJCdeUi<W@5CmK5BcQjSk0L[j^k`;=L3;LdiJ2nj::iI
UF?A>]D=95jD9?a=K\_@OJGde;i<W@5nmJ5BcQ_SkdL[j^kf;@L3;LViJ4CCmb1U
CkpghgiR<dH7gTM8QBkNK4JUn\E>6<LL:2YHJ6cFQRA2W\6FT0Ug`aVKZZi`Q]N0
GCRcc5Fmkni8ZLR50\M9::>cJh__;KWa3BB4m6WIGFSHCLio\Jeh_Qbfc0:TTn:]
i0hgCHBDXbd8VFR=f>A9Y:ahJh5C8]>aFB>4m6WLGFDHCLiojJ9h_Qb8c03TTn:]
F0PgCHB4Xbg9ff0]2LcqVYoHflc=oDJfmh7878\5=1kml6n;<o;6n^5\]]j=SJ6L
2^mUM>>cH>@UdaJGOL:36To143GB[b_Slh4OH1X>1Y8X;WZVRc]CEf5MYjmL;jAQ
^eM:W`]3fJMOYMQHCK9IVbXbH^Kg[@Nk;^[<H\X>nY8dVg\2Rc]CEf5MljmE;jAQ
^eM:W`]3\JMEYMQHCK9IVbXb>^KO76PFjZ8mp=d4NU=;agc?Idi3;RVOQXVABbk`
VV:XVVdm05Y>J8=GQ]DLXUD?mkdE197h=moJ0CbZhF@kdKh:L=UbUGTNaXU=`h=I
\nA]dp`9IC6^qoNm@KHL$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DBFRBN(Q, QB, D, CKB, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CKB, RB;
   supply1 vcc;

   wire d_CKB, d_D;
   wire d_RB;

//Function Block
`protected
kQEPRSQ:5DT^<F1MD^d6U7daB5k2U=p`jePePg9=N=TLD6b[=V8L?BcJNlSnQ8[O
k?AUGiDYY3ni2Tc:8_q]>hU>fUOY^9I=]TSSHhiTe[T?[6W1TH^UYWWpL2PIAPqk
_T<aZ<2P47=moGK]T]420bZC>p>S4k_J[NPKIk;NE;]HIVQ9U_ZTVp]W[oGM\;;B
fHiYL?mWA50YU1RYgVL@@75Pe02jhU7bR2p]7d2`4aQO>eETdAjG4h7C9aQ@O7HL
5hIFVSc9h]e9MAh4J2jeDL@SYALZ3ZYnnm5mde]73hFE9;:qS4i`6_3kOIcF3N1n
6DHY<<hm?T5JF4gVpE7noUX2pTe6RDCqZ8eg=EUhKNRP@Af;[RSRB;YZ1OakJjG9
H2hh83i3K^A?5:aJN_kDEZD5HX2GgIY;T2LTIg7H@a`0fh;eC[^QR@AK`nNGlA<Z
TkKLoIkcBYV1VIqALgYo\3mZ=b[1hN`ej:T1TUM?ojTLFg98Go[;iT?cYJIT60CY
N\?CFeVo0T9C=LNS6mB3=SGm1F0\ma:>;TlCYX9YA<go^cHE^Z]a_6H?_b^Pm9pm
BM7:Lk;Fc`=3[lE^EOfE7XGWWSF;3C__3S3YFOPeZ_CV0bSm2:KW6im>h>WNnm\m
FMG:=8ne?JmUe>d\:cT8m9^XkA>ACnGm4fFp_]kPljo0A9He<TkB3W43;IKoMYFK
MMT^Xl[@LWe=C5=mCJdff5XnA\m5G6pZMNaV`jgI?T=^V]7o6m=ZJ[D=N>eO8HGJ
3R0KlPbXiWiWlo21j5nQIO:e6=06]g`nW_jN0kUDKB0LViNOKgn5oi\j=OhSB5_e
8ICGhFkKDp:JN>4Mq<SGG=]1QD?\]48g`GJ\no4;KKXA7APEA^n:_ENpgV`LYWLC
URjZn3NcfFOEf1Z]`[eBCFSDO6ECpicg=D@NHaWa:f\N2j6nA3hiUA`^PPT3m6El
WmR^mKU``CdgG1=g@aa[n<YJkG_W>g``_MLTfi;lK`j0a7E969[M^`9UDoT3g`6V
k^bDWI:J9=X8lR]iJ`1=Q@__A8H9h<So6O^_qG9f8UH35hhlFkcP6L9;lJ_dhUZ^
:iQQJ?Lnl2=@1OTTB[1l^Fk_5c^RNqWnaleNgNP;Oj]f4V:e?6eFn;ALVcH?]Ki6
`\F\84ofMLILWgCG6L4Fdi66Ym3M60W3Blb;N@4kbgMPe<jE457T^7Z8>^U:3eZW
O\?`l=fF5NDoK:7lM0RdhP;^eil7]SaTV0L5VY`GJqJ9ZfdApRD63>2V=BoYhb3<
QB]T4LLIJ<9D5jhVGRB<K?=SU;XDq<<E@G94ieGlB:M2>m`Fno[Q2PNJ:[<bU6n9
=W3kjf<5^pHhVNcb98FV7KK:e[<0LTnl;eX;C42Rg_DDO3@5Q4A`b280^\9VmUMD
bK<eBl9;_GlI@XYSaB89o[\RGlT\E1EdZUV1M`TcD19_cF2kR0@oO3\`McW6OD1f
6M^WgQLhT`o:^7e2pV>7eKPmLTJ_JkeLUZK<CR5W:_g<P6cI_3iCg0]DRW>p6MX@
GWp6mT5mO:EcRCI1`7U56>a::0Z@3ADIZTo^m[PokqiAD?BRme]3KEnSX_<j]5TT
Wnj^M]EhG62o6M^Iql:`<DRhcXmBB?nkESM4eAlN9Sof2cGDhib:8ObpJ_PlD?g\
ii6MBl7eLbnBfXGf5jf<^UOTc;YR[adRJHV@8:N860[AS>0m;8FL@7ID<iiLE[<9
<7pDJmTM=j?`FHk:jFGNCQo?[;:lo;bZ\=^TSUf1<:iZeTj=AfBmHU28SOl?^@h_
dTYCI9Phf0p29Hf4G6\IhFjSP:c]U?^6YUNcgFoOAXkS9PH6PV8M8\P\C1iV\IeK
DVOohG:^3_<MdHZGOn_Pooq`;;iMPS$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DBFRSBN(Q, QB, D, CKB, RB, SB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CKB, RB, SB;

   wire d_CKB, d_D;
   wire d_RB, d_SB;

//Function Block
`protected
=@2S>SQ:5DT^<\cM]^WF8kRll7h`G]dV<dJIIdP54[^pc:nhH?iB>@LnCQjZk^@[
F1E8>^Wgi42P\ZkV[O]HW^CKd[F<RA2Gi:91C;6pd3l4AOD4TGOEVI@bGRB:fmLV
W0qW6PU7?qBWF^PffmCj0L7F89Vjf`?3OG9:qTjmmFceZWc:fA[l5cGKW3i`1J5]
lp45?l^4h>T<Gl3:f>acRJCKD8WO\EXT1]hY<cg7:LdK]\e?YAX_KGbW_0YU[b:h
fih8;EW_X8_mWMjGpQTm7ii@Z[b<>``O434KDBL:VR4AV6GDTl8ojW5fHP9fii0g
V?5R7HfUYDiheEJp8Gb;oHM7GTO;OLXVZBSVoo3oM6jYI7:ifK2Y`YO7DckBKnPj
p6WZ2@Qj7l>B2;@d2?1IPOO>n]f9`kgmjee;j0`>pYn\C2FMYPZ[WfHA74jhHU5^
D8FN3>HR4B6jp0570<U<C0>5>UXLQUJW=iZ7TAlR`8[\^pNKYTmMPi6oJENQDO2S
=R6L9^hL3RomQ3`Taf5CbFk?fNT<qX8^[ID:Cn9bbHN3P2MjY^n:Xm5C@3Z5nNNk
_b55I]OK;pUMeI2DShJb`aAh=FPb1@\5oeBYe4]Wb2W@1X@]AgXO^1T_e6=XTNQ^
4hqaL0DBBB_i4DnkojioHGmNm6JXDPkgBl@=oWmWgId@5hcj\QC0nJYk3Y7K3OYd
8T5eDTh86JhgT^2ID>gDCg1JJGfGIl2>SZboZ1g]hIcfN3qa\^?0E0qW74ImKlJh
Y`[2]JdCVK`4afGe^jcICoX9>Q>^ie8@L8=XEfTC84XdMkK6gO=p^O^:Y8q]CRa2
k>NA`k9[i9oG^PG@24IRASXHO8Q1\<FQ_8Q:8MQ_IeWGUQVlm<h^kNcWoZ<`P4T@
hX[>bYUDWYg:FfQ7[R[E\f<<?6X>I>]fS7XV=l@:?p5ca`0nIEPJV=<A>M@ShVR9
4clI@]ajAUUZ;Cnm8`LEO=\kY1M0Vi\ojdQk>oMCB1H9>ZVaVCK=\S2ldV[CgB3Y
Wb`i@jn1nADgGT@jYGWNbnP3_q7FDA:o_nhdb<Q73L@B7RA>IN_<FZaQ0L;Bk5Af
Nffc2pE_5gN\oVbSb^j9PU97Q<d=\UIdEHSm\a?0QGWcY;Djf_P[QSCck<nS2:[@
UMN:<lEl5BN6InTlh<L^S7;<e98n^SC7[j]TEA6Wb[p1OBicTPg31\^Z^fd\D67A
^l[Ug@WHi]<Fc6G3@HFmTl>1^3K@ATG8<@F=NWnSJBQH7cQo`OYo426Y^?LB7M^0
oMg2I0JVhn_^eF<nYGAbepCekSc7cPCWf3:06IKMhadW0`08;V@o_XL[YT3Bkk:j
TkMlOcXafB;lkBe4WCXZI1iaF=[QdA1Hi0>0kcRo^l?X]OgRnlMD2b6`6jPDZBqF
:LmOMnS5cYS3<5c5eWD047LR<F1C5Kh^abdD`Wb_belCb3;HUc_NJG:<MdVOW0EF
HLfOXC;cTBo3MUbQ\XF76ci5h9HUZmLhgnd^op>f[0^@p6:L^7>O:eXNQn\lEJZT
bX]YJiCgoc]<7g8<i\2pPDZ4QH@HF[4P[=DJ<:Jg[f9aSE6P@VgA5afAp5CiOh8V
?4mQb`AVU04g3oF[^<BTN?GEoW;g]mN]<GL5c=CfcKPAFT\0hUK]nFGPLFTH=ZP`
Ag1lhXJH@_ZcOJI]GWDYNaGEk`bD<L_MK:Y;iCoJlGW8O5?C[]_OYoQnNNfk3=?m
j[3fQOk1I3WEqhU9l;P`ED8n_5HPB:[=l=_eKfb4Cb4pOle02aU>`cJ2SCeUAbKM
;Rk2d4ML?d=Z6U5f1Dlkca^QYU]_mokL_O>cUTnGENSSOBk[kMcUY=[?`3AJnFN^
SamX9\jHkn\8\e4_\gcQ]R;@aXC9d3SWAm3XGUh\ZY888::gU?9KF9:co<g4[jc=
[6^p89^mYJqRbZF9]i6P=LMl]g:fbLBFR8b>k:iO5Jc^`?YAWlF]iTpQ[F=Y<H\;
Q1`VnfK4:MQ6OX2UK8IBd8NgZ\iRl2RUfQLp[aV@<Lg[h;5A=I9C>cb^6SLK93``
1X0[ecl5jn;;ZRTqfGKf=D[Yk\5E9E:e1F3FTUH@<;ldWRBc8L3mUhjQd01q>1C]
\83PUaRf@F5>`EGiZO6YM4^gfQV@h<>AW^<^YEMhlTeeQ:2ka?E=JmiF=eJ5>@eS
UjUCaTe]MYV4S[0Z08JS6695HnAQkH_52La2];dfEa\^b]6S_>1KO`SAP]45U2kh
3=BQ@>qD<02?aY0eCk<5eh]cXIT2CV8aodRLRo8l1e:XfCLZO:mA_fG1A:cK=oSi
7K<TI]WJ7GC>>418Z<N_GaZkhJ?WPJ96QoeYhX5Zb[RhG>@_O:8J;GgmoWOISOfI
`P^JF_A_8KP1Q<q\Zi6b?qlFBfA]_FXXTSbgWWDlEk>DGWRA2`lYJSqF<TjXH[So
YNdaOfl\YS9f5PJ8AJ?oVILc7BW:3qg\F:Q8i]d;EHeMLhPae7f`4^^5D2m:O>[7
gXBjq5P6fOhD]m?N0ZBjkO3NJKmF:A6OAGSml>?T<XbQqP@g4@:I;ODWD4Jc;g?[
C6djk6Fm==R5ZSA5cLc2qkh_eT5A^R=mLg`ho3eIY9k1?<f@e8EH8Q_Bj`kIM2\N
flJGGX=8cH_\DeT<Fek\EOjPL3Q>YO9p1S6c7G7kGcH<NTU]M]6S7m3efCIPXMF=
i9pXY45i6dR7@L2XTA5JhaW\RS3I=mcCIeY@?CURN>DEVf=140d1V]6oRJk=D_lN
TffP>>VZN^JYVp46HWdfVaRB5F:lel^W@Km6A5d4HQlm5i^d[A?dYW9444Z@iag5
<_k;eP93mG?16U[im7UfZ5E7bqG0Pf4iFe`n4LgK9IUFJI=mJ>hO2ES9necVIDR[
K<\F3?8]hQ<>8>fM;Q45=6?ko@oW;EbYdU2oDq0f3_ni8$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DBHRBN(Q, QB, D, CKB, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CKB, RB;

   wire d_CKB, d_D;
   wire d_RB;

//Function Block
`protected
E^SZeSQH5DT^<okD\m[TdQ?1k_I]?KZ`^0fFClPNlQj^A=GeWe<f44FIp_>YOZfO
5\;O==a\NC<FEmJ1BY2^eij_6k7e0QG84B`6Oh<X?eh9cl^SFcc`=qViU^FZPVWR
UP1?[kR5A2A]B;97XnS5oTEO@[g;cp4aTNj`q@i_S2^^k:E4@B<jZP1`mhl\h3lp
g]?TfOC3F@WU84Lfhmo8GL39AAJqZMb6TRU6a`2RUVPNiGDdXMBGmn<`:^65RYp:
94Hl@4GPGC^J7>352R7eUR9S@Ig9oU]mc`\>`<91`jHd9NhnYjQmFLQ]bc6?ZMNf
Jap2KJ7fIZND<Z0W4Qoc4=T6eM@_JUeLQh0pL4>>faVp^SSiH`qH6E<iI2j8[a_h
BZF\K4D[6OgSTY[KD]gL\bmLnU;LV2Qg@g4j1I^=6GDe7R>`2ATI8Rjf4fNo=N2f
e9`_93__l[FIe__Ji=NC]=388D6nRg9bkpBe]AeSl6PGFb4oj:MV`YI>f@79WJ@;
K94W;DcS[S`<Q3AdoYa=[HQj9@6l81ToG1K>6i:D]5=mRnFJ<:<bn50\S4Qj]N;F
QgCUZC77Z:lTK]BL?qPMR__hlQnKL?H<YYUPWYW@T^7[GUZWTe24M2=lc\`nfOcN
3k;b2lNFJ@nR5;@hJj^OSP99bS1`5^F3n_lM2@KaqVjW[09[?9<P`i<nJ]_8kf<k
506@jIAJo]T;9V<b@NIkDjFd>\YFndlL2`ANYm_g6;9W^Q;H]jASDeLIENZ@G@BO
OIX3qL1GKOlZ`1U>;=cZ1N?02MH;4:2?g<<WgDJY<V_\G6fmV0R5I50kPP3J9ADZ
A7H@Q4o8Z7Q9YfTl1ied7VEH[K3Rpgj33JDiR6=dgR<<p>8KC`l33bPeCQMeXV^h
4aH=42=lN1ZTM[YiWS:8o@dQ2Z[OOf@lWXd?njAA7d^PMQJP^n1n;mBfR:i:S>MJ
m5E^9\RZ>qoUCm[=pc?H\3_NCGI4RH9A?`HX^m9;0\S4P<\a[Hhm6YfSp_eU6XTV
ZbLeHn6;;WRQ<aJl35:g3e@cKFlZVGJqnlZJh_G>1Z\d[UYE_eL2j]l4W]4YEP8]
\oNDgoZmdkFX]I5LD^mGNOZk=B@BN7;mnoeLIOPnSa[@FIa6eTYQ=`ZoTf^VdCEA
]RYNMjY8PNUG<NjZ`<EVLf1c08cCFMlW?EUcAF`AOB`qYLfVF6`D\Y7PcjThEYBX
4`?6Ze[3jA<k5A81Z[IFbjeHQNqnAmFo5>40fcB]mL2K3gZEjbM4hXoeGoP\hUja
nDNhMVC@GVCXj8M02iL9c2SU<7Nn\5D<5b`\ki[`nH[l3bLXl`BhKRLID>f@o2kP
eIQ6d?:WnfT4l^UZ@m2<VI@3\G;?<bhE9`;j1mpjh4UcSpafE=lbc:IXmhco\8^0
R`<KLbJ<oPRAD0KkLM65b4ajMeq\;NSYZ0=;0Q_eU^Q;L[\k:H<1Nfl5[DHVi<kV
I1o71IeqCRcm9f0OKa[?Y8PJf:cl:ChEa8bD8A;]=S;WPTCKkI<JTb497_j7JEIG
\Gf5<FIBlfbQTdcEo;V7UPWYIMBKL2POAYfo2=F>oYoj_7MV:f\=`\\SJ[Po@MgX
BD;ZqTH?>h=p_1IM<KZWm`LEj5V:EUSJP[`m@aUE`0TlF;`ClJ=q9m34bRbXD3P:
EC4a?;dQTRNS4_lSZDQZS5P=RlpRacPS3m9P>ZW6j[Y^O\Q3@l^5:H5WOk714kjQ
m^WV`BN9o6:^LT^BSg_2IMK?TB]L1qk\`J\3:f3Efih0@g;NbCF[`>iL40o1;Nhb
S1<ai\`90<<I359FIEUmoRmID3FC0j1LLC[Rj0hO7p6R]eV?1_BNeY=<fS<fcUY1
bTjEVIZkPUPVaHj@TEOE2nm36EJQoeVK:332ONd=GB^d?2infZEJq]i]9Nc@$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DBHRBS(Q, QB, D, CKB, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CKB, RB;

   wire d_CKB, d_D;
   wire d_RB;

//Function Block
`protected
U;dKbSQd5DT^<cbDdX7LVg\1Eb=nQT=ZdN@QBoS=PgY56IOgYbkF;PL[N<38X<E6
^ah^BApJGiEQOlZCl2MV^BF9afnXJc[CJIP6>]2a36lYRpole8EC95`VGcS0kHSG
gH32h12LS0dN<KD55GWl6U78>TW[LCL6WRfM\`AWJLmVJc26qc:0=fGqkjX;5m16
GKM2:8AjYmUdnBO=C8pTg?9ZKBi:bD>E2D92RUTb6jPTlVp<P=ed2@e^<ZKe^VMC
NFMQ702Yig<UZZ<0EIZ^3h9nHMj4falF\G;5H:Dp]GD5jo>^o9HoZjYa8:<mVYSZ
SGmD>mdn?98G^Y>gL2^[k9Yk7NW0WD<@Pb_;Zl<YSGnq9<<<XM=PEUj_Jj9joB5c
iS:EW[TC20Z\q[:b02H0pA[\e=9pSPWc1_\Aid;[mlKQ0@AJWm5:nG1m?dnm_^7<
16i?GM^dmWLJDMPg3efC;b@ZSK4J2KOEYVi`3cem;V1iF:;MC:gI2oHMkC15PZ=A
KFO2omna=apj:cT\m`4jRP30@Gb2R7C^BWQa6_JQ3hkXI?iIJh:MVl9B\WkhAA1e
V:CWYGnRE8H_W0Ff1lk\S<Hn0?Qj7]@@?G]RjP8=MaGe2ijW_`CZ_Wifc=p\R4eC
Wi4ceS:>[><:ZdB:V2e\dDc7`go\oVC\MY0dZI\UflAPH`l=d76ELh0Y^1]_DX]i
U8nC\Me5i4`e]KIO:Ni2cpUGK`KDMQK8EmdQPMVY8436;ecEH59?`f\aZ`H>K9L5
BljV;V_hoG]96<f\iY4TXCgFiHS\cUnIl>fdBZ=9Q6Y3=XZ5;pCfhleT8M<FinjT
<PGoA7Fi?qJLD]K8K6H5boJBPMj8cP^9gd`o2dJhDHhRG?;R8W;H;3h59gb_ia;H
D[H7:Y8=BWBiOBe9F[[LeZ62kXm>?I3[<q?U5M@i_`3Vl5DnJJP6IKP<E[W=g1`R
30[a8jgOl86@o`6ZB]HoC:`<I]d:Ec871HB^==QFPPb=U5nc8m_bo8?=1gfA5cpS
cK4c1qBiW:U<DH8[2BGoSSbTnLQfRh<MHk@_A>2OH0fNhq_V1]aS9G[4XLCjZ9U5
2^O3X\K9:EX=QVYD\8p:hdiF1MVXE`n<\S4[EcM?HcooP9Z1MO`GaWWg892WOjUQ
F5aQ4[GjLikef]^mgCD:h[`gf;CB8C3RGK6oIP_3ga>;9>\VUJ?T?Yi>7CHblmNZ
AcU_MSWa4:0]ejRb2EUCPa6AQ@o?]<p59H<l_7P_\T5Ug[^gQYB6]k@kZLFU2qAA
`4S\_S0[g5YOgk@6g6T]=Q62HQXlkiW0mgI4T2ig:j6Do\d^L9_`Rj1`Roe0[iAd
n<;N<I]\DVTKTiXZ:NMUU7i8_ZYQf;1ZZl5m?=S_C8@Ek5NFA>XY9\<2DefH6?6Y
FlUNCO=E4<]Plqk<@^;>qgeO6<hlb^4c3Fi71BJl>moD<dH2dd_nobMi];G]6;Ic
Sp=Q9l=__Tk]GD:OVf:3NR9hUQ`87<B>HhcLRQS`HEG7T]pW@Q;ThJQi=j[5AjFT
Nfj5=Xbf31\>DCfe5>47oXdM_7R0Jk4=RJmUW8K`LQ0h4Kf<17k7Xh`Rd6Z^BajY
jHFj]]L46l3f<;27CjAbhDmBok[lNK]D:Og_]De8VCcp2HnKXMqFMj?3]==PA2SB
X::mUOS2O]YV@=Xf>S:nQO=3mdq\4DoJXB<T8YU>O6G3`fgLYV`;hESW?DW0NDQO
c\h>9TqncEl_DOOGaORKMCc3BROLNo5eFOMYWZEG8H^OlpmP=S9l<?:Jj3bFIK6R
Yf<9i3JHWd@d`<VKHBE;[<i37<_Lj;<0O>V<[`DlL<o2CmKhC8cAl<dF7qP0:XKD
b9ENlZJF?HN]lIOJm6;TcAc?YL^\^RaW^JW=e\UeO42@=ABI5Zi4<45R88TB:MS]
Xd1hqH<mHDcNcT8C]2JHQlFHGnflX9l:3H62dR6aqHJNV`IC$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DBZRBN(Q, QB, D, TD, CKB, SEL, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CKB, TD, SEL, RB;
   supply1 vcc;
   reg D_flag;
   wire d_CKB, d_D, d_SEL, d_TD, D_flag1;
   wire d_RB;

//Function Block
`protected
P6ShDSQV5DT^<k3aL^OdYDSgqJW^2JYY9a7Jgo8SQ5jf<=J_=U62V2i9l;PpR::J
m]I5i?5WR_?K?g8_efkb2PPq4i^fjDpl[?Pe:m[lV<N22<?G^UbLKCcD3KnbVB=1
378q0LL<\6m39GnlghHal@@b9IMh9MqQ18Q=hLBLn^GSNV4B3X=8P0@DPLq[LZgU
?4?^Kbe1Y3^ngadLcefgI[7edg:ROCj@_8fPCJMkhZ@Pd3e8ae^?Hd7>Sc4pHoJ=
E4`33]\5I>kC@6nm7GRJ`5oT1?4375[;T_jngl`_4[Nm?i:iQbGWYHY9Y[C0C=N=
QT_24CpDGTCnh]g_E^]fm:5?2cjGMQ[V6k23A<_qEQdedl\dehI9\PENY9l=WeJB
L[QQVogC6Om?2<Zc=5aiLc`M<5D:00\f6RnpcMU0U1[7R@mX_UnJimemMBUQ1h9c
1k@DpY]Fk][VWK<n`L<mCD:J<HbIREKE]N3imZHkGldqG5X@1XPHVOM`d9b?OWUA
]kUgcVMC`Ni3ceam0>kfbmHOVQLoF[0FTNpl4M<ih6qaWd>>kdlm4L0cM]JfSPEn
EPA`VioFE?qI?n;`lMV@>fodIn95c=k8AOmm2pfG]`Pa1qL[T4lYM[?kS9LGIE8\
RgTNEn_n>pj:aSP\]pn0EQfm4pHEh;>4pWk`_WUj<O<C]9Xgnh[=0g^e7p?>5A;1
;7QhWS8inVb0KUVcCh:Dee8KS17N_Ko4;Hbf?3MO7n8VCPQdDRBVjGV[A8X2FSJE
d\[h9d_o\f61Ag:@V2o35NX;WGGZokALj_lnaJ4@qj`AZ6mV:cDQ6KmcUDI`1UPU
L4ZQZEdcBV6mg[_ooAC67oCCo@aJ\I4HZY8clQbV]^\65N35618X]l]`Z2_=3LA1
WSabU_;i?E`d6kMO\cT_2EgWp;2K4A[iImk?Kc97;>h=mXcFWlB;_i;d[C7B1?`Z
l5n^9\L3@95_:6=1ASQBB8k0Q;eK<Ak1I:[:o6YoK;Y3e<?l7GAB^?eT>D]c]qXW
bghXAc<`L<6<>JMUJM\f`1bLXIR<B?Y[D`7168RR7_YiL>QEf`0?OHlPHa=eOLB5
3aQ1eSk4I1_<N=39SD?=]<1E6P6RoLo?9IP>ZEWkpHLF6F<qUk]SN>4mH14HWc]j
dBAhaDYLQCQc;nDdaB:D1Jp9dVRMmRBiI:VGWm?IYBfV4`N]FX6E;GEVX[Tp\G<c
K`j[YCQSjJahoE:T]K59=aok^Ca4@5;6\8^jp4aXF3c;c>Eb0cC4kom8_\A[;G\`
a2JYH^Ma5Z:0DR8@6H]aRqX\o;cBT\B2__8:5[a7GNUBEMc7<3;XQHFgogJlQqZi
doh<mO:DH48PN<Vhh4VDY7\Z]Fh`F9dERSTQMqo6I5iTIM@nbBgQd]Ze03lO[AYZ
i[Mn^o_LL9[nqni9LeoN]2c5YI9;ZgCA8lc;0:5AKFMmU]GB99OTgOj<_g;W60::
Q6Ll`aRK=nN5anTb^FQPI7E7;0]f7lT42B[JcK3G8Z_QX0DhOP_W\3dk<?PfMUVL
>1^VcnCaanKdfYCP:U8EXI^PUf<S9I0qYMOT]iOGbBR\m48OXBRIec`;?2>7o@CB
57Pi@S9aA>HSRBeXCkM>W\Ye72WQ?\caYQ<T6403Z>P5dRUKY[02X1Z[P`ReN4E6
^jBM08Q?7]DUALLGXZHMTC_>=9>:Ao^DYW?2kKDBMX0H_\gVK5BSPWq]=SYY\NC`
7G[cPmPFhD2a]K?WSl[KZ>X@deU>5SZD:d``coImeM?AHg:P\nA34[>`dJjI_4[Z
LI[=U];RS]>7:OL`4gcWFCI6hjbNL[5I=jcM3hE7[m_@9J2;Lg7V?TAYcNkW\_K?
R4n\NdA;28jqT?ZZ<clYSbLn=8@El\nDVXLbAJjAL\f6H[Dj0nm3o:K1o[a6Z5Pg
E8H[8WV:9>KZAlMa87\fA_H1n1Oi<I?7EKN\DLl=lmPi?jVb``D2YCIS>Yg[_[DN
T6G<oGYba:`H1lVQZLbSnkH:=NH8pVBDC:UaI7hRO6GGRXLY:lHB0@MP_1gROA^i
a25_>OnGmVcAULSIO]e[lHII6d_m9H\XBlhG8E2HG@n`:`9n=<RjfMR>aT7kf=8Y
1LHonZ6HdkeUbC]m5\Af2><BT:8M6S\^FNo3i?B06FJK7aM?S`=nqUV39c?8gj9K
=Q10PH2cXg`CX65<hoNM1QGb^dT0:[ileYRC8HBQ?ld8TqL2:JPeRRZNEbfZSZW6
7?<MQhU1laODSDidTThcBHK9gKX?X1_kUdh@^BTLbW?JEmNo>XXTUgIP@WBBCQ]n
bklEE7g`KhfDkEdWoO1gL@Y<cY1@n7`4M6^Q0jJ3UAnilC@JKaaTTRXgi\I_oaN;
XT=ScK=BGq?jM?HBp752;1X[Chm9hRYQ>OgTBMo6V=V2Iij[RLicO^JLeI;KqMgV
jkE`Oa@9c9O_c:5N9=0AYA5X@HA:Tl6jS<GGboCDqS0?7@LcNBA7Hm:XXK2]RBYc
lZ3ZRJlX_U2=3Gf35E9^JiZKE7h2B7Xho@2QA4fL^l_YMK5GPjL=;6lY4ViJAg1i
WJK6B4hIfSH5OVG8WjZQm0S@VcC4A[ZTK[T8YbBMA@FY<fFVIGinqdPS9iJpdPKT
RQYE=agj>fO\RI]K86FLci;XS@YfX^PEm=qa6Y<H<aAHUF1LmSN6OI^Q<dSD?:KK
4I99HV<@ihY7@hjU>:MoGTpmM^:<>BdgJkFWJa8W@fcYIQZ_WI`@5<R`ILi[_Kp1
>`F[H?mX@]Ge:EOOT3BI8XY@5V9?ZnTeKm\SS5qc^5;5WMEgJ3>9@ZU^IKn>QRCo
iIfIeQPT;gI6F0kG3kdHOBh2H7:GZP2g3fmPU9I\^GoT4Ta`apMQoPkDW]\=Y0;m
7<4if`T^g_5FK@LDJRCU:LqI12>56H6ojMDNN9oLViF>HdJOfCdWEVck84RRX2\:
bH0OK6TMiJ>K?7;?@E5QSf@\6ih5HOK[kLpI3ndFEL0Ro1?2nKjTdSlPOnLfW9C2
X_nf=C3W9IjV7OZ3AoN4N7dPfiLlMe>CS_B<RIckdo^KHiqAN3Q`iZ$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DBZRSBN(Q, QB, D, TD, CKB, SEL, RB, SB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, TD, CKB, RB, SB, SEL;
   reg D_flag;
   wire d_CKB, d_D, d_SEL, d_TD, D_flag1;
   wire d_RB, d_SB;

//Function Block
`protected
<[MZQSQd5DT^<F;XJj2l3740?S:eNVje3F@AGPpHYAHPoJ_Y[Q`X`R9OZh`<4m<4
QO]f3MZ[WCQdCUo]?fJ=;D@qD=mKj;J8l6`\i\P9eehH[8HU`Sk041@7o]Jo>KZF
q9T^1ngp7Aaj=R:^SkJd\g320YWTHEkiWHFGRRiY1lkMqY82KX<>QfUDf=@42\3]
S2e>:k@q0o3\OBHmdJag4Q]Pn2eOPcmDTKDApac7?@g7CCLS0X@jA[hZhYKo0:>=
]>;@88K`EFMNd82_LP_A^U<IXLNY?2MKXTYeJ?hL@7;D6CY2q]PdPY`I97EE6>j[
X`B^HUjcBB17X3dR7<dO=P;R:37o3QG<nqHG\8JQ=Mc\43;R0WiVVg4V8jJ<T:F8
>K?H<YE9RqclG_`Z\X]Q;9_<P_Sk5Z51X@j>eA6M:^A2Wq;Ro;Nd7@1dYON?cAq[
;4_<?5\dW_4hfKE4G6m@0hR<E=AJP[?qNEW4gOI>1Kc3S46Q=o57EUi^@IZWin:V
C<1dMe<7?`01fd`\@OGg7oH=12<q2jmQFNXSNkLaEWDN\GES10KjY>VKIaEfe2Y6
lA\LH]W11hqiRf^mGQX?fKJNKa]f=KlX2g29eA6j@e7LCob;NbGQGX\q?VjWcHVi
MR_G7BjH?64L<RB>AUD7HgPbq8EN:UHFB@nFmn5a42H`_BZR2Eo00e>[RIiU>3Ep
WV\^_14p_XJmXRCml^>TUkB@k1X<@@IecZHddSQp_QT9375>X<0b666I0;_16]kj
B]qJMVnO_3IClf95eqWnfQaY:qOc^:d3c6`<jF@14H:RfA:mGMg9Iq1[6;3];p1a
eAfdV`iMoJZ15;PkKHGkH9nT?iZ0P8f0AOHmAPPAQ[O71C>ZF]>dQ9qSj<hBS3]M
]Z1K[iTE]X45PIVZ=AgoWUUblnSFcSM[C4d3o5kgDSF0_5AXH]BVnl36e\`ZmmES
UICHnL`XL`Gm\cKhR<KeGF8oSlWOFSj:fApm6J0LcApV18]N`P>kY:W@dBRZbTqY
^B7`lp3o2e2?9I>FF]SYBK8CmBZAIC`iRgT3En7XSBWQji=3U3FTYif2KoHUjHMY
bCN;OoTn16kSIXfl?ohCE4IP7Xba:LWN5]]d1n0:AM9CV33h_g\Dq^ASJ1R]o\BH
iP?ga]MJc=Y>6SmRSXnEYj;<AQ6nM]i9X8HdNHL5gS0_iH49maQ6Ie5hCP1A^nod
8>bdQg49KZVX^T[L6@WXI6OWJnPkH<a63IC6q6;80Z8I3@I_K@^G76VOT_B]dMYX
\9;4UJ7G471ZnKeJcSU0S@m]R9Kd1L`HiB`AC?b9mH2>?na1Tn^X7i[Lh=`D6`U^
c^6d2lg2U5M@;p\?QaXHA^GHmfcWfA@IGOAFFc2LF48:7=gKY@Zh>^0k3BHP1X[h
:8OlKZeSQ:CVCA\GQ>XN][?kJo\hY^;Na[2YimI7;ZKld7W;G<6IpB9N_OKT\WLb
F[d9Im^X@GQ7I<WE=h5G<KgMWKVeVUUCCkfi`aY3^M[QFgK;Z9RKOBTN1OH1NIOL
A<5b>ISWZ]NoKonUaF`\WEn7ep8Tk<9318BM[U;[:1RT>U?;U^Nm@hImcV2<eLea
T;HQO7>b22^N0`oY6d=CQ`keebV\FFdR4I\2E>k[1I5BLX0Ib>^10V=\_;U@[hXA
J83Cp2@`elX=>\RJa4L`9Nl4]R;:5fk[V1bdVJKBR`DNcd3:j9XoX1UKBbbKm7DL
ph1\CKMqjbWH_YDmFJ7adBXPm4J5>oVN<GRXU@\O4S1?1mp8SZo9X\9ld5j3Lh1H
k[okZH\FJb3cORY=X9BpiBQ>PEC_1T^6Y1JikSZVJ9T4mJ1GBhjD4gDaO0Ckp8BD
8S2Lg=OL3<][>gnBn;8eidP@B5dkGC?VECBKpZY@4PnXlF=eVVB[W`HL\j4[aV;X
4B=>G9K\SeGMqJWFUP`RR:JALI;H@NNQd3W40Zo13Qo[a2aDM_IpYn^c1QU4>k6W
2H^kaZkH3Uq@T:_5kRLYJeXMIgP08Hfk@1EN[7`HlGo3B:6b[VUgL7ci0jSD9>8R
kS5SK_5VUbNQP^Y^Pj=\SUD]\L]`X^?@Fl9Bi01b=VDOAi_EVn34PC0?m72en4JH
3[W8jfT?YPWgA;R9nEGSC24RXdUo8XZB<6Roi0MLjqOEHJaNDMX3lU3RoYYRZRiO
9GmbR65:C4LB@L`CZ0<Jmm`LG5`f<Kl_GceROWQDcEON=e=CDm;eNecjLd0kQ`HV
UPO?=i`IUS=o5mCa>3OIgBXZkgj7BZ^_7S>9PQNK6PHb6WgWMFc3RHRQ5\G]o:ID
;3B[b>KoPFhoFSlPpXO@LUZ9_0c?@PTD`S:M4<3iik`0[LT5_XDR22?bia0G>9;I
NI^1[EOU6aGX@PeOnBnNchXjO;E7aKM^36D[@`G2SD\bL:LiL68jA>5nY5>\WIg0
LJ5dQd_;@l=c9WPefWcb[hQeL11]I9E`gZA9[I\:lRZ05P^@GpSQG\X`DcLBDPR=
\1fQ:PDCHPR1G:LVISCbR]Jl?>6gmDd0gohYZJ>5kk5G\hN9GjN;Q2IFV7Hg7b@5
G2HRM_BNDUIoodk3MF5A4c8aQ8UcKSXoX8`bKZSAnamNQ5WEOSRC^PfWa`X\E=K<
`XaN]Q6LYGgeS>XWGQqTWkLf`Q5Lg;Yl0VhU38;jHI=>a?UllgGOPTVcdSVR1dgB
N;W:Pb<hoGdJTNcg4dh?1;d65fHMdHbN5Af4k0N;VbRB;UJ=j@BhUMFSBjKl]i2<
Y:R0KciHX=c6<4FjLG[m;BZGmBWbK;d9<P3H5Dn7hJmGMAfP;7dn=Mc;[Qp5l5J1
i7@>gJXcaJJLbNQgf[@bf9JXAXGoBS^MYm3Dc=cVPWR5DfJ8QA?iEbj2a4R7HFc5
Y96b8I4;7ES?P[]VH8DS;jDCCQjB8CmG[:BA2DfV?]Md?6C=BPWZ:o\9FQ5a0l\<
0DO`\J[kH1H>BDZTllQ1DRe=oJ[gCC11bcpFQTC2IqE4dhE>JWC:iaK:APXbLe9d
B72m\h@AgjIcaeJ;kBj1Lp3Oh3[m1a=V:F^XnghVYibiFLR\ELOjUC:I9;IdJ]nk
V`q\MU@6F[@F@5K6NeQ0fI9M]HIKPCfM07oMNMKa?_pRX\C`b:YPaGnYfVIA`bf7
5oG0UgS7ZMoVo=GcOjRNE7pP<EkGUQhLN9?I247?QiAO<o5=W6VE\@OIlW@d^>TK
MKqdng:g8D11Hcf\MIcZlKgHm7^0aSneeU14105N0U5]B<beKWY6:Oa@:6<6577C
A]Zd<eV9oiTOe0[_ahm`^gHeRl_S=VXU_lAeLd0L>X>FE\QF>JWWV`9S0k`eXL_9
Lj2K\0?I5^c<8DiPRJpN0L>1FUnTlR?F>Mm3T@I7fa28m\Y8gNIhdWbFa<L1boXU
A46>?b?Td8Sl<74FJM5liK?2@gGIlcHbYU\cHiY7Ib5AWa1AHX3kUY97YX67>\iT
im^`>9^5iQ\Z\4Z<JC02K1?jK:YnBd`qK<hb>lp6^I`Zh^3cWYQOm>?<m=0miSBn
`R31P;0]OBZSAeSo554Scj\qMGB`j51bPbc_XDBcKnncWcUK5bU5@3H?AhYNM9qZ
fH`\jC<JVP\13A_P?No32UiJjUjS;BAAYcI^Aq;3f86:jjEjj3cQHGO`ACAIJ4Bj
>Vb_0MEcf^n3bpiDDKVDjFLUim?_f6jZQfjU@KgAVlO7H`7d?^B47q;Gl:12FHGR
Wm<68GO[D<55WI:O20jH^99J?LVTE\a65bCBKVMWdU^5HnjWHnQ1YH;=[agZ^GNb
qIMDm1G_hiXnGM^JiFklM>O=_Pi]X^kSZR9]>:KlP>Y<P77;f1`CQAA[c7Sb<;dT
@:6mk]hE@9eqcIi9UZ2>RAW;6RmW[:H[SMXEI94DZ_NeSQL9kBKS9KSdNI:WRXcS
4ecZ7R4V\kiTpFRC:fZBFZ298:`4D?<3dDJ25diO<IYB27e0[R8i;eV?Lhg3J^mS
T7gbDZE0SJ7jf;Q0SZL8;Qdjq0NleZKW1DeD_fOlR>K;MjD:ggN?jn3YJc`0Zd=k
RF<G8NL?0XJj9_8ZAKaX4k8EoLdX\\R4>;j:pMh_:SEf$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DELA(O, I);

  output O;
  input I;

  parameter error_limit = (7.11:7.11:7.11);
  reg warn_flag;
  reg outact_flag;
  reg O_recover_flag;
  reg O_;  
  real old_time;  
  real delta_time;
  real outact_time;
  real unknown_time;
  real O_recover_time;

`protected
ADCa^SQd5DT^<jFhEM4c8`B<H`9ePnkde@UV1TJ2_3BS>YV;NkMq`\^TTTnG37k9
GGjERbcPcYE2?kYETN0okIT2\0TkHEWl2Vg_7<[RQ]4meQCF6Mnl[i`6p2:LhP=O
;U7kUD@n<LoYc^AG6I<IZjF?3o\gJT:@Z9NY2gl:fZ52Dq`QlmgTpUmUP``paZZT
dAZKVc\KaO1ZVBD0G^poioFOB>lTU6bGaE91<GMoEe`qhHTa@\VpDXM3dD0:8T0`
ImReH2G:Ti^3lNoEglcqgf:QJhmTH=Nm\J4ZI1=@KGjQNk<q0LL5ED7SC22TBEY5
;8^FEoB0A^Vqo:3[K`@pKB0[FOh?4`ogfkZ8[Cbh:FPWP=MpMU:dXX]pMG<Zlo]A
E3oV?ESUG:N6Vb8f09pPCdQK9Hn7d`h0f^keF4?Z73EVBIJpLU3`]@]A_5LZNZ0<
hi=R87n@=jo_BY\iqJ37?JY2pL=G2a8lnoV@<]g\6Pkp;=dB<>2pCYJSPF=20RkN
`oJ>=GjJDBYHMbO[Hji==ckFg^JMA^beSmH52kg1o_p;bnTlFg3H8jLR[A4>=IQM
SYAMZijmA7eFGepf7S0hDP67o_;aHHbcd\_Y_0\k^h>kAVGWLGGB2p0_>SZk00fg
@RI0iD@j<gHIN;napXg:TBkF4S70_4>qfL;L[jH0lI`^bkOc8ZMPV2mqR^dV>D4q
4Xn;MnZSfgEWOegE7lX\f@oAQ];UG1CYkm;G7m5eMYVUbMTUl]pkDl\_DN11iAR4
`iDM4V25RFgklUKgPK79AePeVE`PDOeW8Mb1G=06H=j<[oJKgD;CYgWjC3bYbAil
e2p76\2386q?jjA0P6]KW1@lo]QIF2I7^=khgl`JALQYHkE6=d0GTZ8QAN<0YgST
HU<Wj;IcQKGP8A:U>Ql8bS6CB;Xq`SP_5<AQKkHGj<@D3Ci]FdZ7Y12Q9P4B:Tg@
0RBQ:FHFk]3Xl4Dga4jhYZ>0EFPT`m\UqbDcEen`GCL`E8:];f7RS6<D7@XTU1Tc
7Rn3e=nA@Jb<4:<27G1d3j]9D2\]:7;dQbU;J10=F\1X3\G87eJ1f24aKGiHhphQ
3fOGLY_o12ZDGb`]Yh=O?fV<_1=<OId]Glh@Y?TXAlO@NXP6SL`C]GlS\4_BD49f
JW8J>B32e:Zjo7N7RVFinEVC2ClAmkONa>:k;ncn9P7d@6PUZh?RP8hCX@nX<XCO
6pO6_g2ngLA]bOk93JMh9pU@UWc=FpHEGP6Y2q0RZL`Kg26BYbFR`BLl7\Z]\POc
2K[mDB39;_a]fUonPEVPM4k>3hAT@\m2aaWRWLYmV7;BF6nWHYp=:bf_i`pS;5\4
:hBFJN5[^90HQV]Lcp[=L]cnRD0RN6VVS>dN6JQT46K>qZ9WgWI6==IcaQOjn1CM
i^[cB7=]HXHIk<FGQ@l9PbDM@f>e0_PkB_gUI3D=jd:W@?b`29DDD@>kRbmVFU1p
5@^h9B:HVO[agnhn>17X<FnqLK2:fGf0odEhjQV7o^Kn:Z3e>6B`nVnjUopjR=G?
LTq8XaMJmP8lnnbgL;eL;<8D@OkB=91gOiA7@5W<n68l8bj^CTB0D?]94`[i<1=L
\B7Pm06AcJ00Y_9emh1p?:;mFX\`;lnWgdNlXBn`;3oG57AFZl?_VcNZnD34nN?6
m\_S3h3[f[aX=5D]_MeJ?6oJp@_9>ZR4A<m;jb>o_jm8KTfPY5iA=PST2:l[ToEL
lFHHVY5;Ua63O\iLBIDJmhgYV@PXR3RYNQ[SbHCc9DXB=:__VJTMXp[1YAWfkdX1
W52I4bd@JWJ5L>T1Jk@2Gb:AdOcZ;JhM<k7Vee=Tk`M>l4fX>UfMB73oAA`<\M;5
a42]GK\F7_\E\7TBL49Uj73BD6C\K21168MORP=;V\;f=[R1UlhBmOi6_pnAj=L?
V3nnRFR2>1UX=SkG5X\GMW<hpTXNI3i@pPHdOb?eqMZOR3KfphX2gle4j5M:3F^D
:q71@3[k7DMDl^5f1n6BU45gH1PQQUkK6qfDHo23jqK<L_Zkp[gLGdfnflbgc>RX
NFALdjX7jPQFa6_RG2dJ;_?15E[VoK2`4<]1a3_MhlQHj0<KKqPFE35IaQPTAMTH
?U3lq2LNQS?ApYASnTS0Aa=A8]3em^cJLQ4mZak5A<[qmJ`n2iYqQe2S:REioEY[
Skm\99bL>Bc4_^1HkmV1aVmd?dX<1_e67G@8c9`<kXJ7:ApQg9\S]h]6;A9AB6ja
2E56mTn]E4?0d_XnMZ^`RjPOMP1G07Y^IOXq86Vj3AIp1_c`LfTSo_nK]BG;blU6
Pk1`JBllMd10fIgG?f7qdZ6aO86qJEe4?Pd7I>KYdDJcJQHBo3>Z`6hJ?\MNC4qB
1jTnVepiGn\7VW`_09E]5UEG?=WN4[nHoF6OkB2ZN03inV5Q62q;6LG07[qi;I4X
cae]LDWSAncN;hM19AjQBAnE6fog@aLX[C@`:[_;Mb<QWZh7BnkQiPS;ZhoD3k?f
l7q1BH4EjqeFfAN?KOP`VkAL41qaNP@^iWqG]T=M4NjTCfhO;Sn64M36YCGqeA[T
NlC<2@\aYk2f25MXmJdeAgViQoCpomZBnGU5@1F53eY;j?UjlMo7e@@05WIeWF[O
VcVpYNBDG5]3mPiVFGMfDKEN\7^oN6]6Ve<;<_=dg3Ek^moKDGOM[dLEbO=L4^c5
I;UpQOJ_XE]q?BOnXHbfq4FhDVCHG:g]E`n:EbREd^Z0CTgjKpD<j\7kUo=d\S_N
_aaDeFB8:9phGLUdiKcqCZFKJ][pi7fO5^>q:38A;=p;17Z=YMi1]AK58@q2X9eA
nFe:W42oBkXCRZMh6LIU=iic6Wec3<eM6Lh[jcc>AbK9[QAG:6lHk1KM>`H9g4Ka
c:><naQYjcZIW5PDL]bcLS>?kIQ6TJ:AODDCO^[4\Dq76VJTbM==@lHcW0JDF[l`
okMWHZgWYW0EN[h9DUD]40b:S1ZeK:^f7GF_VR?T?6hKn5Q\30`WgmfbVWI\V__3
elDp=gnFn_K$
`endprotected
endmodule
`endcelldefine



//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DELB(O, I);

  output O;
  input I;

  parameter error_limit = (23.80:23.80:23.80);
  reg warn_flag;
  reg outact_flag;
  reg O_recover_flag;
  reg O_;  
  real old_time;  
  real delta_time;
  real outact_time;
  real unknown_time;
  real O_recover_time;

`protected
Rn3k5SQH5DT^<U:aBnf=dURIhjmJ:J7L3J]BlFNO50MLUVT3RfQbT3idRbMB7@WG
pjgii98`nN`aI@Y2ecZAUJ>3FHHUgZcc>?0q^[9?j_@Eg_J8`e^foA2iB]Ze>I5<
2f?eOXOKL2ALTJX0=OQKUh@[4Cd<1UQO9K`Q>HlKk9OEq3kaVC:pf[bNC:p4neg9
eSoeednB8j?MO=KJQq]>4LTIGHeaMn?5L7X?[K=Hi7qINabSS[qngSiIekWMZcgK
Na>_U<QDZ0He<Ok5?nqDOUf\KijT=Mk=mWjdMJ_0L3`k]Jp[gR71J0M5ebAFlJQo
Bn`0RZ^=_>pWGh;ODfqGT2jVOG2kiBR54kj>c:UV\@HO48ZP3:^XE0o^4LJ0I_RS
14O3]CM0MNdelHJIO=q;=XAg^[q@61J]7Q\oOIEhNX;<f5=KNaBRJq]l8aMna5OB
@FW=YH]D_8;S72_>80p4JdbFYo;mm7UR?EKV;eYA3C9T`h1>0bd\jHJ=HALA?bHh
0FX\=L?S7NB3:BUPo]c8;9DF24fpU;o;9`bEZ?>d:a5UbaL1>jkfGlXEUGYfpCF^
?l:9qWb0nIbeZZiFCS56dk>q3O6CXZBpdjSj2_MN47dlG5SdY[HNE6^Iol[`JGYG
2JZiiOo;CQ<Y?g\SKcg2JlpIl3gSM6:Wbo@HhX`3F2f^B>?foQN7b@nbcCqjLX8I
1@Jd83DKf]b:dSl60LJ`dJQnlq5jIJ?TUGmFScL_Ln2VB7[D?fLbpmH@M>N7H6EC
4<bp44eEm?djCB[`Z6YT\Q[MlWepD0_=][iGQ=_iIF@VSjDdGfFO1hP`_OSi\VhF
oNQpcG5K`]Pq;_OZ=T[3[i@mZl]6FK?K>PXlFb2Wk3S4]afAYHAD^O5\_YIfd8@>
Jdi4?_g;ePb]E74kPM<8KZ@;U;8q=OGbOZ9p@DOBiN1kjmOFE=9cRLXiMec?>>\T
1Q;9Kcjp1:VC=^o;X[Gc`Z223icWbG0B4YMMg76<UhbiDf]P=TW_VS4ZMhfb;0Dd
05f?h=XQZH`I[<FXh@E90BBdpR_5iIG]V6TUEg1cIBa2EWMIF:m<YYfCP8;XN^1n
aB=KY\mX_@kHl[b5>IgT[_6C?RAFUq3F3>Vh:R`4I`2k0n:LW]R;F?O12FL1N@7L
bHk8:8j<kA;a@n1J12QB34hn^3cZVi32JX4GAOeR[k3H45hO\Z_>ahP9ZopES[7X
@d@2@?d4F<[AR>ghCDHkha:SEa2dM:i6FFc8fJ`<^d?19eH=iEUJajCZ9@9C5V_3
b__XB5U4ce[c;JP2?0;k>b3PH`nKX<@39SC[Km3>IO\1CI<?jljn5gORDYZ^UeqY
798Ml`qk6oUBN;p\RPg5JLZ1d_1SA1VYZ`<`1<L1;IS?1WoM>gEGm7ZCmZS5W8dc
fnEijgE7DK4PICak_hXX9jVClH?pP7ieTj:Te]bo3Mm7o1<R\UfdA3;4^7hW=6jT
KI4bgm7297:Dc\CePe`=bb_\p6amkF_[pDJ8SGM@3jDAe1`o?af;4giqZTJa0Pnh
Co>Yi9V0C3kD>eXETYqnCgL3Ij<I`0U5PMoP<b6;K?LcoCnD_dbmXO9O66n3jeB;
Z0HcX[>Q2InRh^j[2bT]HN]E5fm[bMaj[;m^YpU@kEgS1dI]H6?JHEoJ?OMkP_GT
VUFbh5EGL^^@Am@:kAiS?\:;3lHlj3YDPOlhf<5Aq79MKF<X=_jZY=;;HlHV9?Oi
q@bQC]EWq;MGJ_VQbl4bdA_]PmN[]0o_Ca;_V\[ZHj92UABjjX?ka:eLL1A6hB=L
m2CGjQ26X^7f0RMJ<h>Gc\C_KpK^^_ae[9KN?R^=FO3lE`3LK9DFILZIMTGh<dBB
TCMmQ^>9E`;A\UbH0RGigg7b>HKA0fqOo\`hg2a0^hVU[ifF<mb`ZSR?ZlYg=5nQ
gLXBA5dNYYTR``H@Qd0^dc;k[:RUjdZOcZoe1hT_Si6<1o@g1g;]1GnA>HYp>QU7
2G5G^legRTcY>6jU<@Jbm;\Z@Mei<7DT98>@SY9N2eIgCAT=EK>b5]3bbj\G2>Kp
JO7=;[jFW5<FKSYEgaoX76YncHUa<mQ_SOomc16HRM[cRb;N3R5TnAKNjJTORLh4
k2[@c\be53:jKm;VaGRHh?jkcJ>lI1OM=QY^AGNK8>0ZS:193Y8b9j75gmn;RYP[
TN6p2HkaGY?pP0b`WkCqM2dbi\:q`0lFEITeC:SP<NAHqXWQ967`gCEa[aQI8O5:
JJYS\mAVkco3pP`8T35Pqb>g^0VpfaE8=C65;36:6A:IecqiR]@A=j1bJjFhSbAh
B78EM>DR=:`DF\3DG2:W`CTFG5:=kP85PaW[9J?2TTZi=pBfFcML]qcd_61@W4kS
I;^cR:76NYb6`XdBRSa=pAC0@1C5q8:Y0DTP^;^M@16aWXY?]edl3n`9AOXGI3G3
f1Pl=IC?\eG7[>F@kc\6Aj@q]Bk:87JFSQ8\XUD5?OF>cV0Yg`AZ`BDh=TLGeBY4
UM<CdP0N>j2^p[nF>Ll=[1L?@A>3N\BLEdHKg\XDdOK^GRK7nC[\jj_7:hdQl93N
R1=FbpI\]F7UHp[0HG@A3qZ\d2UMHhEfD]lZCaK7AGD95am3I<M1X4hOpk[jS@`K
po_E9Fn9^9m48_1S:alBohl7c2<aQm^07cWDOSfj=I6<pL;WhXXaqOlLfL7m3gK3
5K[Zk2lpBhK;j7pGhRbnn41DHP77:m7qk>QGNi@q:4N3Ko8nm5SM;aGg=>=qN7Xe
BWo65^CWG>W[cCa<F<TRp67aoH7CLCENAo[Nb[VBfWCJ6c=?7a`=pN3:aF=GoY<_
fV@3cEBO09\i_G=e:Y3U2\>FaBc9p@`3[WVAd\<DP4Wk?F:HdFTFgCiedI?@l@G0
G?7`Qh<q2330CUjqi`jL11EZq_D?656]7PU@T5AP0W@SfDGjkYQH3qNc81:Qdg9j
[K8GL]Y29A1:>Gq\NOeJi^OqkN;_eUW=1JB4Lfo5nlP5n^8qGTmYQ6Qp8VnT9HAp
BdT\U_pbcd4FC\9kBP:TiiV>=6LVZePRQ\<P\0emn^`6:OG:OmG1a<_d;RaF7BNm
d;6bo0IiHBgSFPe3KO?;O?QP:Q:TbF`Z>7GBm5hH?mMBBXNf>dkH1<TUojpbihRo
H;HMUVaH5oQobdYC[?Z2caJljD2`0^@\h@DmmZX:1YQ`dGNCLm@8ZX\iEN4o8HkZ
6dCJ=TREIO1MkA9ZC:TRongq`b8fkRJ4gCARI2:kA[IDL?0i:jJA_@3LQ0I0^TY9
UL0oM:4AiSdiAjFO6i]5\@bpJ9KEAOh$
`endprotected
endmodule
`endcelldefine



//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DELC(O, I);

  output O;
  input I;

  parameter error_limit = (43.14:43.14:43.14);
  reg warn_flag;
  reg outact_flag;
  reg O_recover_flag;
  reg O_;  
  real old_time;  
  real delta_time;
  real outact_time;
  real unknown_time;
  real O_recover_time;

`protected
IG\ncSQV5DT^<DBR_oig;L41JjDa4AT3IB6=YT6YWA>BG\\?hjo3Pl6aT1afQH6k
6Q8ck4FnB;\k2h=qj\a5LNQ9\;Ljd^nZQL?ADQ0]dE]FB>2TN182HV?<3Jb<T4i<
KkJKZOGbiQk7q27^7jMKOHL1WO9>;lPRiS:N`VX@mnO\XoX=pS;ggYmp9830:7pn
6nJQ=]>EYL0[Z@PGF1:O4q7>0Y2eR^b[VeRcN`<gKhD?c;qGbiGcckpfYi6leeUH
1GB`hNBQQN@Pm?49Nf?7oVpP\M]CTVPha0LLk1Nga?aAWIYBOSqY@E`WGgW@b:hE
Pf>>O5MKmTq>4mDRb?mf=S;R6QCg_ZP5;H8eg[q8A45dggp\4g`DiEp7[C:>M_<i
on7?EGJoJ@4VHLPS^p^5N:0RSXmN;`X5DYci9m>FO6;RGUpXkB[U\PWI<6V9jP:0
4`4`N[1CQg]\N1q=aDeY1::;l>dV<cHC^\8W97HFbS4ddFYp]G6<lk_pOS=X@2kg
OGX@NhH1lBpmYX9[QCq1Ff5`^dbVKc:F_hc^FXFm\LdXSSF1iTk3J?;08E9H:HBf
>1`5BB9JGqD\JUU76A=PSGUCd7_NAbKcZdN@_[2;kD9g[p\nj<mZ9L]GfX>U9:Tc
4Y>GDZ=Iq72`fPDX2g^GFCVp5_ahebCg8;4@KkSDiK]n[GlqC=ddOZN[CFlaiOJa
Shln9]WPc`ZU\YX[P5QGZ7>IKNNaRaqi:O7bKgqZBDZnR97e6>B7O3d5ofmk^S9U
_UbM0Lf^JMZ]C0EnkH8XhliaQF`K^Z^5k5YmL77WgnCEfjln`>E;;Uq51k]NioqQ
@5BUGI0oPMTC]7ei1W`N?hBBZUUX4`\hA0S<QPU\\?2]flYYZnJ5W;QgVWoZI_5Y
RL_:S8Dm6abCN`\pOe2o?HXA1oI06i;bS;MSG0VUhOFGPh^b6:IooL<@_T8OQLim
YPenf^J<ln:gFH4IOiUWqUV@R`X0ZUbNN8NgjTN9>oV5g7@]:V0F9k:ESL4YU>^3
b^GQRO^R<A:4=7gXQ2:E@U4chI@gLKaH@oDWZZD8[0ZEEKSYDpTC2OoT[i2dfWoo
JK=k;hiY1]a8AM0XiP>=^R4jgS6b0e`V:9>RVfIL5iP92qU556RlVPPMeR`\PREL
Q8eO0\ZY;8[=3<?;L9hl5X]<=JYj\7oGFmlAYU9;_Xff2`1B_W;5_`27\K`Ocae^
cEWn:fZTAJd_=SjIAGXc<?L=PG_Qi;okJkYcBJ5W:Z=Lj37k@qOYe>HB9q@6C1CI
BqGhE6P^=`FI0df@PadX7@o5a;;A3M3B`Ai\BbNeVZUh_WTbZHW\]c\PolHl3RF1
EoSb3ESm40MBo@pUBcWV:Sd9cT:YZf:^\nnIDlB<4aYiJ9k\IPcHC0[?WocYBbFi
^kV5E[XdTnR>4HNA:hqZaf5^l]q1W:Ce;CQ8XND5J62U\\RkAq5`04]FA2`;:nie
07nMCbVUdnGKpn?Q1g_69ilODneB_3=M7oKgf_agXHgDAARbU<jCHj8Y`bA7`7m]
5NfcMPA;:@IJW[<gco06c>0jOj>FgmWpcRiYNP:Q>46QoJfRkC>oa3ZplRXSHj=q
;L\P_o?L`fVfL_c?qJQX=?]FJGnCI2MbHREU:Y]A_84Q>o4MHV<N?eJ5AhEdPkXL
R7NGS^;G;[`<jZIBaG6K]XPK=01Z<^R\nqd0n0E7MmIH5HRcU\W<KSgg[;MioH0W
khFMmZ^>=OQ0;8eCIZC8Xa`SZIZ^R]igldd2m0p^DAHmYb:4P^A^W9[g<9E;jFdV
3LIK\=@VGkmhhokd?YBM_9kfX=W?c^3\Ta2dbmS^LEXX6o7Qo`9mH`o1;VbKJR>G
6Y1qTeE3]S7GdC<:R5B1hW^dRmKaeAc3ga4ViXJ39i=3=2>BFC7JAioPWU<il7K4
MciLiDH0>0YOeI@RRL:eMZZi6e71e=aD3Q_dXLLdD7<FK@;;MFm>AeWY_VC4<<;O
VV?X[J4pl1D1VI_pNo40Xho5B?`Q[Hl0`PPRDXA@PVXB]So?N3Bc24ka8AY3O2]N
GIZOfB1:jaDC>epE1`R;eGqoTBI5\[q9PP[9lOh6<jgRYD=q4k6Cbk7fHnoT\Y^f
@^e5WP]a2j>QdTLqFeYo8@e8SMGZee<l51^_;?gYF\P_HcPbKngcCd6?IJHX1nqO
l2mXM3qEd_j9BpL0Va@hk0_;1`Y15Qg^p:Lih=WS`\=HcaichM=9_g6[3oN57\GI
9QkainTgEfl57CQ1oe1SV87D8Mj0E_?W4p@I?d7m@qV:o=8WT3Mf6g1GTkTn^m7d
7ijVFh^bp19:_JNWqAk:3Jaj3Rk15=B^dSlcK7RUWd`D:C<DA_0LJkBZC_IFEE22
Y9hfJ10HBAlqoD75?1D17VV^hOU9BJKEINE]c5IkC6873ME\<NEM`VSiMD\kZD5D
pSnIN;cJp8_mkQMn]JbIW`oHHcUdK2WTg;C3dmS8JXU7O8<Wfqk5QWb`Aq8;;m>]
Cl42I?3;?niX\g\dFP?mdSJZab9QpRZVD5Y8pf0Baf[Z3OLlSh4:m2L^KJ4DlTU^
VOK7Z\\Uo87b90Lbq:7:S1c_FCjdX3;HHUIQ83PjX53JgYCpDWedoZ1qTZ8l6kp=
NMOSS7PdabWQmL8pTU]4_@K6=`DFjjj<oT_5h[:\doJl4aI;I00e2]V;HMjiSRlG
l63q^ZOI0ZQqWOj9OeDbnWAl2Vcl68LAFUKnqPo?]adSk0RgH>a?HcQD;aH=h39W
OaL_q[nNe?O=1ioBoP3Ul4fSeIc3ZnUkYCYY=eP7mW]MqdQ_CS;>?oYo;7GN22bF
6EDX;Iba;OdL_p0g^GSYnqJFCQQY^dqOoB34dCLeOIo51kRHT9M?HmSkaGlqnY<3
`QXKKSKk9]F?<kYQ]2bnp3A2k^SUHq<j_PIoeiL>26dPb_GlX_MMhH]m:UiZ;:\D
Ng`^cB83gK0n^b3XkQpZ[d:4g1p`EVc9B^pA6Cec0p2hhXjgYhHKYNi]\[4C\>D6
[TcBTgDa0V2IL=dEo<e1QRm=P7fOE^VdbNAOBlE3b`V7`[pLg`J15Oc<KbR0Pj]F
S]P@JDR:FVX>^nk3INdQ:2o>D>hPaaIfFmk3GL?[V_NMGMPd>TmNh?eE2X;h1dS;
^`ZLNYhPA[HlSj2gK\C_Q64ZE6CCf2n^^fpg1JY1VFHJSaI=5f`?kY;IVCFo;ka\
G3Mk2:;jY]TA@5ZPng>8cQ;Z6\RLf]U:KcchkSLl>>bV2OM]3T@Sc800S:dHe8_p
K6DT7Da$
`endprotected
endmodule
`endcelldefine



//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFCLRBN(Q, QB, D, CK, RB, LD);
   reg flag; // Notifier flag
   reg  D_flag1, LD_flag1, RB_flag1;
   wire D_flag, LD_flag, RB_flag;
   output Q, QB;
   input D, CK, RB, LD;
   supply1 vcc;

   wire d_CK, d_D, d_LD, d_RB;

//Function Block
`protected
<[V9dSQ:5DT^<3jbD`>FD@JF>UlQRSFgpa3PTS3c0NZYGL0A5LcXG7^MejRYK4\0
^L<[kD4`Y[DRWLegn>0Sqc]<f=aL3X1_bJM@8R0FFWfek^@1qTJ`bCPp]BM:<Y=n
3?<PQ[Rmd6Z@_aYZghASSh@pc:`NTJ71QQ^3WcU;:[WAUXKPV1MRL83]FBpfo?\3
35iQZBlN7KRQV22ZUh0l1V[4O:20dp2o3h81bc5HcJk0gYk6Mn1ENf5dq;b=JV43
Dk_>PV3f[@1jA<j:Ncd8qR>cgCTZMkf77UB9<H`fMZcQ^8Fd3TkiZV@>1\jb;NZQ
`TVIKjFLmjSiL2NHSCM^b<CCG[Kg9[CTTq=O27dO_3G@M7Ia;>mOYn[o_EOd:PGe
[;oEIp[8_m7o_H;C4l_fhNl<H0`HbVNdWkdDjJM?X26SSafC15Y6IIp]\B]@A4Qi
LHmWLQO30UaEFSQ]gEF593jW@MLLoQ3JQSPIZ1YC\8>qd=[26lnVA3M=`aYD7[Kl
3faAQ8\n@^=WM`pOMYfNkCo0F]Y@G_3W4e\YMm3oi>IeB?M;d3LqXdO3DQ9lhPeo
KURAL\EIcQ@RHTIXn1kFPJ3[plJT\JFnX;]WCfoVO@7h8YemO;Z[pP2;mT;AqV1V
A6N?8OHYF7eobo?EC=jadPWQhhm\hp74DfF3bd``3Omc^TgdeO1@nnEfJ5Y@PRSD
Go>NGmFa\6PN:\48T<C2=Jmnp7B8@GUDk[YcBbAkb7?Q7n0::?dNbNT6qKYFdlF[
qbQHUoeC9Ea;7Kj<?`_3eQ<gCUYMYq;:gB40`9n:jKb`]@LBOfGhm]P]LGBDaqHW
2NB21p`HfJejiB0KDB<AI3I`454TNMZ4c=Ob>hpeBWR6VQqZlog6=[6bRU3nY?3C
6lldWS2\eUmI9E_NEGOlmKk4Nb[>X]ibYqaCFA@HO1@S6\J?9m`^mKHXT2gOeE9Z
35p5dW>iHapbC<]mQTH_5S]k?>K2Ko?kI9jCMgXYAV@qXKTLUA^Y`5Nbfb\bPZ=U
qA>N3kIHqY?M;bfn3cL0M?YN?qSKQOE3RpO2D<R\>P@ZE:YmjnH_XDTF5bHZqdQG
43R6oNJl1F9:TkXnR6`Fm;HW8Fkjjp_O<S2n<pMWM6PN[F`JYa@Q:Mg_:P9>Oha5
d?l\B92o`qP^o3A3CmHKmoEWALBYbPS`>j^hW4A<=NpX2@_e?2qCMUV^_Qpl2J_D
=qQGGMe@1jTn^_mNo84LFo[R9]=oeX]8K1W4^mgTCe4P=jMm5kl\9dnBk0Sfmo:g
83mGS9C1=MaTV=_FSYcmn:onXiH[K6LFSEVVd0ehIGW862pUhak`0jW<[^R>\oC2
BDO2F<@1^4Y7m>2jEf;OF<jnkZkaaal]Ya]iS`g@R3^fH;GOR`Y65TiLMdO\lDmd
@3f5Fe\D;FRJ\^:3nJ1CW8na\[koSqhb;BK`93j\En>K7HL86kO8CU6m4[ecS^UZ
?n[78CeXO3;S\BElYeU@XKqjDZnCIqCAoDNN@DO;4=RnVn<HTS>_D5NQL_c9bX=:
0<e2pRGW=F6KlgU4kF8F[J`LfA2[Encgc0hG;H>>p@YV1aCBlBjA]MSmPbkHU263
JNKcL2iVB2RP\c[fpdoJoUf[T]@FGgO;NAU`6jTQP52nl<C:j3f\9pe4K`F`ARD7
XADA2Rb\eYe^=]YoBkP;ldReVXI>LqAlK:Q\d0hVaIg^\EK9fOc]K9aV]>Q:nW8f
;]pVSBhD^AJ4PY<I@72AS^_``gCZQn?X>Y;01YD^@;]YC]n4nf\nF2G>P2=nP1mX
lGQ3B:60[TOgL7ci9j5e9>8RkmUSL_oVUD]7NL5o_ElS[j5YBEFNJ\_?i5@5C1;C
[0jGhF6hnVS^PePX?q4XMiVJjRiijbDakQi5oUaidU:HKHdI6H3aLNhhEU^5F4GG
ch]l[RSo6f0fVfDc?00I4GEeWdGoo@AM6h5e151R?<7Na2n:dZ:oHZ:6kK`:4D[_
8Qd4_ORl8EKTMX3NTOGl[Yo9>a<iimddqNmkPQg]kW8kdW^[dadZjh^dZ=U^NL0C
C7YE>@dSG>8eW>Ka=kmI_hLkJG>;HXUOVq=D=CTBb[T:<DSS:=8W0lAbWX\Z_][>
>YBWhhF2`>d1<eK>eG?j6??Ti2BW;Z8PFS=jWaM6;5jAl;HTVl02]:I2JGK_DY[3
?MA_ZU=ZJ6H5;?_RMCWY^YBA2ii56<`>iK=WbO^mXGDJ9[Qf2;RYbZL0pha[oCVm
[60VJZ[2_1EKPGgQd0CGJ;IS@kQHa\_h[R2XZcKZ\e32imfG`S<:LR3\<h[?5?Cc
P]g4RKoWAPA^F:4HC?cVCIXSjK?@Ta4JVP[g8RTef8^@UBHg[MnOW?QP:h2a]gkK
48@@GO4^YSXPPH0q87QEGNM\YkXY`EIc6n4d8HT_@o5;aoQTIFFdFg=0f<G7H8LQ
Bk@Q_oo<n0M`S6nk8aLE<T@FIgIP^XgMVV^A5GMEN9]INC6b2LL]PDG`@hJMbeH>
LCF3eRaiW:9P6dnBeU:X2mOa;PgE\haj;`p=cOMR<P2>5Z\=NM`ijR[BeB2_<?8d
UlcMNhLe9kYO7NWb]QLWa;5UDSi`;_aSF8G=bTSh3D:o:gnGSeKfSb4KT6J=?SQl
5[hP^P09\n:3FRK@eH4mR9\6e]6_YVh<Q48g`1HjnP4a>>ZhYmCH1pR`g9>CqA<5
kBCM@mYcbmL020@a>EP4OI2\o:@d^=mf6;7q2Rmg>HmJ9lh`Ra76k>>hK0CeA1WF
TP6bU4GmNWFPZm95?>B@QG39m:UiqLYCj<fJU;>7P5CcDB[FZ]Xk7Bj8ohfbeoUL
TOTp7V4NCS8g]0QcO`aH?SONL42cDWYTJ=7<ERni`\aJHOf[UQ3En`mFojR^AT\6
LHh5[1NH?lf@^Yp_c1Aed=deTdL\=j38aVHcleKhWS3B_O`nTkKkZT6e2MW2C3g0
3<mK^iQlG]QL0=fEC6P\=qmcFA]fL$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFCRBN(Q, QB, D, CK, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, RB;
   supply1 vcc;

   wire d_CK, d_D, d_RB;

//Function Block
`protected
aObDoSQV5DT^<JhM7S@]f_J0i4;4m\KGIdL^QC\ETS;m]Ip@ZSX>HMOn_RVoT2hg
4jqM1IGQieXaG78dd3LHoPiV[@Iqm5BbXMqHf6=IPRd8F1I[6I=LiG7NSPk@7pI@
In_0`_eH\O_[dME9nhll022:Zq:4F[gLh14gU`QI^FHn1nGd\WGVc>nYTW1PUFmF
Kl8M=9h_^g?YdSjb0GVl75JjZJ8RjMG_j0UTELpPQ:3n:KB5AkU^N\HT@Y0hZGgL
H\PccN<9@AWIGYpcc\0E[?qhE_@Y=pPC0@YDLOUm6cgj1?80=9lK>U^CU^^QOH9g
454Fj:>>p_ATc]O]_eWVX36FTcMinIjo8k7\ZYCCbjmGG>;QQi;BS[e^@f7OCPA2
@L8]Cb_I<Di;8SZJ=?_kB7:ok9132V]Oe2=cj@][gAXPh3oSVKXZAq3R4>::NMnJ
_5^Se7nW<XQT0PNnU]7iO]lHSeaYOa@AZZIA;2e=PjC2Vf>N;[H;P14kb=h4M?O2
c^=^mJo19TO]UJU2Pi`fX3VCJ>25F6CXi`0<q2;<S46p[DH4_@L^hTSh\91agTY?
TdcnY>FQeP2X9eK]G>pP@AK[Q?c1JQAUVZj8_P3O7ogoX77P:7KTOhq6\JGVj?NG
W_1P6LHKIhLV21_1^L4dXd0ENDX]0hp5Jb30[<Y310V3En3:8ncR;E3[QiYVbENH
;0?p3e7]Z7>VP?\nIH`_o>MWS@_V[80mM^9e_3S98b]cXH68XJ6mSYR6<]Vd5Lao
S;=hg8]7UKI8En?dj4DkEh@I>X?nTj8^`Zki7UWYSTfoIV2AfnT`6hob=Hj2RHch
f<Vc75<2jLKTpKK<<gYdJn7nO<gVVePEWcG_n<8XK3S<gD\=qEKbj:EQT<b=9TcZ
O4P0bhZlc>?On]FZal7ml2XJ50>SCk=fE@fOQUnb<V2X<HWLlb0YMN9;^`82eJ^^
WkE?QUR@6;:RffO`n4A8iQkMKGT_LjC^ULggkHgTXEi2\aT0IXQ5`JM3ap17DZ^:
@lAlZ2Z^6h`gMQ@a\9X>3=blW`;[mhc1kGk4k?Q5HM?fTE0@IMFH6cBIoT1lWk5a
gO2YT3:7om=HC]C8HIhh`lcF=`J4c878_T:LiY4o;8CXj[L9>j]hlKa3;3Jbc>W@
\1_9pj:l<=1_?hcNR1?8FS5DSPh<@=ciS91>HYXHFUNXH8oAU]QDA6d:`<mY4F;h
j8Q]Oj?305HmHaXeUhP5UmD<JCl]ihJPhb\<FNg3Qh2NZ`BcNI6AVc_T3PV_RoP>
6e2?PFWIKhOm^>>q]UX3F85W[JCJDEfF::lb[>m[k`15WIp>W5R_KpBhOk1`J;Y]
CnZbdj3O7kM29cVD4`J>L2DbVTK6q[R<J_8Y\kdc1ASVC:Yl9C0TF6ZEHi_l9enO
dH@pBCiiFLOF3JMin1Pgmg7cZM]CSFSBI\2eVb[MbXaKbRo4=T0<SSRcI[6Hcm@c
XC^dOYlS@I\<;Iq<ZamcEOCi8RXKoTIP]IU2Cb5][ecPAaoGRC8X8I0j=d?F0_]5
J_fbOao1UFCTG?@Q5[6I^pRRVPeDV8Pc9N@3fg_C?PpbajB\S;$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFFN(Q, QB, D, CK);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
m\fTiSQ:5DT^<Uo:MXgJUSkG]dX0hc2X9Q<YU_o29R[LC>aJPmfaCZJ9Jk=pcN7;
cPZN]\@DB4jDm]CZOMTS6Fo@>[J0jTeJqWAWmeAgf1o7WUX^[mDqI4UdO6qd7`=k
56D0Rlc9e>aT0EKE8_]K7q;DIgHPAe?icg9fnTA2>7Eo^cJ67qMIfSFPoL6^Se7W
dVK=KOha]Yo>c1X8VLRMSHA8a]EnoQYM18aG_8=ZnbQ^fJ4Q9:G;P=7>V<7DZgBO
qno`Kfj_pbLd7emq]FnBCQ7<O:3BXX\>30TJ5KTo8IJLIOHF3HDJj`_EUfdcCBOo
ODOdKC[Idn@@3hKNiPmLFfYThePfnOdDMlMDkf`5@dPdZ;ITY7LaIBHYOl]3pQiZ
jIIlfKK5KRMWVI@63fV2_mg;ki5I[U312]mRYf`E=dSBj@k74fAX4`DeWnmhUCZC
gI?K5NVnR2OF3h:f]4U00X2MEgn<Y4MBG6=_1HYJbG6pi\:SD_a7\fg\J9`J7DQk
aDOem:YMWBoJ8_qJJa<[epYVZclOSDRJBHgVAmXYjLe\C^CmOaDkm[R2NbmhqMSc
_gn\][[mF`D:4=4B4dYWHFjFk=d?@88OqUEbECK`GoJ2DkTTbfAc8Ro4KM>HWWAH
2GaE`FJkWEl]BOdb8?QZH`nXbRE3Bck2_iH^oH9hJB79PVdVHQ4]D_LgSa[6;cSM
dGZmS1YEjb<_i226JID3Q4bYMb24;d8HjpU<:0NSOKadjCCDN7m>PddQMa0hN=>C
fegSnU:2ahCmgkVMDN`<AU3L>ehngBe[SnU;FV=M1IHH@Z4eKgGU<4Q<CFRJcnF?
dJ8KBaYKW]9h5=[Rdk]XMmiSH1SQ@E7`RCqXd>jh`qDd:9`9>9B>T[_X[5NQ@AAc
V0M9Cf5P1:Ne>F:Xp9g_G3W@8TRD5YO?hC:1V\VJ=iB=P@HMkKETJS6pn<f3CX^c
nhOM_QgF>74j2OeRZ<HJlPFOVE<_Rjlm5Gg>UQcm@^Xbb<T407qi`?3CYXW^ZSbS
]m`=]oNnTc:d;0RRPkhO<OmZJaj[JNYf@9_jeQ_I>TnAH<J:^@5P_<2efD?[XpI=
NK`PW_oSoonLTW7oNRB4bCZdNcADcmCjYVJR3YDk8mgFH[l^gf9:M4Pm[ElSNm3g
GlYOF;Y=pha4ZK[]$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFFP(Q, QB, D, CK);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
<DL4USQH5DT^<Fj:=QOo]akJLUdHJIjje;WoH?anK^^1QbjAIRajDJ=:B:9Gg4M4
I9hXmhMkqT<H5h06nV]IR>RqLT=I]1Rba0=kO0:Qmm<jBLdNc<glE2\Dj^<Lmg5O
j?WQ69l?b8iCj1gp<ldBnDp7B?e>7NV`HWUhe9Ohm\MW^WdklpPkXbH\SWmKFB;Z
<RFoI:h<DAK:1p0KH]9dem;h?HLHUH0flk?b6iRY9=KYiOCKL^ok]Hd>\oQ9K`CX
_l@MJ0W:nL<PjLTfb5Tb\GmOhP7QqKVR8I;9phodd:L`gCgC:VPZH6i^>3Gj<I1P
38]Y4>IlBSTmA5<1npJd3h?9qScmCJ\@H5`UiE;9G4RB@5EZ14i[c@6=Z30H^XcI
>;cnFM9EBRLNWI?X[Pb[jZZF3M[:FdV:iVleI@@GoTEMDBZT3JGI`KfC4c2_5G[c
9T46Vqk5iEf5XQ10^BMgf0RM7@7Mni;=mZIY1GQdYI\nhJ0Y]kP@\i9M82m30h5A
J@W2eD55`I`D^@JaijL6\jeP[LVmmc6>AH`GMNiO75:dl5@7OX0:q6H7TLBpA?k]
9XJ?KJ`:m;I606fH[ZXnTDRPAk_K38iJ9\plAU:X7^c>?Q7S=7XRbXq7JAllglD3
o]aFEZYBPlaQiTcD<oPho>9X;0p?W8^RBiRVJZ^93K_GR;=4<dI^fn`Jl_5TCXMo
da<EjV^JT>K?Jck@]_aMnU_<:c?d`V_8`8^P[efI2O>DNQ2APHAJ9lIfcX\C6ZDh
R37T]`U8eK]^4]bWSbJ^S?kDK0GqHdF3F7f<[G>?H1?ENHlOKE=c6Ug6VbLfn>kO
[UUXnkMkcaafdKTR77X8W9F9676ZV\L90<eN<6WePA=T_WKK_g?`_X]SVbeffU@U
c@k^E5j]c^`PKWFmgR16b@ekq>1D0EnpAl:BLV@FCD:^k3aU;6Rci[\3K>Q37dcO
D<UDG<ROG]_L0OJp9?7^LRCO\Zm[`2Y9a?8dX7VIlS`EZ9B]F]NW]mq:Ejl10Z\W
XhZjDOIXDXdP7XUA0_VS]L6HDokknqXgPLVSmQ14nanRm\iE]2hJ7PVLZA]_9B4a
CIX3@Zajc=[MW96dKl>RZbMRi1jF^T9;YCin:alWpP]o1B5F7odGS2BUP^FC?;0X
Q^DbkVC]hcE9q^3CO1ZAHAJoVX=X2WoBohL]=n9c91UTo1ILCLA3@:<o1;liYIfU
6E1dWSKO`h==eNc4eg=qJXdDY\P$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFFRBN(Q, QB, D, CK, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, RB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
ZZnQhSQd5DT^<FYl@93[glT:bDaqGL]AUljMkD@N]^gP<?K@>@9^Oe7EW;WaqF1>
TmM<RW6A68A8\\fFQdDAa@jd\];;Wd2I=HHgEY^YUDK27hT6VJ;iJEQ@qF:D9?6p
aS1BhSWDh<h`U5`2K_eeUaA^iHq6jP_YbGhSjk^Gb^lS=_j4oO`lAUp8KiE6D>ab
Xj<kV<qSF`ThTQ3abWf9@7ZBX>jLdZL_jKHh0j0kge?De[;E[UGC_iYHZYSnd[oW
8kN]J9A7B5ae@M5<2]AOk4pRPP]Hm=qEN;=nZpLd@?BDFH65V__h1nV]iCf42i01
D1dT>6\WfFTHG1bM8MKZF^P^IT6V1d^QaB]XoaBFC_\Q_bF?G3I>7UFalXCLB9ho
\PA3:_HjBcN;Gm]gKkq>2AH9:BL=KZ_ilB6583MU;cYkM6SPgUBG]NVFQn:;PB1]
j9j_6681lDG`9;cV6b\b9CF>=5m1agA>]7<VFf4ocgX5kR8ZYBcOnHL;l02Bho>P
:pD58B0NGDYc=NM5k3?BeG=e17IRO\34aOS_kPZE7cF\aMf[_9ig?Uob59`USod5
06DC8F0k;9^d<[I5d6;1lkML6\cloOBdg;7XAOq0>VhDCnU<2gHlCAi_SZ58:ikm
OR<DEd:XBfi7K6c1e?07ERFHW:\L3mYiiI92MRf1T^gahmlHUJ\FCn_:iGmcRQ`[
9H8i4Vcok3b@4K\;VqG:IO^@p?\4GTBgA:h\8OnZ786_E7TGDjbA?7i8k\VS0pB@
URWhS0QHUj?B[]V:beFHA_:YEB1WCmBCVTVSRV3_>[0doXRJB2hLffbEF_87?HqR
X\C`n:JAaG:YfhX\`G3CkBhTOE0@\giZ;aqnFFb_4:QVkY6djj?oiO1gQ5oK[n1j
EYcCUEU^H2_Li6JngTmfKUiY6P`^F[IIC=R>>7gc3dDPH[0`ClOXOJham>_T`D5T
ncI1a\SB0:^EHf:9W]m@36eXQCk\[R0Ua^QB`\FW1]kq1ND;1g[iHD6:GCW81VK[
Ta]kETQK6E;A1jF72PhTEQ6N<nlV<gW^JEWPJ8D<7m@;N<0MbEL?hG:VDdKn<Pbg
CDgGKSiP<:m;n1JBeN_CWWmJ9KCE=EkDoKBRYTo`YR^9nSRZ4kIRpK9F3]Cp6^><
IFgi;c6CPD=]F7VFfg?3[i<`:WiXAQ7JUYJnO=q7MhO80hg;6g57F?^80E:C:VID
oS\d`?W96MEXHjIjiq>f49h1X4RMhX0[X[7\@4p<M=8B9Y?=IA[V?OWS:98AYk>\
i207TT9mHMX>60d5K[;5`1dYLjE1];OVEcnNhg;[MX9XA;9jVFhL2j;N?HJ>>O=d
^?V:YJZN0bEHWPEX\5lNbe2FOP]Bh70UAMT`0F@n1hq8jQdnQqnle5GKPQ3aiM@X
Le^4Ol7Yml\>T87CDAb_:Yp2E]?GQjF8n9OVo=N><25igbCfn>m7DnXP3c2IKqT<
7`bl_4gn:X4:\8L9KfM`R:]o3Sj?eL<l:`pNDHG53?4bnocQa;JlX6ZFGKY>]lTh
SaZUj4fPhIRXFGgMoVNl]h19WTYPU<XH9T^[64hJ<HAE`q:MA`J^@J@:\AIG4II@
Q>?e_lKd@ai6WTKA:doeRF;C;Xb8?N6mDPIOI7]N^DUk9RDkgSVEPLCLqD1T]J[K
USnD0AgKdaSO:c8BEVWU\cM73BHR=PUg3fJ;^71mWZfAMOMHCBQPRfcDB2iQ=mlq
n_bL6nQ@OTf7_9;Zg4q=LHHL`i$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFFRBP(Q, QB, D, CK, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, RB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
L36YYSQ:5DT^<`VX8S^RX2OA6^kKEW0emOHnfeQepOC0RF3_m@97IonC0_g^:f:j
c7OX3KY9fd=KoF=\Y9I8_DQ3Xd^_8\P;aXk5G=11GqfSB1:Q63LONT^GF1U`>>43
eSk9<WLBI>i1hqKcEncnq90MD8R`K>`PG8JO7CR2Do:Gg`Xp<U66[c1l5k0jBECS
VB;lb@LYPXhq4QEb_Cj;6keAiJWYELQh5L_;:MgY4o;KCXA[5S;a_Fgh52:f[EMe
J\5<\lZFojNK`YYOI\KZYh3V\jepe:?oagMqF1KLg<pb\`1:ELQ1:>ECD[ANXnL9
Cf@hU:]dFLW2Ij?mBIh4]gC[[TcnU\\XA;6fU8`G<\=FIc0B_I5dEhK`d76O2obL
N2d>`m>nVRGO38CP[5>TD4GqfcEhG4;b]Ka[0X8ABDVG=SSgD8<8j][e:?6XLfWC
>en0]`@K[oS?O2;b6AJYjYCQEc]C<_k@G76iRfKY>c_=hROY=<]7miaU_6niW3GD
kDHZX4q>YPNXR9o4<A11alC:oKVm6oEMBR[YRlJnj\YY6@>R;ndEY3AU@EjobhS7
aDoZ2Z_>CP@X<WPQZ]MNT^:I?HP=Z2=j^>AVa^V@`3IqLEhDNEY7dEh]XWSGKRKO
j;2Gg7ko?]EnZPaWI[d?Y\4KLHPKKOg928SOiASVaCIY?KSHp=QG?c;WaIEP2<o<
4RAccSAhV<XV2jDKF>aHEJ3ELGXaG`:C1D?6^PRTb2IF@ZiH<mARU<N^PE9RFoo6
`VHIR1<K^n`Y2Mk`c;KM_Kbb5kNq<T3VC5p5_8Q\[IhhmB?PMQ7CV_aHlGOm^5j@
IS7DI_ApgI`O0_RO3?Kc2J`ZnW\em[\JOUiA12cS\anqCV?ileGX6ge;U^7a:Ma;
^j;Z\cD1]J0fPXWd<<Km]JZFBHS7Z:lCTj;YQ3ZMkg2;YT7<<md`:P3H>mZ]YACY
nh\Z42>3Ei1HIMdR8M]3W<MHLMb;A5Y@e<Ug@P:CnTDTMB5SE1oRq\BmUkBH]X51
Hn_BQ2?OO4LcPJSaHTVOMV37B^AW3nj7XDC?jJCjWpiCkVn=VMi7Zh54Wa0mbRRH
>aXIW2hM3ENUfB[ER3\U6kWBY^NFSFIR[]O;>AY`Bn403ePAB>?;?F_A=`Hb`Y\k
4^[kX7fmN_7RoJ<F@f84gBL@hn>:D^PAh[nkOiE`9QD5goi0>jpIJQ3H:qF@U]B2
YBkICPIn0P0o=iif`MlQMm4:mm3olAW6MTOdql\e`kOVgF1ol;MZ>Q^L>`No:6hW
eN_68_Cmj7J1S]1pRo:j^OVlS23nRKSoW<i_o:dhQSZfdUL\7JdM>aqhQHn[QW@I
7WLV0@YI<N=m::LSlV_G]E8K1c`9ec4o3lSI>Ci>ET>0=VHM1ZW05Z7`AP[3<B@B
aD;UK`ZUC03=<0PnBaMeYN6PQ[_@hQD3CenXH?IcAR5?LlDhkIm^nCE8l`q]?8I7
Wq3E]42e8S8_b<8b>3[i845_jigJ6?;OWBgX:1p>I]N6ZJA_Ve7Lk9nk_mVNO:k?
;bBUTB3GlD:X4p3oRVmnEVf13B7e`0HZD8H^HYX_N`YKT6:5>Ap0Hib]\lGXC5Cm
d83>]66b\k_IbK83ndM\RY14_n>gGhTi3cHH`CMe>N70W5>CHLon@EkmKkn_Rq9>
f7EbAAc7fBZ8DD]aD9@4jQ3JE9UiNXioBGb=_RX`c9<IKj=U24M?Zn\_20Fn[6hd
oeMXc771pIbhA]NecZ2P[Q:Z?VRKF]T\^In\`;dUh`Edej;l<X?R[cWMA;T]@SB;
n3]BT?=880K7MCd@j9@p<92Q4XCE_?_4chV\AYQlSj7W\N\^nRdZV5>21Xac5:1p
>]2]D:J$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFFRBS(Q, QB, D, CK, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, RB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
0e[_hSQH5DT^<I\bcL`8K<IHT2Hd3jkN`5iUM8?[^8AX8K8`o;N?16q2PVinCDnN
?C8n?8[kfamM[d[XJdP^dX_JJ70AF37_=>U\NhP4m9Qlh<0lApE;CAH]_Xo<fjlX
O`V7GmT`q9EDd?6p0[0OFb4GGhi?`06lQC@8eZAEiHq<9=9?ON[^aO]HD8TL`RB?
KhRl9cqH9i311IDK=IUBQ?XMb3EXImTfMFfLm71__K>h^ENVdR=<Z<9GagKZo1RH
2b;F6bBE^Sh>l3K6hlWFDapLZ;<l:f996eXmM[7D<2=TT6CR]f@lW_TNd=iLiad;
adBj5IJOO4TXlpJZPAnSIqWYo5Q?pd^Oh7B7f9J;bcBhJ@Obj0=;TFAm;dbJQXIJ
BW2nVA`bh8PJJ0KHN]`TenmNIKGA@T1e@M?HG\eGS=5DSP_i2_d89P4=V6W;NdBi
1@5iF<;\Eq^lP[P5_ae]MgoMl_jO[Fe^OciK5j4@8X3I2\FIS6;UdhH_aSYJ\I:L
HAQLkT>M>58n6<aQZFI[0OlJe@nW]X7=l]E^V6JZHSgdTQUk\jO03S`cpSM7[ZS3
9V6<QZeB:gEao`G31_N^R6b@`4TXmn=@dMOea=Q;V;U_kGL3B9VW5j8N8Sa7[ZOH
iNBQ8am>T`k99OXSi\X]5LiD=[hScpS2\Di\ohWEW6a]>6FS;jVXb=Nn=VTi?W2;
Z:j=jl365K:XOUbmO:MdmM_>Q13`I]]cUUod1kPcic5]_YM1^g<cWJSaINH7[Y7h
aUMcV30iqJlVgZ1pn3RA6Y?nQkG?2;ElHE_9LQnTWNRNChd:E1TgqX@N_MDeG3<`
KVRjV;SRbV`m`4dcVCOe_n35qNh\knD@ae9fl0[IWp=5Xh2\h;eDHb7Hcg>PO19C
VUhHdn2<P?1DQQ5hoAShPm]5C=IF8>4L1>2DSNgB59R>D?n^OP7W3LI2\b][d>U`
mQaQGb4TeKg=k=[RAH<Gh^NKNN<nD9Sah9HeBYQid`Sm]<Vn]Hpi`01<Kd4GDYjj
;hV^ED0A:3C[oD?64[bfa[=eaNQRHGZ4nOHF8[ZS@7<g>9Ee31>jZZ[JI`AWPYfK
F3M@XG?bE]T0F]Sn;a8aZ9>5<J1g23OHQjo]43ZTTVf8[_<YbTel5n31lJ\pK4OD
ZBp`j7F_`0ERS4<693[b8RNeUjl<8g\_NNK3@YF?hnbEQqWlTSQ;]>6@keF6Ilo_
T0Jm<i8K><9OCCKPF8KB3gXUDIR\WNDEnYfkblFTSq>h10P>2M2Q<CI^G4d21WP6
H<K8:IbG6e;LZ9CNglCXq?JhDi8Pd0oXCVE;214EWbKJBRhYWREn_`Eg=<9`R_n5
6lQ:XBFDPVgD7nKljoe:Q5ki?5ocY54E@4\5A@Z\B18CL^AoAe^30OXdoGcNP6WL
2caYOdL^0lXKWP2lL6Wfnh[aq;f@l@cq^U;GTTGAEFTXR`EJ@>2@2>nVc]no\\22
M_09qkG1cfhIQP2=@1oKiEMF5PFJHQafFBab94GZ=4WqXJikSGRcH4R6gEEFj]ho
B?_\]neKU6XkK\WBpbXgfLWdJaWUh?@ATgE5Ko]\;W66:=hfdH;X4IKJ6I7de\J<
7Ni>L4@aiVHM9XUiY]PLGD22hfPpD_I_=U1j2?9;VQMP`b8Gf7d8PJ07KX2hbHCa
bS?HlgR\@H0B90>U]ihm[mj3EZ7_q9[gAfnCmnm1<hYPAg_0JCGUhW6HDQKc3F\>
CM5[PnOKPCgI9:iBOPOHUIF>N[JO^H8;U2SPWNmpZ1B]]h_:fN2PHIZOc6P`^^aU
U2bMImN66UF[I=`78m`cGcjY3P5D1[\cE;4WW?8=ZbfIDmpJDTZQc@$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFFRBT(Q, QB, D, CK, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, RB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
\RTQ6SQd5DT^<^I`I2Ua3[>f`6H6CjS7T4oAQ4J?`fOXU38gQM;1C4^GglO\JKWG
Fh1q@ZA`_0OLA5XT?oU75G;2T@WL?N[;mU_Q7^R0C5d[A=60YnT\?iTd?c?Fpd`<
NMk81g7=`FH4C8d2HB^7]ggHf43cn2HpH1oHHmpgP3?ZB1`7al1S]OmbePNMc9c]
1q:LTC[o@Z[DA<3Y1[Gk^gY<Y616<p?2oO`>_SQjUE3[l1877aTGgBX90CcRWUTa
=>OXZa6T4X6ki:9LLE9I9IFUabmD60lIDT2752P];R[oPqL[]A4JBq@^N=k3q<<P
AVO1`2fQOQ>QQYlY=NWoH?<^ZfobYneV20^3ec`>=PPXOZ;41^^aV\QBKSH72_[f
k2Y6VeWBAkm>]fc3288DJf2:Ko]8^nU`<=Xdo0^Bdp2dU^B7be8SCWD[IXMBJmAe
<TokRZ:9oN=1<=b@\UT7iI9\JKWQMd^Jd2gB[OjTGi^7gOk]HbWkIR^2=4lh[>]I
h2K<V:H3Z69[HUUi<4FaVMS]pBm`a:MfnWR6W@@dI_H7Oh;]7Q7VYBm`cSTLXf2;
T3oe^mbF2CV3[_]?_]=Q`j_14B5`<:@TGDdB`0e6_WKCZBHaBPk4DAnKBXJdTpQ6
DfV:i7FG7::=:YnUUopfKZTcUM@T2RAG`C0T61Kllb47a97m;a3Y>\YB`6FXBF=Q
36lV=imE3jofohYR9m_YYWJE;KL2UK1f`FWAI\;<EA6fd6T9UP;Skl]G>[:WAq;M
kjEWpagQ5ljT8;[7Se]F8<4IQP8SaSCV_1L14[J?8pP`]VlTK^6UiTWam_X;IFe`
Q3A?9WCbckO_OqES5ieC5AE8>QARc18n?VIO6^SfCA7jM^a`V]@KT7XR?_1HWIab
\o_T^i32fo>H2O3P0RN9QCg`\iV`DUDa<jFo_agS`Tobc<2VW9KW_ILm;bK`kh=^
PJGg6bY\Jl_h1k_1`iHQO8p;5do[HnaARFMQ1XgG4:Bch_f6Y4Y@l^Q3gG[?P89e
_We=^1fX;e<0:0bl?5GSk5d=U^M;2=L2jg>k:Y_^iI9VMD_HIWWF1Q2iJ4K7hm7A
3UngHbh`EB:6>`iD\[dB?:nj4moleL4qWhae_UpLDOTB[Fj\?@A^LkO9=][W=UC8
`5Lko]QZn_4Z0WVglqLBnEh\PEcOYTa?]qOfOgQQgOhoH7@JO_=GG=800P>U6<@1
IkKR:EDQJ\S_pk59dHj0?_GZ?_<D2LhDO26PJ8R<;dbLY4XXFo2L:9l;hOClF_>l
Hmd4_9<mkgnL\WB2EL9b2k2ca3F;bTDb3Mk?I^fTh4@JIkfQnW4hH=a_\N_`cHC[
jjH0e7G<cKadEj=7pH;Dc;epW<1AEY@4>6jLA50MX]8=Y]eBGEYo]7RX3T=LpZ]m
OOhnW3N700foMH]XA?G\b0Pe?ANh4ZIFK28pHbQ>;aJXo_F3RPcBEMBQ_FfOBMIh
LMi1cZ_8pgfB0TfQTQ961O7olSoliHo;E`1I7d:Ec8R1Z<^=bJcK1O\V2E`8aT\l
1SRfel97R4BaRVWmmK^pWBkkkD\A;i2iA_E86aR8<Lc4Sd?Ka]OTeHGPZZ`e`f[4
JL\e:Tbf?HXRS0]8TG33a\FH;nF:_YpLUXW_n2Rk\8?E>c2G7gkRBLdS6[C<hh^7
^[lj37_ljm;ZNf?ck]kUeKDLmiA^<GA^?70oo;_7`plT^1CMUh>5OMS8aW]_?4hk
@Fl1S6S<`c>hUG1\2:P4;i;DqXD2K4`9$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFFRSBN(Q, QB, D, CK, RB, SB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, RB, SB;

   wire d_CK, d_D;
   wire d_RB, d_SB;

//Function Block
`protected
2SX_USQH5DT^<h=`7mIVinqmZGaKZADQ:<Ig:Eco96L76mbfMUXBVgUEi@G3PS7H
al9C7hM<9PD<8nE@<`_[6<NV;RqU_1f?6EkgHoY^ffo2lI1YeIhMZLL=gD=6JDVQ
0PbZab@j^ADY1biaKmOqH@J;Ejqc:`NmVf_4>LmgBeHPB^M`XDV>Oq1Qa1QOJCBA
bWfMYGSX=2fMnlOSd5q5aI3R4WGek;11_:09KNiIGZjOQWQ_37ighX2aYq;>3fW8
KKDN5eLg?SRP\HoI=eZ=C>bK^n5GSY7VE1K9^OFmBo43cH47=XV<_LEl2^LUgU`W
;`]?5=LPf8pARhh\9gBBJ:T8BbWn_WC_17<GJj0k8FXmkTfZ1cpKS5X0BGf<\ceW
b3geca0decm3HX4WcQUc32pXC>Bcb\8EN>cnAmnfaP2?Z^o2_EZ:4^7VXW25Rle5
DUaTmqLbloHHW?>A3[b0=Focm[g[B=b_:nWY`KPbLOn;DRiN]Kq?@Xd_DCjE\5CG
]flPJch<WU32[M8HW93_:gP5JW6QG`;j\A]0178kojDa3ITq\<DfM@4>441Kd`cg
mkA6=<FAl5\W?kKSn839cCQPSiQUU;cOXZfW>;D6q<m9i948<;gVnM8We?L6N]oH
;li1CNo^HC3HgT]GUfG0_:ZLH\;lg?`aTH4@MO<`<PPSP;81A4:>lM6J792=Fn]^
laT4M9LaK]jBlZ\GjMY6qglReSk2qBo;h^WqMQ8jQILPY0f4o?9l7_GBhg4`mbOb
IkLYfe:[0:ATN`T_KX;46gdneIeOUOHBFV3Y]U;gdQOD1gZF?@lQgn\D?3ZhoAo=
LYJZEP5:I>lRdYP^qZknY8cNR5IdNBi][hRg^I>9SFA[Bk==:SmMISC6;^KW>loS
F1hDaIV4NLJ=Za@>Hf5@W1Q<TGV`<:;6d4bcKRm35ob^XU5L<5HDZTSoX]5m@4Bp
b5GmZH[_oM`Sj0DobMh02`BAS8Ed5eC;EDOJaV^5oDO;F\eIla>BaJCNmQ33N2VX
bJGnZO=9aT\WF94k8RPMdH>^CA:@hDo6lRDSqjAI=YM@0630J3L4hY\o\Hh4cm1C
N3mZc\:QVe[\@SA:_K0KdF>NMAoGEb][:b3CC@4iImIIBG6=6BL7ooO0DfOJbK3k
6:k;o=0MKg^]9LWpPU`<=<;[e:PkUGXje`egn:Hlj]l_=DcTPLi^B_SD4ZG8GBnE
4_\@ml?TTFkZIXSaaN;0lkONaKX9ZG;\5oKTJZIV0lP^YjGK]21PdLijp\dDJg:]
NIREnI44cf@GNQMdAAm]_gPm2\[q[19XP4?`7>CjEHg5eVV2:ajNFE_WN[BC=SE?
0nTK]aYIkj`87<9Tk\T_o7jg5inC[i9XPbib80L_PbS6GIWZTB]f;2SY_;7n\02G
8\q=LhCU_p]deIg0dFfo<HLA7GC1ZS\S8:d7l?=^WEe7iWqJofiodm^HFa8j4RLB
<l:4<;OAlMaVkQnL7cqkU1SQII;9P:LnE\C`9P5E?1ol>n62@B]I_E^b_TmVFiiP
_C;U97EXZLd<c`4nDDVDCBFniFK>54l624cgaSIPn14@V_[OJSO;]14OA^@i\hlG
^387f8Tb9eUfKc9HED2gN>I@OeoK2<nmmV9^Xa>qc6Jo><a7Je_nnbFCSR0@ShQR
:U`Rc87C1Xki8hG8BmWmeUh;M=2^IT;AcL3JWo2@hk0ijR`JP_Lm2`D8XD30lhOA
n0\D]cWTL>RSn>eIc=H>ecD7^83G<X?l^=f40H2:Y\\aWnYhhCj@;ZTVPOmRpnk7
iASpB<GnOAOieBJACY8]Ad1famB@l\W^D;NGC9b?IOUXUbp2DhklBd<XK60D=X=4
UOle81jclXS]T1Ao_F;eGni`Qp`GlGWfn[]VYnh`B5BC[SRD76<GnNYCd?8d8OYk
c2agea6FkX>D4pC8;g6b7?8B:[j=g^OSk>UIE9mV<C7RNDaE?<\B^[o4q5U8<25`
M[P2GnIJZK4dH@6<j>3eSSO>@9ZZei_h8kPpSHb`Ha;eA0HA@?oS?9daZV0WajPa
mmmSTS;hJ_U3BZXGN>NP^EhY>=3kP@cgY\hmW6Hg_FQ@0fgIS8lCiWV]:DIX6AK3
eSGR2R?`aHYjcG]l7VR_leamEdVYo:OXDS^8@=Uqh@iQjKlF::Dn2djW3`O58Yc\
0b>7TDEBB8CH8j\W7b5<5nM`:OSVSIkgL;FV\V6<CZfV[\;HEDdJCZOKk67RAYPS
34@kV^B<@ga@X@6?MR9]d?V\dSXJ?icj_]71MGInh;]8q=5_BhQqE<SJbZF9lJTh
DgFF5gJ8CJY]Z0[0lOEWEHTjq8n@]CfISDOC:]H=H<AZB<bCJLJcdWN<_`45W@ap
R3Eh7=MTa>Z;oV3[_cQY<P]WQAD``@iOG]AT\PqGeORjC8h_E\<QX:5nmQTEZWN4
hjGi;lkk^J;NQbR\@GqC0hQTK^X1?26X<i:a]A1V@jWjGf0FiCee9Y9emq]NbV?5
OjR?7??L1\=_2CYkiER@21=jKDOaTS@MC_R`6[^\3h204J=OjGLg<U;OF`=oET60
TE\jpFN[A?VPROaRT[eVnQokHWoG4]=>KUCZm=LSa^dYXa8X8f2hiOao3J]D3P8k
d9OU6@ga3EEhg:^qaAg2T6D\K`^lWkfA3>Ue3Vb=GkbSfd9EbFEKdoaB^0dgm4Gc
oUb]fNaRM7\Z5>K`TC[kKLSig2q;a_?j3CTP52gSJXm26ZOg`ClBh`HkL5?3==^\
]7e3e?HCXF\oH1hj0CWhoE7iln5M=93o9pYgl3bi1$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFFS(Q, QB, D, CK);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
=8F<^SQd5DT^<c3iBgK?;hAB`HgDAh0^k7`q;d0dn]DcJbd27d]eLSYSNN:Ic1Zm
_^QE=@K;>Vb1nK>^Z1b@ajOE=S@liKOi8G9`dgq:_c1j`U<UJChIE6aIWkB2SJAC
Tbn:O\X3EnPh0Ck>5Xhe;@>NS11@2\d::_cV^qMQjNDHp^J8N<Fd?86m17Odj7Yn
g80U?=4qJ4570of?iL]8dX3DI@b6;01^?MPq5ZPVKC8BMQN3UL:Xgd6:H?RdO\7g
j>eb]mZ2YlYg>S9RXWhC_YgPn4Um:?g9EALb<5MLklfbNF1`;=qJf_4coXqmZGeg
1q0h29Z0akRgYj8X?5TU>JR?FcS<DNLaq3g@[k@jl@;PbCGH32Sgd<[In82l[e[6
EHPn;jb]bcIUePBYS1jNiBAS=ZT0hcdWFfHY3oUSWAnUGIIgdGffkYkCa4n\7=:J
:L_XTGZBZBHEQpmPHkM\ofP=^f5kEVec`d1o5<l_j:FGgS@VMR^]Q:ZRWDVGiCjk
^GDUl8P[R=YO4K9Z0n4@037G38?g3`OCjoVf8CXk;aRBk1h]2YXSYiAIGYHcpAQP
1]BqA<SkWWec^b@4?o?X3[^ge?LZNI;RBj::GYS0SIqL52N0LAJLY:FUZ9QXSae1
Gm>fOhEH5lf:j2qHZXaRWW>898l@Yng<h;Q?<:Pc@RV_m>=U^XI<4Kk;W6:YfNR6
f]cW@ZPUXUO_8KHToaKAm;cq`^VZC^Faj3<LT;QldoNWkm=2b;C9H:lN4:HeKI9`
fo<I<@LHLoHUW1AL2oD=@;@4f1AUWcP27bM\FY8Bi;<Y89bhoo0KWbXi9QV]afdR
mR7falT7CE:E:WA13M\8N\<Kpa8fE0C<C7Z^oAhKC2OB=kUA0AINc;^_CeCK;I2D
ACN^aLJUbmY=Yjg6M=LB3\jdM@OGmX`;ARLB?1PCF[<ANkYUEX1PSVDU[]`RG7ZT
S:[TNCdA8V0QE0ICYlho^AK3Wq:C1`?OpTO0[\^4HR?U4MhA:Sahjf0\P52NLXLL
[=U=:<1pViJZ2^P2VWJ@>FIe<MFA\>LJhWdWqGj]jbO9Z0He0B=`IVRF0HPRG4lb
D[3;e5Faem6pIVAf:h@2P`kRcTZIHbdGVaFDRTjehHgaOC3`3=i`T_6c[C8Bjh8i
]LPPm`KENlHZJSa`i5Y3cPqj>AMJd@FE>Q@M=a7L`7JD38=9G^QOhhdflgQJP47>
VZSgRP6@l3M5j`NBZQSSHdUa04SkAWj?hqBf^K:VR$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFFSBN(Q, QB, D, CK, SB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, SB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_SB;

//Function Block
`protected
WfSBLSQd5DT^<ET1G;<Zg^L`DT>?3Yd\cM?e2fW7X\i??8MIq>iJn4m\jiOU@cl?
Jm5fm32NY6Yg5d2TYpE66`Ec8`oaHe:9P@Z:?:RI=BcgblnTDgG@h8TF0=N=WZ<:
Jm23]D3Yae3nO7ohTpO_JbXjpcV?8da[01Oo^hO]hBi?W8PEL7GqbV`]A=LF9G;Y
^NVeQQKg_3i7``\q?D^:^037XLKEZh2^CAoPml]ga:iHXAk]f:0d[9S`I70:1KOP
kkm7J^bV]hF]CITdOX\Q8>FaEcl_GLfpc:U9i=MI_8\:RPQ;P::G[]j24LP[X<od
X2DHbFAXojM:lk=UNFh[p50c5[X`qTXciDCqfoQDSNLK46:9YKETnOUk?VObKLUI
T8<XajD`=Ak6T:h]h_FTZN?:7fgX3QaWbKc56?BC>a:cI0jB@DglX6g`NQH34l6=
1CTAT3QMJPM7bo`IpHe^6`d3\QCNhB0G3W6bRX3_02_a<CB>cdU[54\5K^6ZJk00
34[ZMG=obQCVS0^qV2SR70VhE<;IU4G>Fiil@GYJ@4Z`;8mToiM:k;ZjN:@WNC?9
XZg:n`knQTI>UjiQ3_@DI9lURI4MX2<9RNE<50Df96\<SWnj61XMEenP9`dMY2qj
]4lW3O411ZW@9B2eZ>oOb>_0^4`OG2AVGE4Y<GSjXGP<8nfW3a^:C51];fQ\G;2m
672b3HA1P_S19<6a7_:aRHT_:;Z[5l=adLka=hCqVLW0jFZEg`=A37f2NB[NW<Tg
FK\MI]KKO[e3S]OIcc7m^C6`W\k<OP7B7I[>^_9?VjW0jTY9h`eC`F]onoAj`gQN
TScImKM7Z;2Oe=qVCKhD2pJ\S_aJa_UUIZgDZReKJMVL=23MD\d[MJYK\XpeU@M[
_]HK]a`JK`Lm=YbN=EUd3UL3RX@fIgp<\Nn9W<a2I>ioJVg@ohn_hQSNIKFi?c03
K3Q7H>dfJO5<0g3gok:HE>>eSHTRJ:0JDk_mfoMe4cLCg:2Xe<VBN9>_mh;^GIIk
J9hgV3;N2ZjL3507iH7P?ePj@][LAD1a=3@@YRHpkU1SQII;9P:LnE\C`9P5E?1o
l>n62@B]ImE2bfThVFiijeC3[97EXZ5h<cTAnDDVDCOFFi4U>54lZi4YIaSlPON5
@j_[OJSO;]^YOAo@>f9WdW?2LK?=?>`NILV@R^[PRK\OV]<epL1;I>]9i0>QcId<
O<@V1m1OHk]0Z?[kJ9;UR=;:]bmZg^>`6^P=ZYLlcqDQ72dAqVS:h02lmAf1M0ad
>D2_BN5lnHO8OASKITTBIGl3VHNpOB[a>30df^RVCKo0R^XFHBS]F^CSPU9mOn38
GQ<>ihpL^^e[f;ne]8YCbC_l2W<0f_[1AG]e<:51?Dh_o@mhbkTLN8>JDXTL@oIF
`]9YB^c>l4UVY2;5@52KoDd]h0BHEJM>@e5]M?DeGPLo97h7DMPiC1J4?KE?DmT@
kU?2lGEL_]gp<dd5dGc>aTJe?U5qT:M4a2pIG^:F3`3dPPhnO2NDgN1gA>?JgYl0
@59[=;`[2p^?USjaIfEkad^YGU:bl1H=dhAdggcZR3OUdCqN`O0^;EL^?5WdDj91
UPm4XR1n`d:K30_bnG0qJH9GR1gb66I?a\f?\BL3f=Doq\PQ5MWU:RoDYfGGbVo0
YGQFiDOnFNIQdo;E]017GLBEG\e;nTK2`@kO[JXcX:6kB3_G7DC628TpiBK1=]AH
hR^`d8>[@Xh:lJX?7;[lnf;=JIYkoA;F^<Q8Ag1UPRUCL56j>F[<4C5n8l6cK`I6
4CqTojRXX`Xj8IVn<MZ;ah@36^9o2VhT?b4jc6[_8lihE26>O<i?H67WCnC<hIVR
Z0AXI`1<?pcT\EK9Q$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFTRBN(Q, QZ, D, CK, RB, E);
   reg flag; // Notifier flag
   output QZ;
   output Q;
   input D,CK, E, RB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
Ja=dcSQ:5DT^<W_i_ae62`n5YCEkNg3W^hP=g6Z=W<738Gi8UmnoEjo4GB_F9oq0
OhS[;W7hEI?]^7RY;JO7mQZX:EZUmh_^KpE<oS3WU<]79FKK2NLWbQaIOJSSjXdV
CGla]:29_FOD26GQK1AVP^jK\:gdqSJSFI?qAg72NbAb0Ll=a]UWWVENSMeSih1d
=D5W^<9[PEDVRNnnE@L8Xc\^K49N7Ed0[FVHWF[lU5fW^Uj9gjaph6\`fl\o3B61
7M:9:DcJ^J\d]1qXCb[CWDobFEALde5a=1kAEM\mQffO6Sn7iQe48CSZ`7p;Di<D
f_jO[^]C2ET`WLJ[7E4QTHe`9>Xpg0<?h`ipimSCnkq\FRR>89g8CKGiSRSIS^mk
QnfVNU6L=kJ\n?ha5UJD>a;VlJPqV5mTBE6IMP`B]ikXjK_OL^FiVCVY>_IV[\5I
JOTi4FFR1X_Gc_dmF:1B2A=7bW>T;QTkTSTYYEKJTgX@PC7o@N[AOQn7n12>gh\g
9P1Z7FYEpdJ3B7W40WliYnAGm`@3653[jP\kCNOeLAA1W6X1jiF=V7c7G9T9KKh0
:E4`TE3eO8nmNMVBPkR>e@\iJ5YH_VnTE0E91Fd^;0`G>GGD495liG^plID;mFiR
<mknbNAA^W0JjK^:;5^HIhIOBgIQmfdDLZV\`n8k12ge_gQh1eFc[CRNl8DCmL^f
``Qf:O^Wh9k\L:MdM<^>b6c<P_oNqKb`l_1X2T\oLC\nQIUYado_2LC8EPQ0bGPC
P:T@a_YCY9C@c61Eg7kbHb78\SS@aC`gPDUAZ7XKIlb9CkIX[DJ8CF9YUoNlPK8B
8n9ZGWQpDJWS\aPi0V0EZe0KoDOPHI<cj[F\n]]UCTjK9RPXlLB@TS>I]WDn54_U
OHPGoSD;^CEZPP@1jgmWiAOXjQnnQ;89B4nH@27^iK8^>aHJRXJ>nanNk74;\5:M
8gC`O]KUW_87TQd<I<Z^`;H4??l6LT<b;5Fle]ESPUBH[YlJGBlf7DO94]Y8_`AS
Z7cWoF6PPf1@3I4FqDdCdUEc4KR23;=L\RU4:qG7mTgdpcP@c;CE3c081@SYP8Q?
QE09@KE?<kOIL@Na8qQ]a>mdBYdHeD;RG[BYEhLYh5JRYDFl5=gBLpXi0Y>gWFS`
7@XPlKa791f3caG:JISfU6\5W\NHfcH::LJO_Tk_I7eVk[l94HG9\?d=kOAH9?C0
?D3?_NAV=N][>J]`jUl5EMETd?j[30ofND4Z^FIeb8G7MPaHH=ZW_79Yj6OQdXp<
<dC[0V??ejdoD_Si]aZ5:ci8YcH^?H7E;Ym\MN;HT^I[GPh1=LA<PYcP1b:[16W\
K4]nVoE;GMPem7^V9BTBbHY79mCiIPIRI?7E;F[DB1?Z<5iIfNKXR<ZIgm0R]JYg
oYC:g4cp;UVgSgpR;3MIG\O2[K:`:9;UiSP2MO^_\AXamF:6Ghm3K<3_2p@=SaQj
3>ef^D7eA`5;A0BU:A6AmN?j6b=Y?E:UCUnoq_=P0H<Dh\cOigPUL?U@QHN99jjT
\@SXeemRQqE5W0Ln1IZ7^G3_DiI6df9T<g\h_mkSLlNcZQRdl?oPi@On_@:=FANU
gfXaN^@kDmh=KCoUfla39P1\F2la9<MLhcVi6<idPg^\n3QK\4EZJjPORW<=9oDT
49i?@?kGo\8U=qMl5Thmq0TGQeOn\CVFiW0a0_YL[ZRKC;2o<f@G2V\Ifpo_GZZB
dm;@VJlCeB:Nl\>b6WGg212P=kYFNE;PqU5B<::6fmM[hY8RjOFPl@];>[]oYAn[
8oJ6cq6ShGJ]eVT\T_h\XEnk;;^>80b^F^@TiE`3j@a3iPX\cGgTF6KTb^Km3eUI
?I>Gl\Vm[0JC1HMhq=gOlNnDN[944@7OQVj0=`QZJYbm^So3A5Y<[H2B0>IX94K;
_i:Pah9N[OZ9^]71>Y9`J[HMQ21pRI5Z3F?fb6>h;<jU6goih=Mom9jDq^8W@:2b
Bj6nN@eWdBD;jMdGm>ViP^3VdRVHY1]OSFTPYV`>>9@ek;dR]a\XVnNGloOIAW3:
g9XqWQg4GmE$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFTRBS(Q, QZ, D, CK, RB, E);
   reg flag; // Notifier flag
   output QZ;
   output Q;
   input D,CK, E, RB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
TiRn^SQ:5DT^<mO]E]A469:PS82IY30?^f@\90=EPnB8mm3=9?hG`?8FfiK81Z?i
AUG3iD0E_lDlpXiG8BJEPQFVn:a89bVUPjn6U1FTV;US\BZiG]U2FUih8;W?BEn`
e=NnEdilL1BAmk;=pW[8H6BQIb1l`7@8lWEDQiA2FVNINoV;dP2m69NNkqC1XI^l
p3LDI\l3iIQ98:Tmj;;\iH\P5m9No0m0VH0O0CH:\]RWJ8@3HbF0Sc@eb;i:Ad]j
Nc9X?6N`Wn@hKf;apAIKc^L20a0Y\iAB=XLhdYSUBbLq6:@TWWYBg@fU^289o0hM
[RP>;j4nM7bXp7N2E\aRpE]\?A`pdM1KbcfeKJHXomCoON?2JSmW?;bXNJb[oD5N
c:ekWF`6U7kkP[IAK0:<6oUmDi0BS1PF2BiTdGb?f<KPo`IolQ@Aa`Z7QL]li2>d
SNCOh7;SqPDQjPKJZMQLemZ7bneZLW7KS8GoW]<dPGZReK4cICaZNaFLbk4nf0YS
`enB?K9e5\6[TJRSm57BS2HbVaOWk>DW79O46^V[=5[Da2gd2JiF@beq8UjcagW_
``6h?Ed_6inDeOlXEZ<RC6=MZ@HWY7>B^3VdgJHS1AISPb8[;0=h8eE[8njca@C]
Na@MUPGPFoQn5BnbY>bj=C5ijlL?pX]\0fcZcnR6m9F[Yp]9C^D][ag3HE6][JNR
=[;lUKUTQ:L[B<\=2NTL4M[Kd:G03\85XQTe9_lQVJ6=4F]iC?D_4A`l8XoP^E?4
M_RjVMVFah0C]KlGnOUEplmXf?19anGeoUDSKh5S2WNCiKOl[1?O@hdehM2oi]mO
]=_@Oc`GbU\nA`mJPO5TLQ[ga7TI2]G1P[iKjSCSci2c9Zg:63@0fV7>=V\]bYT1
QeU9A9i9_Aa:LTT88TMf3[T?GB_5i5agAK=lbMBmkbcCZ;Nlj[?L9oAmTJQjD=aZ
?QH_e4`o@O`?bE?moOKo^OVacc<kiqa5a7fGpJ:\DIMTW:I_R6HWC8@F@]J5W1QH
26CDKlU>cpUf<O3G77m]hnFo^U;\77Xc7GL@^a6BVAXZWpOI8`2^K_JfDdghb424
<USM`7?Bec9GDG_C^Ge>9YGF]_MIWd_U[hN_TI93O7T0j2FYBAWYjlU@[NPB1o6L
UIY?If9l:T\V91i@YdZTTVR=KW?]B8>Aon1e;R8CNICYoVcUC480oiqeEGOc:6mO
o[g19IZSo=oFd>[H`fKj3fcXG0lLNMa45N;_PBRLF_Olfk[UC?<mKCjle1JoYfam
FR[NOc_>P3DB9nm`BahdE=1?Q5N4Y8dWVX]l7YfoLOi\GgE1PmJ7V7E_KU\8^0Ap
<E[nT_pAmj9Xik<J<d<mo4VZCAXmYH^NdNlN?jW`BZH<7dBUlqg;16Ae^4=I2Cj6
1qgTRFl=l2J>JPnSYT\Nc=gnoV>eC6i9UUF3WM?KU`9Ap8;chCCmKULa>G@Sg9]P
N2g0J<fP5M@5JIMW:_;h@^K]nieiCQkGb\9dV5X5Y`]9eP?DD;jb0]1Th`I;F4>S
PU]f[C\[5L53MWG:FXnCJc5l`6[WL0ZNWOCUG3WFE\^AJh@\pLGiLFRqGVCcQGWQ
ZVE]LUFZlP9eVm5Q1S5C\H7g>dJDq>[7m0JH2E0b]<G2n8N40gZP3R5mGj<]nZGC
UgMZPh>\e3<^WOd:1R]3kB?C?JI:=6oRf9Bpg;d:MEWcOXkdQgnMX>lmK@L_I40>
6_j8m]nf9dqEbg6k<`7U3\;Ukn8V8a\TJ?BAP9e5:7kTTGBp`fIbY_d?:=J9@XWY
`HBZX[oJT@cMD>X:^k[:Fgih[Ma1:92DBJOIfW]ZifH@;TDS9Ubn;@K^UCpLThT2
T:>dO1:ZnlNT]^hhh^bXJckD`g2VOVY]C0F:`3Rh;EneC<M`U]D<1c97EGGCO>]^
OPIF`q?g]YOSaRABHjlna_o]<5L]?^ma2GV>GG146a[a1jA;j>\g5R8>a^:TMd\3
[Oa\VXG8DNB_pe9Lj_jo$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZCLRBN(Q, QB, D, TD, CK, RB, SEL, LD);
   reg flag; // Notifier flag
   reg  D_flag1, RB_flag1, SEL_flag1, LD_flag1;
   wire D_flag, RB_flag, SEL_flag, LD_flag;
   output Q, QB;
   input D, TD, CK, RB, SEL, LD;
   supply1 vcc;

   wire d_CK, d_D, d_LD, d_RB, d_SEL, d_TD;

//Function Block
`protected
KOj0_SQH5DT^<40YTNjI`7dIB5=15=q7DjJeGV0>l\9Wk[IjQgO4[aWZf=aF`1H[
ZZRbm^WT57VQief6obp;S@m^mcbOOF2B95WV]8>?d0m6N1cXBVZkI7p0PD5cnpoe
WeYCI@EONmm;oHf]lU?5IO\ojaaaGq:0H3cd_T1CLQS1o4?RmWnn9f>Y2[AT@`V4
pMl7RbfYY2lWB:eUFgoGfh0HZ1<X;S_lG5Bq>lUD_D:Kk>>fY5V:4@Y:dJ6Ra233
?6FX?8SXpMnch>eM?Hk18?lUO>VOh5_eFf4JDnhC\@mqG:8W[JhkiNJU=HBZOd9R
n04ZnbqY[EoVIZ1D5S5Kcde?@RbO]nDGkTp;jh5\JDNH\5:<Sg<\S`mYJpHI;?SS
h8dENke\`g:[cHCiFZoI44akjUVG\HH`:Va9L6MPD?W[GGU^[gf=LhfXZZ4OGWV3
94[Qh<p]<FS`;_eTh[fZ?@j9M6kC?gk3:l9ZjIRbcij:6mpc^]QCPeZnm>n_Rla^
jJTnb_gAPQLQKA\ON?Cj_=1JOL:e=73WVkmplZ<GZS\g5Ed3khb8U_dZagk^7:m6
RBH?hm]L`2`SdGhURjf=434Q[NZ^?]Zpe:IaI1;AZ]3O<c[WUU2ecC;HfQQ4eQMI
khqPN5L49\@_B08cG40ELHK@3GIc61AdKJhq_elb_LUDXB5]o`\R>[Bl36L53F=@
[idc^V[Tq^K<VmhEKo@BOBX;?P:8Qig4:e;3nhAZWFZHS2m`q;8D4;Za5hNS[mnF
8Ac\RCO2?<JB4oRkbhb5dp1N[k\GKC>::jTjCVGXKEd\;35gmM0^EQFDOUI6q3dQ
O?K>qbT1D=YIWDPO1??IJXQ9l@8^J<Y^d_S;`B@SeEPX0ONRVUclI5IpOF:_9V>B
V@6fO`fS:EmRVBnJ\DLnVh^c:RDQBSkl`k]Falh5ERAZKROXaK9YZhR3OI1LTWEG
e6S;W`49:EYPqKbTh6[9_NkKlT75KSfFNEn[n?]NM\B1qRVd=]U4qGTV_[Zk@^m;
dUCUH1jh_>EfEbc7Qn99qfk]We6\qDe[n]Em6M7OKN@MF^\eIEX>?kbJ6bCE8J]=
p362aD]N@QNmIF2VIbZgWI007bLWpDk<N@;YpL5?RAH0eHCfE00BcH8DRTBU\aPE
NFb1lFa=_E16hniMQn@6acW2?baaK?UqLONgcW=OiL6D0Pn5RdA3DZWKaT>nL6e>
L@F<iFWYNQ8TlAbMXCOFD>ML9R0^HVpB<GnNd`^o4W>@>]QW8lliC[=FWiJ?3:Kp
k4j>FX\poTMgPlJcdVlFQXF_4@ClhbG<^QK1]gI`q3C[:_O9q<9RYbbkGE_0Y>l4
EXZKapI\?85QFReoNo5Q@`JAbVG4SOI]:_VXpL@1C[KMpDm_SnW<OO1b8WY05<Tc
MKW>NJE=<qY`^TU8PET^^i?ES2k5Ph`@Yb]?T56@Of_epd5?lmASpd:]I0T3@A84
_P;IX2]YnI_i7ED`gA0M<c6pAZS[UTJqh<8_iRlLi<gPKQimNhSX5Qh39nHmcFX\
I8eG@@kc^k9OGSP2j>^d:JcCDKg^MAc;laqiN\E5HWEkD]GbPeGVV^;a@>bH^aJn
6^SkI^d5:CQ6MIq3U460YlpOQa1\NVXOKc`U>AV=2>Dlao^]?4f>L89:`\3bTS@4
8fBGOJLalaMQ6Rc;R>TT8TZQ3>[_A>9LZANqWXDnh=cD4gSYPg`ja\7LX5iU]@6h
6EYBq`@di89l5DacIVKnpPacmKo>p5K8;B>>A=CYX>1h2AVd^j87ZH1ncBMbMpo?
V=TaKpc<9\<FjqcMO4h`qCOF5cY`4i7iS:LW2o?o1\<dLd=LO;Ai1n;0Of0D7=P;
C6FKDNeJP[<A_k2b;0E54ebi]O0fVKlV[YD;>cKH`ZL6eMVAN^S`I@WHMIUmRDSZ
]q<@;4dUhlfQoUV?nWGn7H95`gW>lJ1e;qX1159\<;gkXm\Kh=5KbnaC[0h;k:I@
]@BmA_aZ]7Welin4BGPX9cLo]Eh1A?fOC0jK3jiWG`lB@FdA9J?BN?nN@G4aOo9`
gP0`KVXk7Y]cGn]=pGT0b_lqPSj5m>`]AEJ8E<[F6NoL5nh;H=?2<GG`W2e@WJpH
Cf`b[=DgOE=k1M^_ccVeX21Bf1llUlC^;[qLfmfIhDFj@\V5??WDOZ502me_74KM
[MDFO]j]W9q>HfIAEA6U>@PB@WUla8>o2^4IDc]fknaNg9b45WO5\Y`_]IWqCj^@
N=5RcB[:0MdaH38Rngc6\KDRk2>F@QRgp`d8FHnN]g2bT0FlLW5P@j83J@XRoM_I
3ALkBAY7q;ELbDmFbTL1A<=>RPo0;j9QSG0iSFD^hR?TgqnHQd8\lY8laEW;^ai`
8UnGff40R;XBgcM2Fj@gGhq]:an<EW0IL:MK?_O5EgN392d_hi:LPJL?Rj\\@qG@
95fRPHg<gQ8^eSV8_>9G1>kMVm70Z6@[@><a]qT?Vh^Q^YLYHCL<ZQO38ZEm;f=]
1EF_U5d9J<qbd:1^kM^j>C<5nW9knJgaBjfoV@gVDd=K]T@PjVMWFPK5m>;CeBlO
eQ]^bpK2Wi3gji3jbJ?CiaK^<Cj^[5mU6F_>`_h;2E:gMcRg2VeD[HQPCHc_noC:
hACE1D=cSeUPHk7XKbkf@YFZga9lgGZF5PaAgWm0=jNTeHAOeaR2aYLfQh6mP;Hh
Tn<87nKff^f16I30mm[9e`3]aWCnq[6B[^ABY[e5:ANje5?RRCe\P9IPcMZi_QIF
e0I:1Vo[fX<E@77dGm7e=GMD4_R3P=fYm[a6WH33dlmM919jGg_P3ck:eO<\dflS
b`7\8a?:0Y8KVTAW>TVH1j`3`oJk2[Sb6g1EbJenO[<LX6U1E[[pJ6N=GbOadPAm
^k_WZ3_PhIUfc7N4T_lVA\S0a]ngQl[=MjeicZlGcXlIB=O6bJVDDg_ddebe]kTC
<RI`;8JQW[I56E;VA\BnU3\>c4mL5^92g]9J<Zi^BO80hOfA5>nhRBLFdEIEdF>c
mWLHi5WaRV6FgYq5f7QXBG=77Gc]bPUFf8@L2^NZFT>WT>K2<5Z@j0mOd`fI@Q=X
PBNJCLQCXCQZ72>YY2P1Gg\GXd1CJLDMjnPEaBF?:gkco;@`TK`:QKF2V77eKE]G
Yfg9bL?Nn^MnL<R5M2h1?RQ7OKOjFK]fXKgD^kkWgqMIZ[Y>1KfMmEBlmD8f?]Zj
?hia7g?MS1NMM[gCOF\ZlZ7V4;aFFkgCl16j[BDBGZ9>W]D6nK1Z`0_TR68bO80;
nDI<5`aFlj<ANDZmDTGOb4_l7O_GQF[GET\SaR6:HA;mccD=J5fJT9Dh=KNmV5\G
];4opjTG2o@gEEVCd7LA0h8B`@Z[glg]DYkm<YiRIjhkkEjPO^80Ca;P^Xo?TJYg
3032;@WV_J0VOB_3aOF9@mXk=K0P3[]g9Fj_lj_b740`=cXL[[D]PoP9KkQ:^485
nU_b051^]J:HaE8SQ?_UiB6eR?K<@7`p5kXo[_Z_Y?gVaQKGWZ]0?PRSV8KgWdh1
d]kCBjXjjN9Q30LA3_a:nD[CPC3<5DN1;<YTKlFMGR@VUl`2G3fOC1<932L]IKXL
LNCB`6LQAUnB7G9fHSg\J^Me1gDIBYBC=;gNAm1hTPLGfnGW5@EnEQVBZQqh>V9c
HOA>12L;_cl7WD:4h[:?1iHVC7T^PKOD;^p=DGmV1JOFRG99a4Ej\HfCQK>_PIjY
`80?@`Q@9;WY=E_V<KQ;BLF@\6lJ>R9cbE?3Kd6dhTS[bmml\FHK>:48lOknUgKe
1=i47\>31_AIZ@>3bXA60o9NAmd4^nTC1@>YnOTY2^>WWjice7OCFX:^Oo<d=p17
_W5HMSX`AM1YK?::QTIkMnC`00^W\^P:kj7ml^FdaY^V15YZaP:OGeQ8X_Z=3O1S
kMdWfHX=HkfM0Tf[U_2U2hG<I<6@Va:Q6mPDT8<cDC4P`njIJYG7llWBgbBU8YW3
j78JOV9AJ_p=i1G0Zj;BGMC_;Ef46<CgAo[XCbBoX5C2ChFF01N7F2lN\j:Y`T@V
i^iIB5H^l]<=VoXF:6N^MP8HGJog`OYnb^4LJcO`U8eI;UCf>[>g?:[SUOnGn61>
ATEBV1W9H07?nX?]b4Y3^EHXOW;q4@4mD8p6gW<[UkQ><ABR6Vd[R3^O42QZNgHL
^48pJeFg4SMW2JJ^7k>]GH4i6W@SSmoUmR?>K:=b1mpAkK34@@GD[=5=h8kh37Ik
AeW;5CBQR^Pl0MZ0Pqc9<j9X2i;iekOP7Ff1_XfAGoZR\4=8d^:8LZ`HPM`ola\[
bRTakEcD6@aWYiBV?KAF\@Z9f2]lp9K<G5edD@10jcS7J:CdP2FbP3?e\dRAViZM
VRol5ZO7V6aW@;N=^T8fJcP4=Reij>_8\6TpYZo0cLB$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZCRBN(Q, QB, D, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   reg  D_flag1,RB_flag1,SEL_flag1;
   wire D_flag,RB_flag,SEL_flag;
   output Q, QB;
   input D, TD, CK, SEL, RB;
   supply1 vcc;

   wire d_CK, d_D, d_RB, d_SEL, d_TD;

//Function Block
`protected
<]?>:SQV5DT^<@:Y86dj4?D[Soh<k2\;n[JOIdP5MN^qUKdUE9_0Tb_j<2@;=2TJ
=JC=E`A40[gqR9FDYSDUEe;RMRBen0?fpiTCK6kp<25enNSDVZ[G]FgE;C\=ZcDR
g7Z[0d5q`:THm:f>gV`\BNhKM2[Am`[J9C`HG9]NT^p0WCV8mhB?8k5NW8]XZ525
2jOCY]@kmGUm<qn<4]W6S[H=h;Ih;C:Q\FTfALBVB_R:_giWf1pYPAEm9^amflEf
IaST3;CiM=_3nqm_HKho2PW`3\O\WWeHG2K0BU?NEph0OWhndI2Uf1LkkdlIJYdg
?@`_oW^2joDf_g>`Gf_C<M1IM>YfCR]OS==kB\T;lWFjWF?;BhMfP\p4YHKo=lD_
Kb_i^bPOPAa:84@nhJTlfUlH\J]8C]MSXE:P]U8T9E[_h87d1Wjp`0W[HgamKGgR
<g^A4V^FAd11ThHNRRMSm4<TAliql:J7kTSUCMNKUm6h?LVnPLbBPLEi0\3d_X2M
@^kG<WQ2U_l\PUKbm45kZEkp8GAhLLZjn_D7^`VXJ3?=Jg`kZEcK[_619mp3;NdR
gJcB8bo6ZnZW_1Q9W4Z4MMN<WUOe8dHP5iqcXI37jb8:Z^@<EkXJgeQ=5ASCS5@o
=D0FXp`]_DD?_ZSSD1:V9j@kWF0?J;0N?FQ9J5i_Kdp`W`>5QUJZWX<<DY83T_G6
Inhdc\FpXROD?Zlp\[?^HY76EgUi>Q=?;29?^9P4L?396C8bh0BNdOXnRRZbimFF
l?OQ;VZLSG>pGmnW<>baKj0;Qh;?dOiQLSL_B\?o1hnqj:4WmXDpJ\:\\VXYW\RG
3WOUL>K@YdhkQcUB[ibpO]>J5hJqmfL5hYGfc?<LR2cG4hg>JO0EcR8R]ZUNmf1B
>igdA;cCm1jR6E5E78037ZqLlC^=iA?BUiX=:h98fbJVcT:aCep[Tjek7;qX=RD8
F8l2gPKlE=CD_8Y1[2lEG75?JF7>]l@:gZRD`ea1_RGR]NJkPlH^Mp@lah`=K1E?
IgW\4h:5hEW4Q3l@6b4K?Dq1ZlQ\KXqIB9@0[;N<ecY_npXSH4P]Sd9f2TkFlX1N
2WfLg8djiI>RhipnCR?ZaRph>PjYKcEOi?kR@\8Sd6E4a@aeTfVjPqNFbRZf>pK9
[ha2WIZgSM2QT8:E6<e1Q=`]mFpA^eeFJ01E75^ck?l\UQihhD?J;7akgolHdp>V
FX5Lap8?_dP0m23M8V9FLGWfggE`E_Xc1p?HFGT7OaD^Ca2kD2PHSm<fm?[_Z_]`
Fje`q=\K3Zl=qkB3=[N;p85@McEBlc04T>XVVqDbO:BSqnVIX<>DY^Y98EMacTcR
^f26@?EVF6ih3eJn:@eFOCU^lkd@nL4^n4EENWmUh36PjT9P3bj;SLOIXUbFABGV
9@bTM@14PFQ7\L2=Kg`[F=[gSp>jR4J`49gSW^b\U[MEF27`>ROGbLSP935GSRXn
3E2QcFJkgFFA46U7J^DZVEBUl8C^b;cOFS3a^h@1k>:O<9j=0k]23A655DLHT783
[iCToXcopD>Yk`YqGaid\\UHKWUS@9NE_PEWU;95ENbW5m?lo\<k1Wpg@6f>F6f5
Yoo\`acBT:MdOlVQmVijlZa7?XqDNW?LXbA_]eojn[_m6LF=AgaON;L6LA=fN7XB
j_qi`RGL[HY22S_MIjDgnR74kL25V9DEfWc9cJlpm1:CdVZZ`GPf`fddllBXD6Ah
0?Dk:CGAB^]g8<27pefH5=o;2;90EeHenHGd[SN^1IFOHXe:kqm76=H1VbB^Kl<_
gSPlWo`abMkP@l13LRCTFU_Cp?IH:L;92jFOCQb<=Slo4o5616`::ni_HI5Fhe:?
qPj4bG:VM72bMO697onZdMYXc;0?UhjYZQZA]p27?BjnkOK3PS9@[2HcREnOMg^@
EHG;@lG;7E]j14OehQWHQIPKEmmWcAd2X;>KZUElh\W5f4@A1<ROG6N8jUMejW;j
TZLTEQeMFAn>=hoR9gTEB:hm8Tk;nY]lP0FC1=A_Qhj^YUO3bQ4Pp@=a@n[hhb1D
;cl<K1l?Hm1mZD?TRY@3WJ8k@_i_WB?Q60`ZeeTk:PYL4;61;TJ`Pb\C5UgYi;ld
M]VZ?n`EjKMiH9YUd8WnbKDFi1OnV8f[VBY6BiSkU[Bo:;OdC8l9ieEQ>\k48f14
dR1pLh_\F?hZ5j:=7dQCUj08=7S9\^]4\JG[P`Lna`;8Eka6:O_U^Wn=m0<jBIIO
]a61LG3fXfN?>ncKaS3knE1mh8W?1B40f[M2l?B5K8m3Ui@B@ZCO2VCgT2ZP9>AA
c1enB8CmmCY=bcU>J8_D2Wq6YY:XU\Ye4g5e:309383SFB7@DejoeQLXO6<TB^j0
@NI^5A4[MT^@2=LE<H42_eN6Di?F?4V>e=R;8:`HdZ8VRj:N5V0c]724V51[WD^d
2\HSKVRYLE7@KmA4B3>G8mS6bkmWXXI8EbI3IW<ALomoCpU0>`lH7E16jjjoVLEo
Jjk\_EP@m7@=8AZ]BC0_eY`e;9kfMemjhS1DmP@LA_hSI;]FmJAiG^;4I^fgNlDL
iNaHm6F0;ST]R9VAA^odPijTMNmR\m>cG]dALF\e9S>?5S7GcR1QJClSa;172emU
@9TWI\Lnn93KpN3\KI5WhoNV_SBN\R`hXl?>6XO]fYOoE;:JRp^J8ND1^`<?5f6e
X1a3Racg06S\l:P<NBCTOijo^f7dW4a1=H6j5ng3e=hK5XWSDB7:HS1n5a;`a<M`
<Oa;?Li1J_M8gCCL]ed2]?]:d:UnG\R2>9;999anecfgmJO3IbT44W__\@BZ`XYe
AJH2ieW0Y6f\q5<^H:lo[^Nh1\J]B5^T5i;0^0jF8CIiUJTH[:PE80e7m]0GXP>C
lij20[m7jHnR\74iMVJnSlXaZI@d\\>3nFDPXRdJ78HIK6cU>SU\YFhj]aamT7:K
>m?If`jRHkWdZYh?L]O:R8a7cIlYI5T@=p@jFBW00UKVa1aRhQ<?I7E_j[OYH:8^
>hh9^RQ6n8^\YPMGQe]7MhX6U]<BSXNc@gk2]]Rj`0WAJ]j1A[_K=I8if\Jc?hVg
B`g>M32dUG;OM@I<A@hdL6E=aS\6ho3Zj05BQ[=TCNo6G2V:=WOT^HpUQL7_WqDJ
8S<]deE40DO>:X6ge@9WNYL@^AAN]kkElKURpCc6Od>c[`^DbOR:DVg?HM;@?:BU
\^4bY=]HEQlq]IH]cYW90lKio`fHiQ8R39aL7EP5Z3TKOJUi;YJ6U7TZJmpBkbY]
1oM_cmYH5[Iniag\E:kcjFo6kW<=Mh1LC99T:nG56eSXC51RJ@PheoEjPXVhjF<[
DQY;Op4?jXJ^NO^o?`LHaGgK@PDMI@1mK88?T9`MYmmN\BRCIS?:>iW2UH84T19Y
o5;GVEoJ`Wh7pDdjG9h8$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZN(Q, QB, D, TD, CK, SEL);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, TD, SEL;
   supply1 vcc;

   wire d_CK, d_D, d_SEL, d_TD;

//Function Block
`protected
SM9IGSQd5DT^<jU`=HMZQYP@bLcJgoo2^cMfYG<\lSLBF>l5We<f4miIqY0aOgeM
n\i@ojSZXBKhC@O?Al5@kTY:c=J]aK4=aPi9k3B]qX`PS>Re^dB6^_`8Z_7XK^6>
]k:q>gUgB1pgbZlMJ3Fihf_fH5_O3oEiHLR7^qHQ:7>flmY;OS1Yh0\Wk5@kS<E_
7q4Bmc8<U<h_f7SLbN<^;D>AW5TG\oU?YABG:gmd7RG4jSXe]WE^SE4UJ8m=gcGD
B0J1QKNTbdLmSZq=nIcDD>Il:TNS\L[q=@BHA;8EoM]2U[I;6C_]klT9fkj7@jJC
E]3Bh40\V6]aeE`I6]Nfi:>]QN2;p5V7gTggpP\oZBCq\`l`KXFLkdX]9<lNcQ4U
]7f:g1No2E><XdmW8K3bh?PSl`TQ1=6a?O`U];4nMdL\B`Ko5Eb5J`G_Q:;`hKo9
4UeHTV;JbPMc:m[8eBla8;Z@qAV_ONoJ4nEL><_7oh_elT65[:5ON8mRGEEDf3O<
GLH4=eOGCTLg^Y>VnL7K3GCg<I>MCH5kREIaRY:HK:j;U5UWLhFVD@MI3H7HVBF2
`ba@_gaqWlb@DC_:Q8\@=CYJp`8>?ZXpNO?Ieg;;2[Ko06<>=7hcS;dJ=NeJZ3iE
D^nCGAqnakNb4F;lQ\<_H4_4RC7??VFDHn:I@K\XhTp7S3440Roib<[^4bJkCNHg
;OgJQVmA==;Qb=HOHQapA6FjEFj_a95I1Y=E>Vkn8QS88DK8?@T1kVmnWDpOcbgA
d7Z5HB:gjZkPmo<7If=OMnECV_i2nK^iEipSi>=N>C8CK?CB;Ha<2fe;WWUB2fRM
ogH5S?\p5Lc`li7_KJJ_FddL2b6Iecp5RCVla`dXL=4LhQJEhfdi5fKKcbcifl3k
7T0JC9PLYAnYDLl^jldhBG=NKjj8@SWP1L^?Q4@Kk2NHh50K[Kg_LANfmZ@WARlQ
5S<Mh`FW\calG\Ao?gBjE;EZC7O87?09\0Vd1EOVRBp_Wfb^VjTRLdk_0jW]hJRA
PO0=7bU0WoTjj29EjY60>8Rb`\ln^mQ1l7bE4RFM`=ek@UHI]IKWoH=lDVb01OaR
96mgAT[EEN6ho_Gg94;HX^R11S;oF=keSDT]TE_BART>dRl0\=afSSqMTkhCM00E
2NnFaEj:l>B=;;c0GV9i<2UPGhZonZ039bPE`=?hGbam\35a<:M_c:OWcZT:P=C>
K^TOA[?l\TI7_okoP@m=gFZ2[`ZiV8l>dD;k4Gk3I8=?1E^m9USbOSIVfIj_NMCh
<qYlGQo\9a>;gbXLa@dG<9CaE@[_k7U\G@]VJ_heYVh7E_k?6CH@[iQXB=HJ>c1G
oh3>7^4MY:j]3h5V7bGD5M`5A@:VSRjPRC5:H;BAb5NY7?LEIKQA;3Hl8mhimd^K
DDb>3HbR9]]1p;K6\mPZnkG38@iF?]lcEemXb9h;BHZaSD6;8[[I_S]`Rdg6C<LP
O8ZSlJGFLFiDG;YK\Yk9^=8B3hTIE_?KC=]R>AjF[Y0\KdQEVVRReb2jQWLQ_YMX
>e4;4DBnUiXc8YZH@kKQ^M]`X?UMMqE[KMkdTd`]dB>Nac[5N\^[ETIo9eaS7LZ8
^RGIpdaa9C2:Q:X;UYR^cP?a2;gGj>Q:gHA8f5T>F5CS>1L7kX3JT25Io:lc>R9j
R1Rb0d2a>T[PP>T?GdmVVH\7KanOZ2RPHNL]d2BJQR;k^6[^46\4SjgSkl8=X?nB
;ReBhPYU99?;IJ4>Cjg`Cp36W\mZpUGGhKk]>EKOk9:[SHgeT55SNT1;Jf3XgYYn
:oJqAZjkYj?`NfaJmn2QV>l2UK2BhK]Ua_K2fohjZWqA2g70iOK1NjPllAGF7bgD
SM7jE?:N407ccXH=Xi>]eN9_LdRfo0c<]ba;b[4Xd]J;1Jf^]o0Dlp69:JiZF^RA
[HCiikEBRW88fJc\QBcf=]C00RQO@E]B\RV_o9S[eRNPUQi]On@=[DV>n]5LS]7\
qAMT[GX3$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZP(Q, QB, D, TD, CK, SEL);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, TD, SEL;
   supply1 vcc;

   wire d_CK, d_D, d_SEL, d_TD;

//Function Block
`protected
:kSV0SQV5DT^<Z6h]XjP5?L;ZkP\ea1ge3LQ=l]lZlin\I>l]I8EHPC;Z;\Ga<EH
^aFI7ApM7fing^7ifjHWZFkORhH\]TA0[LQpOLSD09f?LJUU]f@IIXKhFPPW0>@i
4@W3K>Vnf8B:LGOf13oa5a3pVKE0FLpO[bV__bTLOCL:U926CTi9`a<a^pVYAVI^
4PAal2n4cEUS;W`E62?mMq5ABO5T1jDQ3ANj?8;TE^71n`eV@0m3MlUcDFlhl1Wb
97fN<>q[o4a=`@Y9>MJO@1AT?V4c>lITJM2S[KY[F\dV>`ClUYdP<k:m]EFMJ[cJ
J39PW6b5U[80XeAjdG2poE]38YM=CcnW?]A2<]R^FY6_FT<CX34K2hW@Y7SWcWNO
_2UQGZlMn4goF;oApcEGCcZapRV_4X<3O0_GMf97YRb4p3JkXH:pVi2j`3L4T3I@
2[DikgK?<I9CB8OHm@5c1QC1B`PR_EX`0EGKjF6DBhb\?Zh:HNVSeIM?m6;^>cb?
Pj<oZIj7RWONJTgBGR=E3W3XoLb?cS@KqlVS\H3AZ:J4]<lMlMH6OmZja1nV2=;K
XK5;Eee;Y=DK>ef>UJ@R6cFfQOd=^e012m?=CV<3kL6CoCX=h\O^md2ajK3Q[KS@
:VokA5O\2]n:KKepGE0gGepgW4L1S7CGche@SlH0]K;Ui5`<IG7\lEXDcFi=0q\M
1C;0cW:FE^NR6;?T[[_EWbe;7AcDA0EE>pBOE>GYmRamH>ODTp6QS16kThlVj`1M
7l9H6oZ5fLH7;UVA1ATmVdg4B^qN5F2<e:_YE@X`h3`3K4Lj5Ofc7Ue@^gIBVl7\
SqbL6NjFLg1E2Kd6?@JAU>dNaSTh`?bmH8kkdHmBnq`SZcTfj\1YE>k6iaZX9TP6
5IM`qhc`;7i<`CV6^X?JZHj3n>6@mYfl^l1^lTG2?p60D@=TK83S<H[;187RlN>5
[UCk\Zao;C6D_16bX9Q@30A^[l[A>9:L5Z7:7O;JS6]DkXeocJ^U[k0O72e=e5TX
Rb=<7Bke\:Tj3HM?hc[85?JT8@5O6<6kkSl@cVUmaJ?c3_b;eWm@gpT4Z]>Qc26B
FYbFH^oV>ad<FRJ;_3`LafHTFC2GORXBLIBc?L>@j=DnTndA8Fi;OYMRQkJ=2KGb
iD;QO1SoE^i2SWa3\73TKjGbWWBm3iQ[BmV5`]o94@??<AX]1TL2b_a<M1Td@De@
dqX]RKL92XLYNcS2k`2cnCH5c:hhl[HhTi9^j4:C5B^4>iKo48`obfX_eP6UniYW
__JQb7e6R]2lVF@kU[n1;DLkcJNU`AADn1`IA<WBPNL;?RR`?hG_@F2jlWB7]jah
f\8HGbC9gec_pmEfmPh29D?=OcCaTRX;X?aPDH_TA0<ZoMI;fO3CgXZCHZF9`LXB
XfiHEm`MD6lB?Obq45=1niGR?XRWJFHT^>LFoK;7OOnnIa<IY>l]JmI[<gLoXm=6
iKH_8EHI3JlWXc7J?`PB<n`Jnca_Mif7kDm4Hk>SOBcJJV9UedJO5Cf2_KQTB[M[
VJ^TCNH:Ig6BhJWaI9L1j<2aanqU6=RQCJZdH[l0DWZjXWiE9GR7GQid_^MBiVIl
>7l9Qa>KDPg2a9>KbV=A4R2M:8hU0ALoFC3^gBM0ikDcNMIKSii7BBH]cOQ>X5oa
Pk1iXgEl7G`2dIUcXa0Yee5B_fZ79L0Q]WgWmh;mog9p0b0C[5BDW>JQYVISeT:e
Ai_36cH7O5fd[=a_SCjC:T0Bl5lCgBUX`=QE3LM6[mfl<7??3:d>0_5bOmTQLbg9
3I0@:BY\1j`>BEM0Z?YiJL?:kXS]\I@U:Wm04oF:]?InYZ]Y<j;b3KkJh9a8GeVl
q3bF:Uap[Nh0Rf17Q[WjW;Vg:JmXXPS1U`A]UM45?\nDUPp8m]fcnok0\B\Nf@3<
BGcF0F3`kgkSnCWjU9^gJ6lQc3nqF3aA4W4S9o<?\Ae^3KDd6CLbL[LlhFCRSo=]
f9p^NRomdNJ7CkQIU?I^]chH<J[0\1CbhJZX0QnPOL@29j\ZLPdIFmoN3T`k=[WZ
VUJk\coXCR_MEp`C`iC@TWdV^3\c>Z9XWgE<c;nOd715niZ]NHMoEn8oR]<a>@Q\
D[41d;Ho6GO?6;f@ij9eqBMn3?YS$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZRBN(Q, QB, D, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, TD, RB, SEL;
   supply1 vcc;
   reg D_flag;
   wire D_flag1;
   wire d_CK, d_D, d_SEL, d_TD;
   wire d_RB;

//Function Block
`protected
PCYMNSQd5DT^<kNhL^OdYie9pR@QV4lVDZP[m]8BdiFV>1LF`\DqUNA@1l>iVZi]
>;^GXjUhg<e0bL@SkE4oCAOn1A_K2m:Wg79[``ZY2o^i_HTB^27q78S@D2p;Y0d4
4WV:gBn?QBTCkJ89ND[8_>lj:ZFbo<^pD8:Gdj0>@K`80JV^dPEh91fk>?qBE2og
ccML2[1<bMaL`NKLaN[k^MqLnQ7<L3LXA[9gA=5AdZci_7N7UbX54fdLWC8QLHO3
SVlf1aNKBlKnbNOAGMXAf0^iU\ICHQ[2FT2R0q]mRjg;g3PAVI3]b@P@3V]W\G0A
Qoj;[`DM;^bT4=n9EUBcjio`Hh1@eU?Gbq\X[J;Q[ieN=naYTT]<?fbX9d^fjL5^
`_pTJiNY`Xl>=7ME21mhb^0GBQFcOal\H;1j3JiKhpj9i1P\@pmjY79?Ra;jdIY3
_JJK2`:8G2G\Z;o]^pCml7ZBkNBDnKF>TYb8dhCZQYXTBYcQ9p=8I_N8U@I<?mRI
fgaHLA2_4Rj6p<f_J:b7p;P=b^KYlQVQM\oReBIG9c1Pg=3gpDYdfaG6p=3=bFU`
q3igX:`qaPI@CL@8^g>4OF9G<cc7Zh>a?K1eV08bb2I_WIHhd_N]fhqiBK108Rf:
gH<9ODGKaAGTJDf1cWn2A\]JNF>J8GaNDh:mW=^5a07HSKM\9`^;`7TaaY2I`bL;
\]oXY\g2G9OYe_1RCL0oYaofiAgO^aJ=T9AqWiDG4Mi2oSaWn>27g3:CB8oZaKmj
7D@0:M6A@WH1>2BMcaa29`e_2m\9oF[6GY24DT::<`gWRcZF5bUEV;oOY5FEC1C=
1e8Fg09O;6JNb4;[Fkqc^]QJHgo1PAPR5\;fm4im>?Fi46KFZ=2>>7g]3mfPH[0`
Al2eOJ^am__T<D5gE13cZ]QJi^N?1MbAGEI73Y34R_ElYJI\VYInMj[qY5SODZnN
RnCEFPM`i0:mOXK:U5H@LhJKU6DL7=F3pDJbFb_JHKAhh\m7J>9MU2agGKEU7eoj
[;\:YZIZR?SRF@6dY>QWJo5Hi^abKoDehG1o=>kAPCXaN\m7`6hFL1C>19maPmCD
Ej^J5<H?DD1qa<<7d^p1B=XPGBAcVS=HQVWGNTF7aT\R5GAnfk@WlL8qbDPY47K[
ThKmf4JTooO36R0:hofVX<@9@l2pa2]eiVV6NT5\HP4j>4k;K?aRHTc8Yi?oi5bj
\Kiq2AdL15eAYjaAR1T:SI:73cBV0;b6Z_QI]0Xk6dp:fon^QZF4hG9i0L;M;1Cf
FS8T\YY\oEQL:W:f<p5C:U<V8@:H>:i5TVMlB8kKd=XRLG4V_L[TmWpo4RcDU]hU
CGIHmEUn;bVi8SW3g96oeNiKWOKiA]B1WQ=I:H[<8T@h3;SI>]bFm6Qi8aQIQP:\
?d>jf1II\JE6ePe>DKB?TbJ5I`MTBTSc0H3cG_Y4>ika0ih[aBei95eQk\OIZ06M
libb9W0<2aphjHJMBSfFobPFPJGE<L>AL6qX^RhO`B=<cC>C=kl`DEOSWVMGebn2
c844oYn00gHW]W?k7SQ;@dF<V]aaYZj@FB@FJRP4P:K`B^EV7jd;ElbJY9a_KQR0
<0]J]]X:IUNbc3;UDehmX2>P5WO=GW0GAW<NL3IST1L;ag1[QW]@kEp[fXS^loOA
i?XQ0dKU91oUFm]]AJF9;90ASjl;e?`a[<4?R?\eU2bm>j2<dgaV8QGBobj`KAgB
Wn1i5[LH?:\RQAjH9T]02icDfS\]H7ch1VRK\=N[;UDY9@C7:jjMLbF>`T6DcBcF
AS_YYYMAdpG?]5Nnbl@Lcn@OJZIWNAKn`N[ONE_Ik=_nUfXUV_[RfO2TY6l3leD9
5jTg8nU24FHla8diVbVHXlS[PeJ0?Q8DAZZ;H39=lC]hLSRMJ5kIcO_KeZWgogjG
5Am<`O`]d5a:];AaQ_6K^21`BlWkq2B6fYk]c4a<lK_8eVQ]>X?dKmK>mL;d3Mk<
B3HIWA^XZCb`]\T0YkSIGR:k;6jTS2:mBV2?J@GP911HmNe[L_h:]A3<I?[MnH20
61`5;fD<j\XJ@CQ`DO?PKnh5_\DX7]4IV\KQjP?O[gUj=Q84CB:U9q^8L6Uo[A90
_mPcJTQ9<NF:d\NaCb1BnO4B]\@nY^H_NoSo72i=@C\oa>=0^NlMcoNf;P2=C14>
L]P1W\C]GA2ha<c3HP:gjP1bT?ilm8FaASX]M><OHSnN9]?^iSIOJ52JX3G8XS\[
oB_1@HjXPgdc@d94Jgq;leKQGq_j^`9dX?_]\b53b9CUe1oRnI5\l`kiCSFlcXeg
kn=nq?j;Q4Do7d@EIaWTdf^GlOKQ;GT]l5DVO\n8\6W`SaapRShofcES5fVjhTG?
oGFT<c?CeQj7:=4abFn2kQQjNN:PbBA4Ze6QbP49K;hol^>7OV[FD@?H<aXj4D5c
eNBHO`f71mBR=Yb2FWg`>QJMI52A[6BKj3c`>IOM^XQXX@OL2b:@>m>Dp=cB`Z8T
DP9MmVPf[7=\QPY>LdeITZM_Vaegq]>V^S4qd^9hKjBZ^M]T]W>TlDC@7kiHOf\k
gT2@P^0;q]?JLhleHLnmk9;R?EB=FJAg=G]289KgbKLEQ0dpcO>L]@8TaRQhT[\o
NoVcLlA:IO67[_C2mPmO47qH4ij>Yc^?=[?gjb]fj@Fnm^9=@S2dlUJImHh5:ffc
VEf4F>ij;\?3TM16kfVYAHdRi0]3jkJ5`qgg@PGM2?J4@2_Y7RgDS57<_^U4V;UU
NC[JU342SaH>N2n5Vcm<V<7gmC6^b1aADEc`Rmi6J_:?q7BneeVglY;OiPBIE]Y8
mR6Ba[RQfXmE=Nn^Z1CMXMZT5f1gQ7iN1jZl`a<HeKno_JYP<;_qcmYHig=8=7`B
HjnBgE:<o`T:c5=K5_:YOnSph_LA;N]$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZRBP(Q, QB, D, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, TD, RB, SEL;
   supply1 vcc;
   reg D_flag;
   wire D_flag1;
   wire d_CK, d_D, d_SEL, d_TD;
   wire d_RB;

//Function Block
`protected
f;gVESQH5DT^<FT1bBCBok]`PIORDVj@3F3]KPq>ZGM??BRaKFh[Z5ej7oCMU771
1g@gk`B3\5FL>LqT7^BVa3Ej>MBD>;lIGAQc_TZci_?aaK1FnH;QVe9q]hc>S4qn
CYF@ehChAEHmH2WlMe6M?hDUd^iE;\SJfQ@qi?OF2WjCFEaAJjn[8F;:WT4KGQqd
Y>_YUK3\F5Rc6cmXMRh7f\YGe=qFQk@JD^[O_R0i9<6j9GiD<I3lREEXCh\?OSeG
oaDAe`3271NjAORP0<8b?8NBSb9fE:3No:jh1FAK?qeOBI0hUl;@I:mQNm<Wi5[9
Z0oKgq6V?;8Je2HQ<N>X@aRJGR;[Y?aUGL_?fPbaHi9TF5ZH4kG>h2@h^0bO6K=V
=qU8LJMD=cEdWQHX<leL9O<\9<M_C9Pj0ipK5;>gIJYGKYDf@F;^B=_;KLV5c[bX
O6B7k0`?1qg?W6_i0q[YI;U94Q;V3\CWEq7G9W3fQCM78ThNWFll6VGML07:XNYk
9pdK::jmaVZUh_i>Vnl?jh0J3Ponp7YLQE``qM9JcUBh>dUDlg2`RSeHTIII>=n8
pbb`6A^[p\K?0=W2qAOL:JH3C[M<I3T?b]X<TocJ:C>g`PCKKhZ5oihM?Qm5l`S5
q_E@Y`mplT<6VZef]1a\9k1h3Q\I@ef^RZJ8gYe[^PV@[?``?]YJ6BW[Q6eL0`;j
m;IZVDDn^QhBF5S6oGMgNi2LZ@cmDL>nZ3:H:cD<4[EP9>ZE^@MQp0bGRD_];g9`
B7JX0jX[FboZGK=T]fS_TLbeXRl2:EZfNFk;kBKNWm64oMX<>m>aZH]PI>k4jS8\
Diec^KIOmJ>d`Ncc_`L\FX28KFWfLahmAR2qC[cWUMm2EZJG8QV6DX[Q?I@O\g3e
fiU=F<IS2HmXcI0:gd5;H]AMe[8QFBXDiU8nC\c6UeGV4;83AKkRjiEMPn]m84]8
ATE?ZZE@qCbihO>B`>f1NiZ8Z9o5>ZDh9]Y5c1;IS6Jb;G7:oJehE[E1N[JoeDdW
eYXkel20IELqC4fZaa;5eMhDQI0MMJ7CXCZ\FlP7^SOG7[MY9gJT1MUDoNNgc26\
:5QW:F0Lfom\ZoM13ckA]n^SmImMNN<1eRfiNk4X<FC3^T<YYbWJPdp=VMQ8`pW6
^9L>WJh5oTeTiVC2L4>T5iB[OgNShB\4m[ql=EGkAi1=eDb2gl=1B^bUaAV0B2M1
A8G2Q^q^Hf>eV:J=jcRGK_3]93o24?b8MJZ]Xgo:;6[2m2qEX5kP\F\T7S<__Ij3
SimRlQdNlT<1mNU<>4l=Cq[kSN30f5=@0>G=mncMhCPJHic]En4OJDE20A;nq]N5
DMbU@Rkc1mF4BjOO`noIZX6_H>4U>2LF>p?@kdB\2OQbH<GQYZe]93Q?f_hCXVYG
9R=Da10G^AN`ihDXMEW5eX0<eT<SB:c;PF?l_FfVCPA`f@XnLgNI5BJUnLY5kT7`
5Xj_BeSMFIEoiL_;l>3=P:@OdZ`_cSglAf9<X>Za=9[IPBK\da?iLpNeFX2f=mB>
\6A4c@\nJY?ngOqnU5:gUGMW2m]^HZ[VcEjdF_GnYhgPoX\>dU^96@[\L01Z`963
R=5?iH3@M3N=nDOfLamTVdk_RO;G4G`>`iH6g>Q>ENP03B0Y@_EQ^QM3N6m8d`>J
>a9D^LUcE1GmO24[0c>Bi0<<Gd?ClPdbhPp@i>kS6bR9H\Qk<;in>;NG1ROB=KMA
LBm`:QG`E3RXRa4kfOk]YY1b\LaCn5RS:3n[hOT7T;GlRVPF:?J?W]OWmIaUJS;O
NYb;M\NnePgoM_JVfR`COS^CaU]5o9HOX3Rf1BYKWBP]]`V<Z>NBmqNKYTG78=k4
3:m8c_=@\o:L\YcUcZQhe1g5W`iYTN>1gA0OY1f\0KUk`Q9hl^jQoR64S>QI66AB
BTH5a4>WgL3I9L1J=fk7H3A<kEn@9gV7^03ei9ZTh_?5EoU7jfWRhQX=I_9MdO2?
N;lUD8@np?2^5oJ\ZOgXnY=X9iH:_^Yj16hkZklJUD\Y:HG2;adA0lU;0VC`BY2@
;YhKPdT@J?b]=jNk4M2J[U>mQUF_mX=Nb=N:>bo;CE[gS8Lb7DPk=L4D4nf>IbH>
=_WZ_5=cKg]G26gAJ1R4Y9^n6b[ZWgUF6pnS6n?\SC9dSh_UnEc0=;Y3ThJCfGUM
S9joc0SK0Q=h:G>_bQaVB@6[LITK3I0Y76l>L^XXAUkl?fo0UX<BHYdE2D[1cZ;2
PAZN@X^?XMAI\RC=Ag^Gh2SiAGZ1B[4nUPJ`D9<PKkSI7XkLcH6=o=mSnPg=Teqm
Flf1Z\YB`4;[<CV0S8Xba4@g8<hMDARdbGH=Po=\\jC<lmPAW90_GL]XTi^FHmbK
Vd2WYSOpY9Z^;Apgn^3QWdn[a]1hX\m>anU[2_ERF9g9j_5U35TZN5]97qZWBBWH
7P@OiXKYF?f<QAkUEDPghN^4bQ42a:nTiKX7q0TgQIA\GQ>g]G\0\`]=n^bG^DH0
]0UFC07dPhRaPOiANKmjO>C3ebAnRU0IELlCSkQX\PaSCkRcGViScMZ>=9^]g:W0
89IbDhae?JQ4f2fhXj=I]PZ9TD]^d]A>bL73Nd7N73N?AqjZEnemqoP1U\:0OnH9
;Y0:T1UQV;c9\8;IJ5jl;SBIBqM0ZdIb6dJCV_^bWU[g5Q;=9Lmg[KkS2U9oODTP
qQO_::ncJ3jg2fk:k5liTk?I24m07RVL]R`oaOIqbhMg=:O\D`F1`<>nBcVba2kU
8?D\EU8bMAJ82`T67Dci8?aVIbZS0]1km27INkQp=Z5Ik5onIY=;271PeVEg[5l[
e?F0M7S?]<J:GSf\?0O8[DcZmClBYAn6UEGkB58`@Mg>EEF?g1p]R8Ca]7177C9d
OR5jGZa1[PKY^EVOQ?J=EXgKK2dFnEmHbT>X^QjJ8[A0Zik<=^`<aiJ6OeA31p6g
<Ig5U<RjH;fNin4Eh1;044Slai\h:HccL3Whh8<<jOb==_<MXhLlT]a_JJaFh=`n
[STH=TdRq:<^C8?9$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZRBS(Q, QB, D, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, TD, RB, SEL;
   supply1 vcc;
   reg D_flag;
   wire D_flag1;
   wire d_CK, d_D, d_SEL, d_TD;
   wire d_RB;

//Function Block
`protected
IOj0SSQ:5DT^<4kYHi009kDMVh9E1]^_c:UAIi?_K1BZ>YV;@hipYOBbb?[I95k0
SYG:hZc9IMe\g;hnlNVMG8iV[fBHS\mqQg6W?EFnOoLe^FhC40MPB[ald8XdO5l7
q3X>f91q>H3MbM8k?Ei>J=NTjiIS1PV1NBU;B<lC@`jHpkL3RnZmC[0b=3d8_EmK
[72[_Y@pVB\8WHU:3FPbBPeOj6F:Gm7D:Qop=Cc<O^kMeWABhRC27m9XLgOGUN`^
pQi:I[kQ=dkWoJ@0[nQ03emn?B9iYJk1_`^Ja2Y@W8^2f]dAKT1g3Rge4aNDI_3I
L@V`:Uh`mH@@?=[pX8^[TX0g`N4J49L<_ldiUCONA^Rb]lf6IF1B>GngelmHEOB8
RUS4jmn_gYZqEKo6_WZgbnV`V?VG_M50\oF9F;m8k@6:pNfGeJfIaZ6jOSg<J<hf
Wj_[QJF8G<3Q<4AMU@9p=J3A6^bpbDc8f@O<C2?C3jXTE8c[D[eX2GFf<@[pO6Md
N:Z6l:`Q`@FURdFWJO[=M:pEGnc[XCp5`Q\ZT2LK>cW=Xe1?0bAD;^g9AOq6`kZ]
Qo3<NNKNa]GLKg2hb<2F]RKXOD6G]=QGFY>91RLmgao6kjlUYdhGfM`p4KbFS\:p
8;I4UDKq9\4IVNpJ\@O495l\88RH6haf[lX]<JWGERo=LKIM1m0ZbaZ9gDk1GRHO
d[eoXOn<mk^nE[T]AB[iS\FdUA:m3`EGMg3SgH4WmEnf5NCAD7bImj?TPZ8pOSXa
A6AKL3ANTY3E]U]i4H`1\CS:3XV4=PcXDFL6j<Mj`k]Pfgc4CC72fl>1i3D46dI0
_>X]8Pmiio4eXP[MoD]QUbZTOWI^HX5Gj_[^<O^CeMqX=klY[_E:^nEb^k_>]83`
Sck93JelJYcjCfYce3^<o:SPN;_==RoV<RClaDoSNB^XeklYAkCO7VPWeND?4mMl
?1g>XQRSc?@LW[=paOe>iN0;hmmK@jS@7aPli3=^fo>3VYU<mHm<Of?GEIL0E15_
UYNhFA;K2X`SOl3UIZT>AED2Qog^ojVUOC5T89>P@m]8J:[6BEW`UY=Z6^pGAC66
^pT`BBH[OoVb;Ch5YSUkno\CK9\8>OWI210CodqcF8VkcA9eQPgRn[Kg_CamAYaP
1T`iJJL33b^M4G>B8hME2;pEAnc3=b2@f_]?\N>eWNENP>EnfckWNFXf62p_Y_6E
dGRE_2QhkUbRXSoDBRRJU`HNafZ3\IeWG[pA<=kfo>3VYU<KEmCkj]Cd=lPM71E?
iJgeicg:Cqb9mg2?]25eY[^dSoGmERG@>Uj_gf0d3J]K>3Glp9>6ZJ4@g2[<EB^Y
Uk;acJkmDg?D5\^KDIUK1qlGEdTLeJ?T\OkCnmb>H;qW:8[AhfdK8j:]H_UE;]3W
<kS7ge]mJ3``Dfl?j82AbUaO^7>9;Kkk9mYjB3MMedNnh5OcbC]D^2]NOABoKEW\
X3Q08k?AF0VC]bV[JCj;>mLj8M9NdISeQGc?lU>X]M[:3FYVl4MoKoZP71oj_Tpl
Xe18K>3dG06Jj3BLIem6D0M@T?MZ?^>VDXSEiaTff_G:WPOnm3XBjfUV;MNIA\aG
KLYZALkcmAj[X\macEPB:OfMA\nWe3Ac\@heh]Ije^YgI8oe1O7R:SYi`382DYNb
mQA0oRdVcUDO9Nca93qX\9eBb__0C=@1=1hP\HgC4Sd07Z>_==i9OcRa9AR5B7?:
<n]YXigdQmPFUhl@0a99J2a@\3Eeo>LbJbS[7RM:KTUIlYooRFU=74B3Uk\eXFRI
XB]4o=bcVN>:8`NIOf8MQQ5MEI9]TOVeGL:;Hpj]SABa[Z6Uj]^kMP1TmIXCa]PC
k0=SS`f2\\991@l;LE@o>`=U=i8KfIFd_9mmb9gNf>SjgZc`?R8o<4W:6\a`8>^[
lf?i_naJDjJbQg@VbK5VQRBiSSkVEE@klYnAKRRh\YjcC7`PO:OeDTP1p@\SbViS
<dkg0`8SVRK:HnC1a7JO319>ICjhR^gI=77C>L1WLoA:LJRO[JIeMCo=pO6?CXSe
jA8dR3SdTA5mc3km3<45=:12m``j>>7]<=mQC7U5fHFNhHe]^UEb1j[a;OkBbj``
3jXmA69n7^<YPOB;LMALCY<XacPi\0o4<DJ@1]E^c@`\G5h;f:S2]_i]\4I5PnlB
TlU2`eJelNG9jQab[pf<hPh^>3emQ<I6jGjYSQDJi=LY1XFF[ec`0c@<loSEWHQ]
Ub3HkRi;542[]=?0F[i6VgnXQE>5Ij=1gG:D9A7U`A[h2kQVAcW\5ATdXRAeVnOF
En[EfgcK3I0TCTHbG8SFXd:\mIVaXf9eX1>?]LRF1^A@0LqdR\L4MqX?H`YSd4fO
k4HliZa>]e\3J_Hl`chO=^?O3f<5RN]Xq=Pn0ZI^KnSnfc]^09e^36I1kn@Cb`GM
fR6KHjONSA?pWTf]93goa1d]1=WBgXW9ZEKM?MMfCb\1KQNYG9Q?`;SJ>;^ZqSUL
EHfKGLi]KmMTm2lNXbZQZXW^n=jMeF4[14^daD:4LDnZYh7HJR>0L0T\gdJ]:ge;
D_?>G^_OEd\aaUB:egSe2<\kO8C8I0nO@<AJOL:?IcDQ`P68G:3LQVCRjA=@IS\A
<i2QnpYjhf><q[6mFT6j^TQ6f9lfB@Y4S@1WejaY=?6lSd`VFqVD87YJP1:UCHQZ
Ki8o_fIeNh`87e?TDej67FUPp[km7E\[fIng_4?DH07e`lVTXbKIfEeF9AEo5G9q
YnhAkJ]eGZ^c5i_oCQj<ThYiY6?a35^G5l1mFoMPhk7^bnCdfCULo6iB`>;Uea@`
R9RN@m?OLEpVVhHln?Ik6hLc0m>\DCJJS7=EA?6MFEDCWI0A9eZ6_AC?jA\YEqiO
n]I4XSA_nV0iYmZV=NZ?3jTSDjFM3iTkHZhUN5`Q:MinbJ0U5]2hE1FcU::>=[D[
ebVHJJg<pZiGGdIabkP?<07A=`ATPf`95[chHaj8g0P_HYY;SElWUn_Il[PmdW?g
hb:I6Mn]0g3M>\=pT^oT1m]$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZRBT(Q, QB, D, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, TD, RB, SEL;
   supply1 vcc;
   reg D_flag;
   wire D_flag1;
   wire d_CK, d_D, d_SEL, d_TD;
   wire d_RB;

//Function Block
`protected
f>OY5SQH5DT^<dKYSKZn5Xb7_XI5W@5L:GBNWJj459e3`1miR<EoKLnoRbMB75W[
pIcC4R=MH8aQ7PkKgkB016^JI=d\qdiU7ck>hM886;k[<:cCqTB`R7?p9VXTJ;IS
M6;NI3D8GnWmnJQ[a;Emj[0gAB45phI<lSLd?560k4`]H;AFhQLV_AOp>j]Ld;Ec
Gc=dQod_a[hHGn81W_apPB6T[bPQ3RC728ELn4H\44\[D]BGQi?Eo1hXEWN2X[9R
=hGn7E4fMT[eMJnQ?d[;GAJjJVebP[Z0ClqE\EbZ:;gFVDSfO4Ng3SF_@oVa7Y\[
KEI5Ah^^Yf7:e??jcAKCo^J?28DaQapJchHJ`P7A83XHBQ]lBZ0FI>k>=J[TWN8q
D5lCG6TfD@_mk9;^MkE^Di=_A;`UO`hQk0LB=Tpjf[F9F7qmFQ\;hB@BC1hh@7S]
cibB9<Wa>3]cHc@n<dJ^_XZ;^4`TC:ZeO4hpmZgP=XTD<4`2C4:jJ]XoX;egI9nA
\oapCZ`Xf2I;Rh^j3e\5DHLZ^9RRQPp6`0iWN]q\bKBW1H\?aVB@HbGWgd:31g[]
DJpW81JVgmAG8B1HTE6ZM<E@2dXVVH6;]0bJlXO74poVM6^G6q;YAXE:Ep>]4]^n
qK6;fO:GRF8;6I[3<f>N7VLmAY@P2QoTZ?DL6mD1ZTdn=<M0c\BI\Nh`C<nZ8:SG
7Q7SIGXEQc:8N48nKhjbZZ2:IXjeLPMf>hP;DG5WRU]Z@p=KFSHYRE:j_C5FbPG0
?n[2hPR9ekHaC0Z?\_==82`]ljLT@VmaHf=:o>=6kj4_?hod8K?`SXg>^bBo2iVX
l1j8El@=R9USHB?^Ane<jRkced;=p`d^O8]K4TLlQ3ODl@iW?0@;fT_8]F?DE2Cg
TKF1MgiG?1g=][cd4?oEDHf?Q>f=>`A^O8c<BNo<=b\6iCg`W6Zi5XOHQL7_[O<J
Hq;RgJ2m\elmR7_LnGKc676C=MBGG:JoC;:Z2008RPQXcUE8BNCdE:[426CfX0XG
h<6PJ6EiSaPe<DUL`fkEb>0on2B:^CdI=l[lI9@naUQmp3nb7`lpK0XA1nj_;F?@
T;ScFe3c_WM8F0OM_i]H=XmMP_bRScNT2Dq@<`5^KkW2F>HVlaZb\;XF?n\B89=0
?hci^TKqD]N5[89MV9meDQLKY0>g8lTCUQYMT=ZTkh1qEH4bZ>f:D0C7=F94^Ib?
;;fINT@<iR]<BjEWdHWq^L01FC8<8U4YJ4CSUJD=O9M;BjOF=\F\2>j2=Cpmb>a3
9MlXTL]@0H6VkiWb8<_cB1L\R;NmNA139q<>L9I\]o:=>6g1Cdl:dnUOCQ4_J`gG
:nCR]:p9bMe8PPm3bXJWI08L_V;e3N_LG@4`87jV:<>\dQV0mCkO:2N;FfhJ7UYl
j<A8[Tc7[QQ?o]74cH<kRl9i@9SQ7>EVNg>^_jU\jVXlOBW_l?a^I8LBa5T@gLe6
=E=_Y?>bgj_2RoP>kWddXemniMq0QUYng]iodKj_2Umh2^a3b[`33HMGY01RhjTP
51YfHZoVZ8VRWLUpFhB9JA5O6QkHRVSnF1Vh``EfBAPMl9fkTI@G4jmR58<S0o3C
JZ_R;h_G3hDi60QG6_X^=@D[lE\=kWmJ49NVDb[?ThNLNO`Y<E:RUJVR=?m@4\TA
cRGjdOAAn=L>NgA>b=WGi7R99`Hjmaa17YDpY`2_jO3N4MZcg0laS[ma<OY2:>_g
VRJBOQ3>1cX0LZK@m=FQ;g@A[3cg>;6m?94F3UMlB5I>CB_OZ0DM?RgZ@>7fAGS@
5PRGn?JMg;=6R7SWTl=_`]MW>57Z<6_PK_0bV4Rg6I1[jHL>JG]THXqijmIdEQNa
bEa^FiP]5FKWAo1JRbc01X5<FDFe:D7LKnbU7__[mjg[KUWg0^:`9>F8^j5;n:?\
k5=5Lac7kf\EPX=h1DM@\CBCn4j:8jF>JM3a@84Un\RGX]92\R;iJmooEF\A;Emk
?]Qk0_bkPq^dO=MaOGlP@d@c[E=_DCk5cAQ72T]2_LPY<mYYW3Q[2ank6]MmhfRQ
Lf4a`NQdHC^H\H>e<13dSKdILEW@bbH?SVXa=jKE`TNhldfCKQ8aRPlIR2WXfYab
eCT;DXo[=66:dP8J7W\JN@BoF?RH3KamHdplb6BB^CHgiH?BJo^N\BfmnO=N1A[j
fgM6hhkcT8@l4=3@^0?bVfgi`?OP\e=b7E0BH[A5X>iK<EcgS4N2e]9]9hZSZMol
`XV3X][m1;ka@Gfc3ji`IXdS[:?`kC`_:4@FdNkkdkIVc;^bC46=g>Qh[bZEVaUq
46o^FYpPKY[OEe;`Rd?3KZ3FW\LUD:U^nWGlHT0P1TjVJEZ;2p>a_78`0FKoGb4G
aD<BbH\Z6VG2M8flXoOX0[]aI2kbpAAQ:3BF]kg^@oXL>]oKhB5iMW:;kY^D1@Oc
Y>YgA?NSbGa6a\?qSH;7mPF3AJ_`NY20no]2TI^0a@JMm7L5dE8`IGb61<EmfM[:
7aWSNOgP6I03LPE;a=m=<1=d\oeaJ<eM3P3Jm8Mnd5R4;od8anLHn5oO14>K81[b
=_Zl0BGT@3HPT^mPe?QZDIgVp]`X_KYqRfe_8IFIOVoRS5cL=RHc`Ua:nK`keVKk
N]BnpAg9<c4Wnea]`OQE=KYQ5<5772Yn:b^4j80=0jWqGKm>`mme9EJ>>cMV=EX7
W@fn=eo<Le<;Y][<\[q:f4NIeW7ZHhbI2_LDBo6d:?1mLSVNjdLK]81o7[Ec_W@U
cKEc3PD]d;SjJVYKBC=<O[Y:^j^okqRRGaC:EHg2;E@0C9]Y\i]b3GK_RIG`ol?P
ZeH^bRNR;I1^NIc0Yf?O6D;l<a9aj4Z7h^kFS\:jqIRAEZmW48E9_4Ao:;bTRo1J
`U93WOf6Q2HTT>j3RBBma]kMC>HXXkM6:=@dOQ5`Pa;YH[J\4Ygp\B_=T<_e8lf\
h;GlKS\S=OI7l_\SN4GkD5HCT@Ih@fL2jT6gq[IeQX\1$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZRSBN(Q, QB, D, TD, CK, SEL, RB, SB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, TD, SB, SEL, RB;
   reg D_flag;
   wire D_flag1;
   wire d_CK, d_D, d_SEL, d_TD;
   wire d_RB, d_SB;

//Function Block
`protected
1>8T7SQV5DT^<;2K`R[4\9_\CZDjY66;i]oQEYF0=I9eT8[MYJWH2^6a6OAGj`63
Y[`Z]eFJB;\k@Z8pFZ=`OBA==K<UM7ZhOoF9PmGiAePBIMbSMhX[n5c5BE2V[dcN
:bdhI:?`Mfb1]f7U?WpmdDOb=]Rc\l^S7M@Hk9c3LI\lR]]b]AWU2Am6dboH7JqQ
;Oi9mp@DYbJ[M`Yl2`:@9]DTa>90:R`FYZPdBRDT[HpmKiD4ioPNKgHM0GSlcjI2
3:2NZq8@d\<]VHo3;c5;?O>KfZ]RPX4hB:q4M4kOoa80lj54O?6=H0:]CjH6CKVE
b<4\3Tg_8aLg_8AIjL3nDOo^2GQQg3h``om9VnRUdY`Y<f^DDQpZf@QhZc4]V6\F
ZaX=nm_NM_6bX[Z8do;lThA5Pan1jH7C8QlqjCo[5EfHILRMbGMo?A0AW1F51GC:
eoNEe61kh4[pm]n6A_C0B`^Sel0jHLAPM_KR1JLFS9mMO3M1H_gLMlTK>fmKcE^a
I2?g]6AnN>7>LKpVDFRS<7>PMjP]Zla[oFFDli^?k<GUGf=b6WqPSHTI7JRE==S`
Ymg_g=CBgc6?giTcBe=KGmWY<1dO5R21gU7Ec1fjH`l^Bq1nQM\IbOC`4Jb`c^8a
=ATY6R<<VOZnVSE<B7`FBIR1aFaaqX[lQ2>HX4jB5SOOT3o_b6A:GY0<VNh3^mOj
R2C]NK=6Yqm9PJ1I1Sef5Pf1Q_5WeSCfKHgY;`aPSnpX_SA=NSU]fD_GlKBR>C]L
IlH6jPmLh^TW\VZNMqCGK10aD7R0@S5MMmhUdHnW27CGUTG>Id\2h0D36moF3@B9
AqQc2e_FDqDe@`Q_S^G[jYYSGoMfLAIi919ABMgMnpNI3SOm6LR0CSSGbAj2I]g7
Q<YGqLidXlh<qVQomndib?aAmPJn;HT@ZDmO42ebpOU[0fTHB@R4Pk1qZ;H[Maip
UjWUdcS>7DGDbFYL6BH1?6C?aYJDS1RaNbf`lP0DkX;XETmC]=<HhYEQpAWbHfM6
Nc@nEKkF6h11F5>aS24[A\Ggj:oaXX;=bBT1CVg7b4R4Ym[]>GO<1E`T<mn_<gO`
G\E\E=H79lHGK3IQ85S@6o`a2j87flN=j4iHq][7DO]Cq?jl\I_pa3V=_3eY6Tnk
fnXbYXW`J5N2N[9PUfQlE6nG]M`@8C4nB>oj7FR1HYiDiG8JYKnA7AD1@[]]fNM_
;@DOBogNoCSDXeZVeeWWC20_58lki5J6q1B2T;PLWke_nU6X9b7ETOkMH_6bC?`V
6ZD`Jj[X`PFYJ;<bkEYAb3>GQ^GH4Ok6IG]2A]=kENl<mfa2;M_g@AhKUmh4W\3e
iCSi8XP?S`NN5l>qfYEK6Kk8ORgH\GhID_4W[DVL13Qgic7p8QlVg[5EPEA26_2c
cAan]mSFiLT6hf8Xcck2@fA@KCZ=1`CXj7X9J6I@]BGhHI\n=50X\YH>gdGN;_M:
jMJe93?KB3N8SbTF\ggoXHE2q`O[L\AbcYCf;TY?gnNQ_3jLH<VGR2T69mD=ST;2
enb6f;j3f[Ih1^0O^nH`R\B6U`L[l\RXNWB0A5lIG`7=4Fk@[?HXGQ;Im9@`_FLq
Gf5HAk25Z\P5BJFjfKQSY5RaPVbbkB6WDNeBa=nAI:Ue;ej2V6hRES7Lm`3f7oJ?
GI5IA>Rf>;?XUbcTKU@I9cKIjYl1;nL\HmQOp1a9eG0CL5KggKM?F8>d]NHQm\5S
2^Nhm\ZQ?ba8mG[=QU91O3aJ20>1TUF6G@HeTHZHZX?J>0k=5jMca2KY=3:JHihD
;9LHIjDkW4USnAaqehPONDqDLR1_:ZO[aN=kD72IU_Xj9I05_c`X2W@9<5UZ8pf6
4M6T\`HI3:PjKgFNOC4J22Z0I;bB\lMXdlpVYL7H\7RU>ieUY_E3\PoCHTQ5U09k
VgU]6JqkYE5J=LeBfKE99En^e;1l_SgCEDn_^gDKoFgbj6qNc@12BZ?e;Y6PCg0]
_Mm@A=jadgMaUP81k5;emqmDLgVYFBKeWdiEVB^c0MYOn[oZf?_1W`Ula1JIpj4;
ZNVcicoRRM<_h=PMRAhK37Ok7ldXh^PMTEY0HVZHW;41FW\WeC;k1k?[2n5[?OGg
`:4p5kbUbSIdiPOR@MKCWZAibAogM5XF\Q8SdI_Aqa_cfK4l1?[Vj>6?55RJ2]j\
V_nLWcAjMQ[MET^ERPSXLa[o7Qa\9cdPTjmmCW81ePnb5\SRe@4d:\ho^1O^l9TH
F:P<B]VQ]8^?I7B2m;::B>BY51IAeN3KPkjYV=G@YJoZmPQ[N?[6=YHEJ@_lD;lD
=?Om]@MTp5E^nPWLM]DcVN\Ic?FJFZ`_C?GffXBQ8aFg=^L`Hl7<TG\a?0D:o994
QFUN^8da;C1KjA:aE4dKSQn8CGh88c?POdbBM<K^EF98KPKL6IA\B6@5hQOEHbfT
3Z0eDk`KjoL45d6iea4>hgA3HL2\o4]PLLA`TBkX?o;Uql_[F4=?1HbJ_M];Ae;T
kdUg?=]V8WJEgXQ7ZBAmC`J9pA^^c_oRKQ_153LU@b5j96?kmfdL9kBko^F:[5<>
GFi1dAY]>nhd^JY6UdgjK@JYT:o2]aL>9;ZK>MVc?ZeSe0UW5=61j2LVfG2bgER[
Fa^;>ScfdEY5bmM\eZBA^D1f5A5iEeg?PS67\JnF4KX7;E=Gg]LgOGhpF^7m8XYd
13Pal=[68BW=YOecLFABgUKQKm0K\PKcj2L5gWB6JH1aCF3VH:k43<2<eQo1=5jm
I<:YU_M^e3jPdYbT<kZVOLZAi<V>>6@<<HKNJjELhF;DjFgL?D1gGc1oFdWXESR^
il19^?FlhTXfLBFhb0U\geqIORoHFL2M`VgRDN:b_f6C?FJ_k_kge82LiUPC=4hC
2NDnUCE`N\lCM>``Kg5m5M`I?LeIlbo?T_CEg<LGNejB9K]KojGA2T0Mh?E?_8k2
^>CZ]`SO7h2PS4One\m8O4>ID2`So_gLb;d`7S^ST;a=6A5SSGIfl:lJEhjqND7n
CJDQ6j3SQH41Bj5ZkmFT<;<^oJ?WaAD^6bh]dmK=SQ@QFhSX[mj\[Zh\E4eSah:j
]DRiFWAX=kR=@AX`4bL4XXc9Ab2IZV2LNonT`IMA:e8H`cnRmR_aTW0B3PYE4n^H
mLBDFj3ShRV^Lm@T4F`d7NXohL]c_gR1kQLmp^AALLPqg7\7Igh@c:RBCHl0:EKn
R?oL`b[02Y^Q_d_iZhihQTqGUO:5abNU:Gm1=XY:PHUBQ39V[T^8H5HH?=I9[mGJ
EbpV^17UJC0X[9<QcU2AhP8lQ<H8<MmFDPiB7eW=a9P=;G98=JqVR:JbMheH0C\o
klGbCZ@aomB^eQPeI=RhILOZH[]g`pWW_jgJ7_^T4?XDOa61JGP<FJMP?cd<EPdU
1@BZT8laq=Bm1h37I6@i@>FUQ;RF4I[acD<1i32>;<ho2mKN]9ZSCDnSbha8Blm2
Z4C>AS`S:JcF;0DTf]:B]AJmhEB\i?Vj5HU?f[jj\IVn_BFXYWJ_cnH_i6fm_Gjd
]_FXXTMcS<T0K4^nZq3cF40]moF:30e8A:kPl>kh[2HgBSO;:IoBXbHTVe9<K3CA
Z9PUdMnl:TI\_\XK:E]Q2ED1Ui2X9JBDL^<WicbCRM;19g@C@<YIgQLQRH]KdmG9
WL\@LdFB6Dh]<ke8j@fOO9OTPT3Yqe`OLmJp=g4l;i=P8:4GT4K=AI5C<NYXJX82
=CE?^kNJpSEAH[QVI_K2C<aMLPB2NbU7^DEl:?jY9ain0E?p0cRYa^GHSdf77Qa5
k:HlmoX;dWWLDo><LN\kOWp4cIfAEbNJ_A0eke96\7SNdaMFdCmHZCF]MDgG7p33
M=N`1Oi[01j;YUhKHZ>EMC_MBm\Z79HM^JBZ[G<>gOh73O=Y<f1J9kK1pjk6@6Y[
\o`_8Qd=BgV6TXcKZAcLdbRjac5f]Z_ZDYY@QHJaYK>o\GD8\dBM2ga8fLOeJHb0
dl8qbkH;]lZFe7[RRVULDH_eV94::89j?ULY]`4X6<PiDjMh>i=c3Qf0aVR^b3Q\
`@L?WaX1ZJn]>Jpdaa9?DBH\X;IYmd_0Od0^4KmHBPf3ec2@?Ojd<]7GlX6D1DX]
C4ZcXYce^Ilm`m0@h;=ImoG]Eqag?6<GTC:=OSNBGgE[q>T]M89Pbid2AYCfYLDe
L218MGm]UPXS67i]PS@Mi]XCM44S@ZCeP7k0B?EXZSOo7<2ccQ]qT>HUC>C$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZS(Q, QB, D, TD, CK, SEL);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, TD, SEL;
   supply1 vcc;

   wire d_CK, d_D, d_SEL, d_TD;

//Function Block
`protected
<lGSmSQH5DT^<4FbDh8=ECMX>UlQRXV0qb_;\i:VCcK9OMK=mSb8d?foUUC3GqD:
nNJ28ekP3=3ICR?[<M0Daa7Ab:`4__o_RB?0qnM``KQqX4PG_\jk`LJ;4nmfa>PE
2e:^bKpPFC=S640T>W:lh:4;PP;ON0OkZ<pSkI]C3aeG2hh^3;DO8KFg6[aCSogC
97M8dA]OZ1Fe=EM=e;lFAk^70C6di4jVIG`A1HhmeEWaSJ_qgMeXhMjY@7DP@?@_
f8nFC[J@Y@OPZQefm2W?@]TRggKQCAgfFnSO\<]i05<Tq1Aa>VOnpCl_5S8\RoPP
@=d<h7W4pX`\\F<q077\Q?<kd=eKQ[@OUPDA1iETgmXD@^YSf;kJ^a6gnL5UWN<X
6@:LI`VDUQ`XFmDPTET^SPi4[J2\W`ZDiHZ<NJn5G<oEK520\hbbJ:V4G]Gep;[^
j4gA;9ZEfNK5oH3Qom`E8f:@3h[c5Xa32B]L_VVlT?cTcEa8FKd\l>Z\[H_gaMcc
ZCb]2bK\ZSG86RIl?8`hW6ZF4UG9n7^D>e5<<KZ8eQ`pCO_nn=qMFU>JHLDQW1WC
2TKGPRL46DficO8KF`I1Igl\Eq_O>jh?mjbWTk1=I5k]oBP3=4UfS`=cK@0:XpjR
jjTckdf?jVl[oYdjjJ1QL[d[n5TD3KOjMITD4Nqal1P5gJ>ci1<8kUUK[4=eU8gL
j4I4Y`^`1^[A4q;A?XSon3[:l6im=aL\C50DXYCK_OZo:AeH9XNmDq7?944YoE7T
6C?`j\ZncK[K9W\l3KijR3WICOV9Dk;>JD4[181gI34fGLCAQE=?SpC`XXHY@Ga2
;_@cnFT2UDmfVj^?\i=V]f_?^6qUGPf2d[BQ8EjWVSnNG6Z06k`U=EX959ej`D1:
96L;U@61X7_B^aP08^fA6_MH=V]h<AlB^[RYW0D^BQf4gbhRSml<6TFXg7M8he^?
=\k<ER:cA]?3ZCiOeFJIU^16Gng1D<MHPeT`@0p?4L>JZiXZLkooJIK?FNaB9SlR
[Jk[OL;R3?XVCC\S@[l;Zm91eaJ6OajMTjkRLl;8Pi1^E<bE7MLN_7lY?kng\9[?
D\TP_iOTGH02g_FUN7]73UfCoNDTFTc`DY7a3bgm0DcQZfkYL^q:ZmX2L3KZ0Fd0
AKO9ZJ00YC=8VN_]hQH_i>IM;E]^CYAaOTUlS]IYZGli_6aCF6O83:9nEG2X:^YG
@VRNk5kFc04:RXMP5G[l0OTmN:=<IL>BkXkk36YASjSn8eOLUJ``;S6l93k0mpjf
5PhoSX:fK>_XfXiMPB`g:XQI9YEUh=c50eVc\6E3W29nA^NNSo[H?8Y@iWEe`mkh
G3PmhF]WJCg01L4S9WemZLOD3SD;L@H\gmLLj4Nb@Ua3T@]HRfheLHLPYg;d?VEA
_nV1GoO<p6D=>kV[U:;SlKoNgN=h:]o2`UnVcCN2=VXDdC8>H7:In=M^9^=D5YO=
fnOKViZPb6Ml5Om\7I=E@Amj_B;=S?Lmbm;eBm<Rn::n0DnB=6C;Kn0j1mQ63L<a
?A[1fNg64BaU\a^\SDmD0\k;_pJlPYeEcn^Ykk3V5?0mENWjgA]k347JVgJB9HRG
W9HBc:PVW388o_L?067?BmRSW_J[RGe5T=i`llo>Ek2NA8WcU;L3;1@XXf:K66]9
jc1RFiUgl:kLBjJ?Oo[A\KGW=SnEE_hMQ`a=9CJKZepPTN7V9g`LMThEcE3gOA@g
J6oZ1l<HPF^IOHqg4JWE1pXF`?]BcL@A\RmTFkk:`ES^g=KUml@mR0Fe[JE7pLAE
4e0CX3S=Si]\OhHUfT8VDX1nL`FL<\`V6alqc0`aPflW557NPSY>geQn9IEX_fm>
o<i2?Ij\TC^LNFFbHG>YSe4R\bY<8;3IE<:[0<8ZbM^jb;qI[[D39:WF[QAbo][@
ZZl^>8nfJY7kcn7WVZl63O\20FU@iPI0]Lj0kY[KNqcV?8hn^UNMk49UY?R:K6\^
OeOeRD6LX?oM`P8UT1Fgl`R205RXooRMMEf58hn`eVdbC703EGRlpN>[EG:n$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZSBN(Q, QB, D, TD, CK, SEL, SB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, TD, SB, SEL;
   supply1 vcc;
   reg D_flag;
   wire d_CK, d_D, d_SEL, d_TD, D_flag1;
   wire d_SB;

//Function Block
`protected
TJJ0ESQd5DT^<Z8`OLVV4>b`5:117o^;\;HT\C\FTS9T;Iq[QVJ<d_le8dP<Ef2o
a_=T9WjfC_^C9=WRW?fH2ZUF8_]_WQTif7h`=0@U1[^d>]Rn4^EpnhdhUkB5B@c9
\OIS6DWZlLKp=>mHXjpdKEIPZl4Pame[l^6=?99[;2F?W5n5l9=K^1Tpe_6C4L\o
SnV2PBIoV>Vi0gR_ESpF3UU4hRO=T`VXn9a[2LOQC:aVPfqOPLK1EZ@Q3_mchK?\
[`@3KlU6@_XAUKFaJN;UcBo]Qf>nRPmCc09iO=P2@T]4UmQQ324j]=g4W:PNCpHb
SD8g6efcF;lLM9l6fjlg0=jKk03TA?7f6nCjT?JUQf5He?hY^:][OEEgLp`8AP<P
KgVP]2k3n@nGL[@eieT0RR@hA9;EOe>A1PZ_YKEOlNb`kC1P7M<Xiq9\Ho9T1?ZC
j[Y[Dd_K9[VQ6eUeLIB\c1\`q12<Z5<i<lJCm^]R?^R7U;\cii<Q0I4meEOW>4:O
pKom>IF<p0ZYCB5;B^AUkFI`jkVWHGc0blS8RY_9pY6m;GI[Rl1KIoBAX2ZYJ6TV
_Dhp<UlA`H>qeeZmCS2[j`=F;GT@d5Z;\G3m=L1pHWa_B`dqXO5[eAilZh[3OU>Y
G\[aL5]Zoo7Q0Tcn0a3K[]o_]K_l1CWNT[pT4hW^inpGhk[ESq;a=g]14?Pd\DRJ
@UMM>4>UJ6SANj@kd7jX8n]P;G6bP74UhTi6Jd3Lb\dbA]Q7`[Q1Ph:Ae9bK7aBA
EnY2Q:i7>KJG=l]`?kN0gXYkWdLaH=pk:Kb9^[Y>OcZ8<C_mLi>MfZ^?alf_LZcQ
0]iPdBCFI]MeU99\Pf1N5Sa8jcdc[Y`f;L5hGC92[HbY\8Lb_e:6jP15;_N@^@Zm
<QiATEdXOI7I^pXJbfZHFK8E^ZE0EYobQ0aCN7WN=ASI_:WEeR6hJWggWH=1F`Di
Mi<6Dc:lYji;[ZXNbiZ35KRm7B24_82[KEmH_35T]CkJ[Wk]HgBYqc>U738WMO`;
^j<5KMe79aV3ZdM0dq88P2_]1Eo`?:Oi>6Cl]HAnJNd@E6ijBBO?Ra<AlNn9`U_G
^H1`m2Hj?=5Baj0VRC_Bg\K2@81VDMhi@`HYdSUSCBfT[n1RS\jHa6l7LSqGJ7i6
4qbhiXR9UhJ[LE>5I32D>G=Y<YK4_Gk1H0ie=LpcV`UWK;^D72O_?g@5k5o6j0E`
PD^ofKicakq2]5QM;RZkn`ekIX5:Doco2bWmNIldA^JZk7hm_Ipa?IFUm:h:6^?O
oQgIJ@FgPZ<CI?aZkMkOh:M3jp0OB@XBI<`R_=MNIoW00nNdD8AYA2QF]4DlJFe<
qcVeFGl2nMLmZTKYg7LKTHmYS8IRjH5M<Q[SEEYef4aN]aPW7kCRn6?4pbU:Vk;K
I1PU5P^Dk1hHonI^aYcZMeL9hJn:LqD=UYPXf`8F3FE5@@6flXYo:5l90IQ084]@
7G=;=N4j4636?2R4EAZlPa9o>J]H\_FaQH2[11_WSQ_3l[0C?T?>ZOo418TECDN0
a=gT7Nm>5<I>BPU2IOW;7h;VYCZmSWmo@0J4`9UhOEe>WF6XTq1He<V;Q>BmHUJ;
8CiNU=XTWolRmBV9ch=\^YDV9RaG5nZK8LFWFXK6:Y`T75ZYifaOm@X^IGJAhjW2
3HReViEUAXB;lW_iG9kHJ><L2UCnD7mI@So0dceMQ?E]:8m5VoBPd=JEmJhoL60^
Q;Zh@FTW2p[Ik<io93``:mg_cFB36[0MnWaAX94HI:k1<X1]:LP62gM^BaVlBNMi
YSPo99aME5Wb[[@Q4ETRMcSgieXVXH3S3HRUf[n`;L\5lHUL>3f79D1SWJ6X6iIg
7UJ\SXBVd@gZC^o_IOoBE^;6;h]2q2?gc?L[fJ[WEP`^\YE0U;_Y`TCe\XLFgP6k
d0?9P_?HEi>HmeoE`SD>1h6CgSgk];9ofB=Df930Mi5CmIgcSKn>X^Fl7Kh:bh>6
f9`_:cW0?eW\n?@H7QIHDc:;K9n50\SakESQVE70G<[7^GKqBN`MHbRk37oDk>H2
Z6]1eJoD]jIT;^YHRRNbC[R@1konXM8P;JNSQ2C<h8ijXVJSBF^cnRF]miYC5lII
nGbDGN5_3@hC3ZPl=30K[>gd=T<GL=eb:<2_ON=dB09OM\iTGjZ62af\d0UMPnUb
=::RS3gnp9dYn`o`[GIgH@:7@mD8iGQKJ`\hD1P^KjF^Q_@eIaThK:HECcCdCDj@
M6<Z;cWh>gVn4kfPJP1M0T]TifbFjM7Jk\6UiWWPe:On_UQbHl[?NNGXPOkZc5ic
@ATNO=i7EZjNmY=0iI3NBnkGg^ja^Geke8XYFqAB5DX\X`?N<SRYCn\B18]Z=ibJ
_kR0IjObepXhIULmp>?I;4jODbMXjdcEMb6DTPNbb\NZGXDB@d?afLbX^=Xqe;fN
ZDihn;Y4iX5L:achH[SMmKXHMZb6n<X?iBSM97qJ88`QEWjgVO9H`N:UdMIJ@gHe
QKgK6B]59\I:RDRP\MGG29>:KUVgXk_iCm<00:ZZ8IBa`Om0R_kORk;F[_?S[?QJ
3WkCFdCa=8FTI`56Zl^SYGUVA3@8RHAk9E^5fH_Xk8I_[_bICql`;I6kp7@CE0cG
5Bh;I;mZ>CMG2W>P?24qSUT@amj<155\`kgYU9:gfgfP4OjgaGdQoMRgd7qf\T]D
X4Ih:LL3ZX^g@K]Q_gL_:jR`UoZ3AdZ6`p_GD6321jGW5F6>IiNLFRF1giD<DJ??
oFE<]@[_qFFW>VhFA@^i[\TcQ12nDUF2<kFD0WRTnXWacG4Z`7hce1FQeA[MEcmM
IPITleeXP3K`\oY4M?eq4a^lB4L7BELU`7VUH?DbOmKPM_1cZHB\n4ePoH<OREEL
M8WgGh80?VHL7`dbC<UiOk8b_30id6qXcJiN=0@b_TaD`WXcamOf?m1VIKeAD;m@
0==E31SiUgP_g^>:`MG1E7d@E6nalL2V]4Z_7qTS8;H0]iQ[;XIdL7<n2LdCXPC:
n_aMl691OQ=M^LR29fFL@hB?6n99<PJIk06I[O7ZG<7^pTWcNS;h$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZTRBN(Q, QZ, D, TD, CK, SEL, RB, E);
   reg flag; // Notifier flag
   output QZ;
   output Q;
   input D, TD, CK, E, SEL, RB;
   supply1 vcc;
   reg D_flag;
   wire d_CK, d_D, d_SEL, d_TD, D_flag1;
   wire d_RB;

//Function Block
`protected
Q[5DFSQH5DT^<:<D0DC_\H9kYA5RA\Jf^6InnnQ4H5[L?_BZ:of5CZJ9`a\pZH2k
_O@KJBQ3X_Lea57XJJl>;LHB3l]<iJ3PXlnq]iX@]5\P=WiL4U`9AS5W9FYI:;@9
q>?_4ngpVGPbT>f:dbcC0SUhM3DQ\RS8Nf@dR2YeBiVZqbGSCfXEPa;8]>XGhh23
9W:VRfQY>b6NALC<eADSXB@6\:IUn>[OACefj?J;L@Nj;7NogV<97BZIe]HqbDPG
nUdFn<2QPa`[`hG6G4>lbCqHd`[XTX?W:^AkWGL__FGF2R1BfelBi?HpLkJgke\B
=Z]=4aX;C\C[Jd=cj?6DUUIbFSmKZXngh]VEhhXBgUhZGJ<JhoGqSIoenhk9^c:Z
dJ5I=b6o]5dD_X6EL6[epB>i`h:^6mb[E6=Y77RL4Wo66IoS6f2L^i1L`o4qMReF
RY:c<]M1<OF[Ydd@TY6>;22?c[[43l^mf=9lWC[hXUJZXCXVFlkNpW2K996>qTdY
A[l`?j=i[^ke<V7kKJagD^`e>VT:q3EAnJKfVS`1?NMLTg2JZDAPVK`qL=eJ7JIq
@4>6CLO>035YF?6Hba\Xcd:CcSAqS:h5hB9pG;T5fA]EWc9>43@HZUTX3@;UbaGL
7OR?>39m69[Z=:gph4Kd0>Dq\5M<YSqeJ9j\ZTieRhVLPBY^MhNKPL9cJA?dgAKA
72O`RUTB7g2==KgLUff]TYYfO42C<ilo:FDbS8m3lU?kHY6fF_0bVFYRAU4mH5ag
>QEkC?HOT\Eq=HUDSE52^;jbcGPPEL>\Qo\PYi>kC=[IUii<g>b7<=]@E_\LH^>E
l8dFcYLMPbbUh;_GN;MS:?N`i\U7M@MZ]R8Z3Q52InR:>PUo^]1Z`7G9c?qZIoWN
\<C?8VEQGEDJc_lOdKT9V8PqK5eU@528:NZ^KJ<MI`o6clRF:jCD8CMm\eEn28;=
LaBd6`E0jRH4b]Q^4^nC>i7jKFe@@N?ZS0NPlngoKIc\g35QJEcGfbSNZdY\qZl4
Q:_Mi:n5Eeh19@2Rke3NDb=1UEGZWjn@YFPKke5C0mkkC;bbR[NT1\W5W@@lO6_M
F@QC0:4gP[e^FPa?mOUDmN?Y:mTXo;JjDC29?0mpkd;SJ]em?T:\I_Hn>TZfk:bT
gUWlRPc;d`@E>`WKP[efkBOa:NQDAhWLJNlIfc9MHCPS^fgCH9hnl:NTT7UjjUnk
OLC8;leT`8MSW^HIdOdYe@TJTgYb69j:ZF<c4;PD6L:>4>XJNf4284VKE>R^BFb<
5PWUVPIUT<@BSCe@kC3@k7@JfNnh93eD94\CfA1<W>l0hKfgqjD13;dqgh[RYD05
DHFCenmGfNW6c@G[ogLKe@Sh4MXEqYT_:X698O0a;DRY]gJ^JBfEA\HXJGW\4E0<
qcMTfaRHLCABYBgmM12d?<_D9VGSibM15GNPj<3Y:InV70\T>AB\6[^`[Z6p;QcN
dLgR;fHCW49?g;M@>Nf7>`2Wh2ZBOL1ih9iq>9^\W:5h8l7JScGUKAgRH[L:9>UK
k^m6`0gVfaqQ;kGGV6a7WZRR35Z7ZJjO3ROUOYdJf:nb_3W75pYT?Mnbl;4n=\f7
blCAjROPoWK_?Ug;A86i:>qAL61\<dK`X[U<a4DN=5QSk=G1Si5Bc?_L4<lb;H?P
P^AoJ]M6l2@SNC<Yn>Yk=@:OHgT\YRJbenV`>KR83hk\[=3EM3;\ZP7mY5Y=]N4I
Y<2Z?LLLH\Ueelnd0HeaFoY0bY;<K5LJXen?\cgVX8q[`aHg5RHR^Wf>JeJB:SR8
fk^\Ce96@bUeL_LCPP^2dX?<mhg6^OoTMQJRRl@cD1O:5NcPnGeCSODbATiX_GQF
Aj8U[^e`gQbD6eT4O`AgohYC4_G\RG;L5HI2k:9=\Di3M1:imBDQ=YLd891_L2pG
1E7B3d`J?<?cUDA4_6oA6?e^[IfaNl4PIdIV6VJi1_:UP3WP>goUhEIqnk5ITiiW
j;Z<7`;g@^nO[<dRnVbjJmj3@AdX52aOZIFB8j5]TIWUd0NmgDdnJ?^h[VBGYjN\
@a]aVJ^VPbZEcg2bODZl_11Ijj_4h[fFRFd`@if]WOEiQ1ZfjSJEe@`9idK2@[8=
aOH7N_n?j_pXS7n2@4ULUHea^iRmVWJg>CZTm2>SVIA@KJRSYS``@=4]292V8I\O
2jfd?S9iOEEDFTDPFYUOY2H9ElAiP1jKR[<gPoe>hjGl;Lmj@h_6ARlZUdi0QY9f
Ih0CJA55F<Q_HNmI0e?JmM14Wfj7gq26?Hj@N?YB63?nOO:1\E[n<]<1VJlXG@Dj
iKT`FW9jlFB\giX8gC=3ZinPUIXdZ?2OaiUda5^fSM^DBn0UQ;<?8@^;`B^f=lf^
iOoP@Sb[_e3olO[G1A5dAb=a8haGbDl?^5dd3UIOP`R83n6WZ>LQ9Vp<1U7Zfm9A
D7<R3KGj>A0cFfjI6N9P6ZB>nk1SAb\OEAWIS3c\>^GENAVlV:E7VY6Ob_ad6TX<
fn;kn`;Z:9Ci`^9X>V[h36Wb@`c[CDe@An7DKB;ADlAN1S6UVTObkSW;^6XVZQ]J
f>I9?X?eU4ZY4NOa;4:qiKe`Z[QQUgAo]c8K[UKbSM?iB@SF]bT3M_0KNTnq=0VH
4?pgV:V4:?XAQTa3L^U;2l7c[H1MQj=@;`RLW20;ET_:mqJXfCkZa^jiW?AC`CAP
70FUk`25eP5\c?F3XjYYn]=mqZgRnLSW:e2and\27Ah7m3<W5llV3GiV3QcF8Vg`
2H2mmgJ4>Uh10FG;`eRZdOAlmF`1X\``N^Lk^^FFj6OXDFF^4eOa8KoI>I97J28b
14QcDUk;o[Xb=nH\4H6[?lSaU^DJV@l>2pgUD7:3gheM=<@WUJoI_[bgXddgX=g;
3TD2nqE;ZNH1qdGliVF^O3lAZJaajGXmD=fhVH6DN\40POT@<qZg<=JDP[:SWR3N
Y_BN4j=3mgO@keTLQh9O0MU>q^LXg@MR`e_>Dd?S^9n3HNG7@9bYj@iBCi=G:Shp
W>?NGA6[6;`3A]^PGG@imcI7ic]3FMCJOg7qoaJ[ih798=8\b`Og7jaIg`ck1dD:
3;ajY3L6\ARJL2f885@3lFhJ=8?hj>=gg8@c>S_]ZI;8bPqS`d@]Z]jJmc0U`^ll
>hi_boA65K;7>@8HnS>]8G`kEc7T`0j]55DV?=_I?cd2e?FTWF3P_@O_Rqdln5Aj
`ToRh=86OJ>aQ9Je@J`Ze6DibcNAFH\aGW9dXJW`h6doj_Uo=mhZhQKWLBfI54F?
0bRdpI6C8EL`$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DFZTRBS(Q, QZ, D, TD, CK, SEL, RB, E);
   reg flag; // Notifier flag
   output QZ;
   output Q;
   input D, TD, CK, E, SEL, RB;
   supply1 vcc;
   reg D_flag;
   wire d_CK, d_D, d_SEL, d_TD, D_flag1;
   wire d_RB;

//Function Block
`protected
nN;G9SQd5DT^<]cR^eEoR<6gne>O2\]SVeTCX:6;cmgcXiRV\fSS<jlYBS3\53`2
I9hXmfgHp]S<NG\[UVeN@ke<K1TJi=WoC5fCf?\nqb`R>RbYA2f=@N<cEQo[KSWi
Fd_UTHnn[TWP8ZiC0?og>k]h0A`9C6o@gqO9NQ_Mp9`@PkCL=YZoTER4nNa8VUoZ
NVUE<jC5^4KQ4q?9:<1ERS3V4]c`[e;0of`B;YUCWFUIK@Ufb0GREA4TkS2LYeF]
EUSl2KYTc^OGTXGFD7YXWMC?5a\Sq6Xl4nGedPO<fEnN3k@hblW6:TdqDK]KemD:
;PHY85L6L10D1Tj\b]X\k<AIqh3FN[^nT6nL2jcfR5o`SZgWTmV:LlYNR7bf]PL2
HYXVXNo`:@nTkjb@XFn]pdXB?:FaBkIAY`Z;TmdDB;MQI\Vmfk`hkp`QO2HjnB5=
h[HkXh7QV>R=b2;5MS4G5O83cRq;n[gif`KbHF\6\SR3nbjFehnRSTX]:cM@=6g>
XqQZl97F`qZ]n]?DNA5<026CHU6N<U1\P_dUEIY:8p0S9nOMGlEk9S[n5>[nGW1c
KdgKq2glH346qV5[J7emBm]87NSOV6hQL1I[I8L1q8kn`Q`[q;?ji<?XF3]<H`PI
acaVC9`=ejchRVfY?@B4WTglijGmTa0;ghB3nMcn9iOV<0b]lDAQpfQ1PGF4qd5D
P9KpYKRl7>fcHT:\L3mYP^ICGMRWD>g9Ig\Dib4gSC1K9SP9Q0IP3[0QO;IL@d9F
LFYQP6IUF\`[D7[<aKNR;;Om?048J6h>anl35d]@[L2jKj]7q1TQRPgZ9Ul?ej:n
o0ebhg?Hl[49PX7iLG92PPF^Jgl9P;71qi0;WV@g<bDFR0l:Mf2F<`oCgif[<aZW
RI=HU>;iTNH]k35433ZbO:@:Z4]KWRH[D;4Ih`cobZni`Ge_Ho]]IEo1o_6eHg7o
HTVaE^289R:J[fmpT`C8aMSFf38LcUai;6XREk07WP3@4N]1@V<Z2fBmX?=PFdlH
1MkXbF9>kEQj6K7:TgCVal7FDBH<mKhAJFBMRQBXAgY4b\BM22^npZl4Q:Q@n:KU
OSei092?0Qk\k5BDM[bSP5D=UjOKNU;dJW0fX;RGT:iL0gW0UE2F9Z_4c:SaEd[5
<8h91D5Hg=SH0lRRW7lHABJKa[Vp7>7oMiG:[VUQ[f<28WgA@5@E=G]4hmULZEAd
m\OEWb@@A?MGXBMY6d]LA>ga3e;22M:Lgiha=NO8Nj6Pn1M4HN0\EcfYD17lHG5G
BW1d0>nmV=0gdF3G1KK0D@GhK537O@3I3bX_4YEPlK<BX?`E5c@hVC]MZm_cP7>F
B[?W0RA;maS5d?R?AACU11d=3^52ng\oT5:op7?JPSQqC^iN`aFm;LhOgU>j=EI`
JQM>kGc4Wc`=6m:\qMPJM\<?o`c2@VjHL?4SA9KLDDfJTcn?dWg]q^7R7HmS5j7V
;7WU37nBV<^gbY`A[a:`6kESXV>`p]j<JC6EVCjf\9]\8\iHjH1>>mBdgIkfekM8
23@UBXPPEC7`ZojYU8opLXcZ^dlP3CQKPRU;fA7Q=m3oT=47`b19b@f9OXq`P>]N
deAFSI4RZJ]4PbSfd>K>@cW;d;Nm3GHE?qkZdC8L`g3MJA1?o:DQ[kUoS0=N]AK@
:Y_57ZqfBkanMdFB_klg3UNHX>7SXT_CRV??X4c_G_<RZR4lg0KEKP5XTJiOillE
l:`AjAEDc8niNaU9nANQ5aYG9`K_A1\1YXVQKX];f[_X_W@8j@CK:R72NdaY:cn7
C@0C_R\\0laJ1iAiiok4BX_@0@qSiD;L5>h^7ekMFe[;fD0fk4TnE6e7Mgde?T^>
fP\Qb?kS>7[^kM::XVnRc9lD;64PP;Y26HA<;b:X?:YjCZ?>==VMGSNL]mYi]4kA
?2Z=L`UY250PSX\Jd5\kmc5]0FfNbm5>bhXO2=1aNA@=_mpK7lXaIA<n2o^YOTCY
B4;]OM_TI\:HM6IH39K=MZW474;l_:dUMKmNRhJ7bfg_kc45]6kPZ>=>=V>9NBoj
9PlOZ1DBRR]>g7lIMWSO=k;I29:XHggkId1hdl1BEi:`6d4;nk@K9In\bAT>nG>B
8pV_[:N2EV[0Tk\U8cKB<ZEi4kldECjSjGg6>>B=dFid>2eG=6QcLUj7UR<1USRZ
2Tmjjk;P6e78JP7^aN4U5[GIFV\8>`Wbfbe8H4FmD4S60`g1am`3YQ9oEBTnhfkk
aOeol^_=aWSMOfJcmcB?qdb\FAWFSI2O?h5\9VIHOWlkH[^^dn42;803ecMK3ig9
2DZcd;:U6dlWo0\_b3BXQd5;^T_TS7l[A=@JUn76m`2m6oEA`SHE?A>Roig9\Na[
F6AU\Y6oZ2RLobNm;gM60mNhk42URbMNIc]Ah3m`jHLKbp=N1>Elo9D=Fai15FJ\
UIUGP]o5jaM@0TDTWWnR7QXA;3F^5D@0hMF66lRl004JJMnA:Z?>7KbaMM833\Wc
nHn?NlR[e89Ci9@GIcdL87aMOCdIiQ`^1LDO4B7;OT^`meGDia6U2i]37njS]n<G
ccZE]4i^B6pESK0lJg?Yla8D:FnB1CYd0PK;X9EkGATB6WA94PL=gKn<<ncVHnPj
HIg3B\S9HMXpOh`G2>qnXPVn32GW33kb2WUjXc\XB3G2mDYBDA=cE\iGL]U3jqAc
g]JPYmJ\S^ofFS=na96ZNZHFYU]h2blLdo7@oZT9qmm_FgUhAH9:>CXRP29VfIal
:E8<P8XfRNP9@B750`kc;ghG198fZJQGbRT[3^\?A1Z[2;_8CZgfo787MioL^FeI
3_I=TbOOA:XaL3@=P^g[;4PcV1oYedb]IJX7<]IWECXnc^:\apc1@3H]pO<iSAjA
meKGMc<mQ8F]3C2R\2>L?:ZfifVSXqlZXDQSOd^R=<]e]\]lLd[21`IR_Hln4H`g
1D1jhBXRTGnLNaL7`_MT]4fGR:mXq4ggU>68mZFYZ4@c_FPG=<X>=Z2LAQNXSDK[
PUSpGmRZ0oNH5n_f^kiNJO=^Z;3^N0]`T7SNKdhO1mq>24da;T6QV9ZRN04N0l8j
ET3YK`<\KND2dJ`ilPf]cVDcgQnMkXFoX0hAE1jNeO[?6T@bl@:3?qOC1F3k18JU
6nJ>hjoW4eaDA6fKBBC>=I6X^[I85K@9\n3B1EbYZDNZjSOm9<RPFigW?\<;]^@8
qXVIdRkS2=j^\864PBb6@[hGUNYCfV<j7\BN2@HW`ZIR1m<OI[0?:K`Y[SnicCB?
gkI:=B_pTCNfPej$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DLHN(Q, QB, D, CK);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
BknFLSQd5DT^<^biba3aglT:K4NqVcC=:CVE3Xlnl46BJ>VMPC:1O8[o>WjMFUOj
hGLFJo=^4OWKMG55HPiA4hUMqFcfIK>BHa>XTfm\idCmGHDNU4DbK7bF\3BhOUQ^
Nl6D\\MkK<<e6b3jD[cK3[6;GD6`d^oKpVa\9Hmq\j<fE:]RUkGNWoRFE;iSU[@d
11p5VKEeNAb`3NZ3kg:4ojQHl^gAI3pkCWHmnJl7XXKgHl:V@QO1HD8l6fCn4DOe
=?@QJlHeV@Pi\<4nFebO0A?a6@Y_PJHk9>EqTnY_Ze4p@HU7ZBqcKiZZ1fDQ8l@1
oGm]j>`C=Q57SbReRDGNmi3:bk=YVJBSVI:\^nfkNOIkiXq?]1SFn;Ddgm@Rjm:Q
:5Iih2jkOE=\@?lMeGe9WA^JPdQPldhhOCg[[W6W`Wd@8GCF\e]YKH^lQSkH1CoW
_bd:lHJ_iK^J9aR9CQ7HaajVAOgqg\S>m2F9EZ\8WV9Pc_DBnoG_f^MOF]n[;28U
gCHgg^PS5GT@=<bS8\=;^bRnS2W1ON1;3MVTTNlQI\D2LNMJR9k``2K=F8T<Nl8d
VhFRDc=eKnqYa[H>C;bhSX^[coFTfGQ?b6i9NdXWZ[ZMm=N0G^UQ>NS1@W@@6\^P
3<VKlO5Z5N]YcCg@5DQPeRfmHA10>qUdZYnF5PADfCM>]\ZBK>bQG146fUC\oK?K
;RAI1aknh;NYDkYOIUNW0@G>Do>I0Rm_MTE^`hP7]V4g@;@kYFBVEd>iPpWAdjSg
p>hJ<[CaWXS?ZKMHLca22j5^gj[eo<;6iG`OE\Sqo^<310hMJLbZ[eo2B8=Oc>a5
YQO4Z6K85Qb3QbIDAPjnO^A`kG=]U71QNgq?]]^aYZB\5oC:LWKAeNV0N78bOf1o
>F=2GSp3cF4J^XkMO3lQBAbkPl>kh[2HgBSO;:IoG5cH=V\9<lAJA:`PUdMNY:kG
\_\XKZcoQ19D1Ui\V9GgDL^<0K`bFR_;1f`O;lS4`1;YdR<O6k=k1ZkNHfAD47ih
ne8pn;n@8:\XmWX`Ba43JSGSU\>2F8:;7BJ0mGViC56nVU:n3_TkBM5[3Si4U^Xg
T=JU`fXn^NMA:\i8U6US9nOY2A?HN<?@MPE7DY77A>Dmi4cB^SUha9m]n19d?2f4
d`=Hq;W9MZJpc6BT0mkIX=YTg`jOKUbNc<2WIYAa@bJdM]ZJBJp^DnO>MmG9h^Mi
WT\j=;LQnCf8EH_Ohd7ncE7EL]5Jg@dUL_>P0IgNQ6`nm67P3Hl7KiC3Fb1\iqkj
=Z1dRTYN_B3cc\:<`3e^clQUSgmSpaNaMCa1$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DLHP(Q, QB, D, CK);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
M]@i3SQd5DT^<B\bBgfSTIn`6d]8Tc@WmOHnf=5OpZlV\I6;e:I05iX9d0Q6]o<K
8QPqkcJXDNX>bcLdKkpJGRIe=pG6A[^AD1:Henn5l;QPn5Tm5gY7peJF2XMXf@R2
hd7dVjP;7a9E@AbHqldRWS35l;@_`b=X5X9A_W8Wf<TEc`:Z`A3mekEj78m`jTiP
TeJ?@UGAUdZjN7]2;lVKMqlMYEE\Vq?W03O1pd46^W3eBKmcW<d[T\Bi<=f0_bB\
JnZ?4q8_1^jfWA>BW1NjZFjV?dF73`HeBfoaKP4TZW9a^OX016o1gEjQochK5BdG
XV1I=:1]Rb1m>XG[k<9FihgoF8aBGni7BkXJEM5F:>>3Q0jJ7aqD01l=CDo^DjhQ
O=1A>KT>G<SMO_;O34IOMSVKm[j[;7F;Lm=mYn=mk0n:^P0KD=19ODd118ac_]8e
=\YHSFeQ21A>06ajbld6B_RG7?bC>RAWIp?[bNV;T8cZNc=V45TVlf^>O<VeZfh6
F6Lo4DAAI7B]f\B<`1Ue[nZl>LB6EciPZ7Q\<IgM2P;67I[PZ<fnedFPqCP_<Im]
g`A_I>54ljo4W6Ge?^=NiY_a@N\3SC8<deCMK<lN6`e`QhS4Pn1fjg]cI_N5E`UQ
DV2bo_cBL?0[en4ki@1Cqa;RPc1q:lT2@3>C:o_9fK2[]mV87j1<_^:1QnHG86^n
;Iq?mj\SSKag_2ZgGM:i08EKRU@l7Q^DEL7GJ6qdDn7`F3C7gCTAX9IISk_NJL95
TaoKXLUF>Dbk`JZN:VWojPJ9fo13_R8]>@SCDEkfoAc:?2W<LA8odNJVdAK\UM[R
2J6Pn5KF3l`jja2JjH6WmIH0G2IYeBgYU2_129YpF2kCm[<BQ\bW<WX>4neGD^BH
OaMoQC1k]Ph3cWO7\^Dj]EjD9k3nkB`]0ZXG^\lU2hb4DQ@@^G8iFF16C=hQ9@Qj
8hdGA1@;2OgR>LmRAhOAl6>7RAVV7Lfokfim`75Lpbdn]Tmbj`<O`67?Fh@V;j;8
m_e5415NOPgf:8hU9IkFn5e=O:O[go=mIO[^mIe^0E6RcpUl1gZQpIiccg_5i2ea
Ie64n\6_a]oPFDD7LGlA6BhnTV6q3kZO`4Q@=dbZVf\4<dn@P9SknjN6]6S68JgZ
d1emkmjNI6=S;g?]O`Fi9DT[O7NWlk=IH_=6R7pm;nJY1V$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DLHRBN(Q, QB, D, CK, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, RB;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
7[C@WSQd5DT^<joMbcOEHhF3R[VK5<\J5l]Ao8ePoXn`\K8bo;S?L6p6ONfE]P2H
S^[nT:;P[B^]^_O=`A`13?R;Y5DM5pan22L7SH<ORSX?Q[MG5Yd^>M\koEeg;Dh\
?VBBB`>]PJlgU`^3P0eL;R`04FY_R8:f<iH;ApOYm4:?pB37i<RDTJRXh>M=R7d_
RVH_3MQq^7R@PMKEZh2^PKH9=]_9HeSPmKJp^6_S7[]1YVcG1DBFNkG5dB]WncFF
L30hd:TdJ`_3QWFA<?AfCh5OmL18LM_6l58>53U=3^p0\i:ln7H\?EEAMU\XN6L6
Dj0Z2Ypi2Qk1W=qe3jaP1p^@m=Q0=:n08OM?dIaPbA26=O3[Z\[246VKlEoeiQkk
@ligZ_J32Pg0WTb\U[jIF13`>RUEJWOfc_G=X8knUDicThNl[1<GkckVkA3Qj??Y
olqGD^K85Xi5fbeKWDQ<Gg47J4n9D0?Tm[`]K:d<NWP2B3kZkCQU[X;]HkXWBoLc
YD2\0NW>>EJeGQ6i_gVXE`MgmlaG[Inh>a;o<6^GK_kZYP:AVp:9Qi?8ScV`c4Bk
K\n@T\7nb_1iJCgMI9B[GXJWeX\Tf^28h;5PcHNbaU:Z]AlXlG?7g6S\`Qb3PReC
RfQ_Kh9cpmT@93d1PXmYMOGkViII2ff9E=BV@=R1g3QLODleBYkgN86N>KOacYnq
c:h?^;Ujhm4Xl5W9IdZOB<;]JT1R<YM_]j9G]=PKdDDfJPG42dnP=OR@CK6c]<TS
CafUn1Q`egV^[BmAJVM\nn41@F9qaS`hkH4=GhHWC1^fojEY>Z\[Kkg``QNcS2TO
Od=fmicgA0;=L69OJWn98<Fg_jOjZ5N]YcCg@5DQPBAKJRYbT`8qW7G]TdGcSm=Y
VgAnLeFnHQ@BLDGSBBFkNm`L@WhOK_Jaeo5Ak<^_S?>_QWCeLKOb<>X5X^<ee\I]
Pm]cIA[5:cG>725dq_VmFkSpn[eQKG?mP^d5@U=M=<F?0FdQ\BJTnXo>CEV@BmpF
Mj?lE=5DYGMloJEE6Cm2EV\67OP<j>KoReqCcCU]ldPC`5`@TjhI]TJ=a0XQdbkh
0?_Xe=X4G0:09IH7G_i8I4d0RnAEaSSdcRVRDAeHmGIbS;@CP:n3iha=]iPNK6>B
HE:D2Jo:Qe1dJU`^TNiLMKEMIm1c>_IVQV5KM\Qb1`3qHHhNEAZgaJ=XI9Qf><UP
AcmCi3HX<bTDIE=CeTK0Q2l1fZb^GQBo;H8gH_E<dJDSgnhY2odi^8aYfhLJ018T
>2AVho8c];OM@I2g9_5TjnP^[[PTPeE2mL5RZ<88Ud?ba=f2RLV<qC7a^>d<D2:N
[T;K2gTYH2c;\6FRM[UB`HO=P^_CpfQ@ALapR5l]5I3PIP37nM^I<^8bL0g[o5a`
`ZXEL\cQle@eIf6q`>KZYiKN_`W[gEdRKmOo3[OXGgM9Ljcm7eKC0P\PEefpK>_g
gmPjK9;JIJbi>IOL0HVJA_RSgTa;^gQ=`K3oYWWI1Bf1UFjO?IZNYeTkjJP@i:H7
RO=;<W<TjSfgJXO;a1;ZC3\T\6k>Ed0:;FJHSY>5_L8>0`?HD;FK^=q_7<9V4p2l
<31gWW=jKN_A^6cm:94_ah8LjbLooaJ>U_=6qFhDNNK^hM2[oGAhnhDcog:?0AB@
7LcaV:DWI7HpUa4K7@gXmESlWg=KHTO1Xi_]7=CXS>Ub?JQbJ87oXHWK3Nfa]4NN
d2N\mYnMnHC;I?1J95@kbmpk=@f_>f:nK`GYQHqck`OV[^@Xh3^Y=?>XnSKG>?5m
oYL90<UTJ_T0C[?YDaiUmM:@@Pl30aW7Kh;4lMB?9jjgE8JmBp>8S9?;9$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DLHRBP(Q, QB, D, CK, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, RB;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
V<NA9SQ:5DT^<3Il;=1jh894EfhD=267mHlIkmS@<UO=YQ2TOa:OM17i\aOdJKWG
@GGqXFH6=25Z1c2U0IX6:[;7;6ID;lk1>UTNSn60REe\B46P4dbBq@CQnI;^QecY
Z3QO@li_]A<V>0ddaQj6b494D;_NP1QqBWd3I?q6l9?@eYBAZ6NFT`cO7FgDDn5[
BpXon3`1WV@2SUaE9HmCmnBcolZmMq;h2NhMY;0Z]Q_mliB9FjPLGkJcRF]N>XEo
cf0?B5HH<fi=;07JlS:RRWUdBXPVRImLbO8lp>]ScC;9pYOM:\6p__AY7j6Vm<Vh
Q2YVI0M5Qm_92bBhDjV4SiYDE^Sn_@XoU<SbEMh6j`YY\lWjjMVoQhA2c_iqCk0n
fE]e=Qa36fVI]4DLWnlBf@cA?ndYGJ3N_G4Om6W03iK4_ZLIjV4Y2Ube<mb:<ZO]
c>_iKgS9c49:JW6B0SoBajPG2Mk\ae;_THER<V>kpC@X2hdc]H44=><K\=GKG>i6
DBiPC4SDaaLkIoTJme;:dHJYRD0fYDY?KHMcPM]\]j_ChmDQYBDAoC8DoNL6DT^?
TMgYD:KVfNb<l4[bGgF4jB]pEVSaP72og``S=EFAQSEOB;@?XMmKWf4jK;_R0VN8
_4_`QbZ:@@=hL61K6cO@iG7U5QS=W_jeY]70WBRiC@n0B:eJlCqNf8Hf@SFKPSWN
U:UJ9cQ]@YbZ;RHc>7a0NUfE2PXcZ26;LF<2?5\?3\iW0OehOAo2[<<5lN<aJ_j9
jDBlm>3Gd_Y2C`pmjfR1T=R?F1m;GEnNK@:91K5D:T2c3kLgndf1hAU@eG^EB?:h
3GfXY`V=K<`O0?hGN6Ff:Inn4G36ko=5nL?bI8pW_JJ?BA>mV<?>EajGBfUVcG5E
QYL9=Oe`Q>gCTHAk>YBiKHa]OJ;AoP_VPBDo6G2=H2c_X;_FDjQ4_j4MIU8aJ;7<
UW5p6ATebDpb2HlMGU\I0^XGi`ghQ[XiP9E4<BVgV9[ViA[:=qfIN4\XeLPGJQ\b
g`E:YHZcm[OeSS1jMbih759MQXHo=mkBY=Nm0BXXR=N[:7O::lA__33Hq`Ojm^HN
:g?LQ79e]H91jTC3l^O@i3EoG]]5pYdZJTTaK[OImCP9iHgAAMFdko7CfO4ogOmQ
?ELZcEY<[W3cHJWYQmdlCC2GOMmBAYbRG=VgDSLg5Ign@8kASdP4QVcWjG[CU?1?
kM]W0e7Ul@cS^WkFYWHkeN[=:UG?CNDS;=E80qmUK>l3DlTSOK=Lb0I`9Ek<J_0=
gcVo]n0\4U_1cH]QM7djH6QL:nLjX^b<5WIX0adg327YMK\<7dnlQU0SlH3Y;<m:
F6[o05LdRa@5Zbm_W69K1m3TY<ZTVn@GC?YF^Vc02W:?Ehq4JG]6\pBn2gjQ=XGn
CE[ggF?h0Ja38M[LZPS1eo;8jQ@[83h>Tpf3Z=onlI<g=_:8nnRN06cOaY1>2KRI
]_ZRhVa<anK<TpRhi>47DO<dC=\=>LVcSgC>PXVO<Vqc9<j^Sb]?iV[D]<[6a_Pd
9@kNWdnIH]?;KW4HVPT`o8Q:[bUHY^CY9S2l8G3FZlA@fX=R`ZMFdPV[ZN_\WL@G
D]<7\LhbO?BlTIS\`[\\cc<JeCdP`aeBSnT\OpachnEmpP0@mVg3g^PC[Zhf5:m>
K5^FfE21JQRQ`dPY:@0qNh2hBcA\=8nN6bK\mD_FHYQS0oKM>OK7\NT4UBpinGl8
4joTW28OKn=o?QC[O:`f4?`VmcP3A\=Shi^Zk<hdilT[a<5:iE@1=S?R0\b\eO2T
8a:A9qj`WW]J98N3TdhKXFOhOkm@Hekng@X[^n\c`_VPPR:ZN]8^5?F\?o<mg34<
Y=JcWJE>mj]c0dQCpE`45T3E$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DLHRBS(Q, QB, D, CK, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK, RB;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
`[AU>SQ:5DT^<h=`7mmVRnqkK2TRK=^5^`\WgEWQB^<oXYVPc]^DMl]e1E[D>UHd
J6eBDc\KT?N=9KHGWOHaYRD4^m6qT?U=LT>`;n`fR]oL7;;`\YW_:2IOXSV6cogd
f@k13aTRab^g`YDXb0jh7QOjKT[;pMC=P_Mp3_l?WNdaENG]7OQk>8eBfF<=`0q7
bJ0\17N7jh00[BLgFmWL_fe=ihqa<onL4FNH85?5kIGU<Q_^0O^bW<[UJ=mk<hCO
R32;eCnWfT>U6gk6VepIC>c@JiYF1[RWWgOdSF_PWBZO^XKCAUjTAUL8XY3h0Im]
Gi=h_SI7^0djjOmHUgW9W3kodqMdnl`_QqM8O^D=qU[C;o2RkBWY>fi8;dTGQAKS
GY]:50oONKV:6MG`5I>?Qh\2g<;d=5\B1Oi_kHCj=_mm1Yd:XG3[lH2[=ljmO10E
_L[JaQ547?V7T_5eo[YK`p4>Jk7]V=Z?oQK9_B^\]EQKU7nHBn9aD^:UNAf22DT`
ojSH?UBaQVe?cj[b^:QDnS>T3;S]hB8OMAkg2CH?UYFdH>b0\aIb_Bh[hQWC<9Hf
IfVipXFljOTc1F7V:6\B5Rgd<ehF^Qd8b7ZlJkMJkDoHB_Aa88W1`Bkk?eO<]<:d
^GiFn17Pc\WUo;KOWhf:c\@NHeHNn@SqOgEM:doCT>@M88KXYj8DJF0P>FM[3K8_
J_=SGc6G[^kBJK89l0HhM55HHkica[<gBa:>IC[[CYBQDW1YmLPH]c3>[H9p@4<_
8<`lC7?eFiT1<C6Q9mnMaP`;:=RDgh0[gGj=e@^Xb\;][ZACaS\dOflXRT3_^39:
]L_c?Ch`01O0l[LK>YLpT:nfJVUMGR[XRo3fS2:TUcG9DOROIJVG1?a3JNnBHaTh
fZB9om6V?ikqS<\LfdcLQZ?V;kAVMd=NW9070H^gfJ7]BmEQcC;ChlUn:0eSdJJ1
2MN3i:6f_fCG9L^^E:B:@3Lmc49PF0Ke==bag?LCqG1d2H4pHGYic;=1;UZclQ^b
8]Sd3aGeBoZIETZQhcK3fbp5R6ooPT=9K6\cFKacZHO5_P9[_S8WY91BE`qNIa:l
?NQm;JK4L9ojFW26MI:`NQ6hfL]C3PfiToNGI10bYY]l3Z@D=9HnmQd6]\bdTg^l
SlI^QbiYFf3m^moMTWEHllXYd[KL=n8VQebl[iGB6eQdVAB@^@H@n`]3i2Ti9NkE
cBiq>49O:[0bUY\h?7f\ZB>0>cDT>oFIGd=9Y2eQVkCbYP`kWkYC60:Y^@GnUjTZ
2gWEIF]>[dAKk0jeT=\JEWOA2T]:@?;>03T\05U^_g?gBRLMjl>l\iObbXN^1h[l
1OU]`U2Y^Ok3]McTpSGB7SQpX4M^6GYI\OV:kJA0c6e32NcQ9Rm]k@Q9L396WmN9
bnDpSU^BdEQG\gC9cYma?YeW@EF`UoFJQ`?@Q6<7jJf@Go9pl[KfTMl]OkaWG:XQ
cN9=9R7g3JpCWXYBIW@4_e>5Z>@;Do@A6An>0ccMDLkFha]mm<YdD\3K^JBPj333
9m^G_d^^Jn5bI1hncAZRVYDPYM@lOIcmo^LedM;OamOEGLDY\1cSHC4KT\AUK=DF
G]o=lp]Gb6I?pLVDm]E]]YDASBCJ6d<?8lIa9geXPP33AOo5LIWq<5DJk:DTMoHC
QQDZUndRe6SWcXh^d^KAM^[aGopQ_2?f8BJhBEV^XL\8LhhZK:B\5ZRSm0\Qj9MD
Qf4Lbfo^Y>6oX35=hWhaI^G<1UA^1HS`S]jh=paXj1^bVRa=MCHhVZ7n\GW2m2kV
7kBBbO@h]4a@72aO2BJBbc`JDX5n9A3>T>oY6`8gVF_PnMfnpRUkfeK7$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module DLHS(Q, QB, D, CK);
   reg flag; // Notifier flag
   output Q, QB;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
?YF7XSQH5DT^<?;l9]K[BKlQJ[ghAh0^W1hpLI=T;eMQ1\WaUm0@]W5c6LJXX:`h
oZXq]<YXn7=VBaUeLTLq@Nc<4Mqdkfh1j1M@Pfoc?`;TV59APIgF5pDkYb?EXMhD
\fRR]=Ghl9RIVX:mbp6M<TWIdX7SI?9QTUGLAEFL;`aDMcfjcWE:g`\j1ncP^8kN
Y4E;5BUj^_^ZR:`N_36D]\qUJncIcYT0K9]bIXAi81LEO@;VI?8hl?^jQoZaAiFP
N18_[cXR75YXD4cV`l?FMqMOJ^9e=qSPaDZBq7mNI6i0ZG8;@Le5>8^lKMg4BTb4
2YZ0oA<N=7JFME];dXB7BKmle^8Wc31KEX>3NgS6dmV:;`VCgQFN[:]Gd=OYBJ]4
j1R=F[BM994MX3GClqES85P\8\<9;l]JZUQiSJo`l\Tj>9Y37JVg2dYT7<@mdem;
2ca]:Z?c=kM3R88@fBg4\MBMYM8cXXW>jX\6[R:cYcQhMXPLGg4aVmW5X;Q0go8d
q5\2f=S;bNl[Q>G_k[_iObi\3g0PW8l`OE_=me<2JgeACQg2<m9jk?P3KlM\;ijo
Kn8jWe1een]=H]0<A\[U\0Sq<6Fkgd9d\Al;aUK8Si@<lMTj?dY0[g9@AY3ol<>L
oZM12nHZK6MI6`lQAJ^N<Se@L05LV8?3iU@E0SfmgUa[m<?5[K0pg?SGinpkTH;D
MdRjaZN=SVGR[:hcVg3^m:E4C5D7:2cDiiWc7R3=3B4_;EKPWqG^8JRc\BFEWE75
0lJ5U>iCnUmC:hOc8Icb9KSJpUM<WZacNWWFIV1>egSRbf2d^ESF2=0]1YZZpReO
PFVWRLQKWZAY6L4IYTc^13Y^WZFK\`DGjTlEi[k\7E`S:3d]enE]:lC7eX0]J[GJ
6XAFdkk\[9HMJ<KU]^7IF1VHPZFaHk^O3dgC2_8U]lG48J8D;W9VcTWXKp]=SYJ?
d]QQN4hIQ4BG@AKnUNnTZLG?VUWZ`9G9_iP64Wh_VUm3SdL1W7A01o2WT0Fh]iAn
Q0XL5^M<UR5Y?9e6GmXZVMbPCgTZiP\TIH<44IS0hW149?XQ8oYF40DLkb]bFTp>
hdA^QqlK=KAIL4QmB;AY=E<6QiWFnT>SCF;S2?b]ID0dq>2AHe2]CXdX8GOcBdMZ
S4YdV2M6aZcVe>=EcXN?W:7LPdCGo?W9m20WYkfkHYZ_oXjJRB=WgSJq8l1IEDCq
ahKiJc7[81X_ejbhabahlPLb$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FA1(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;

//Function Block
`protected
Po2HbSQ:5DT^<YERS0\^m@mUDQGkR^Pbce:Ci;<RX\i??HnWq]RKbiJHdkRKVZ\U
`2=JD_GGIDEmmdE=PYZFe:Pc`KhHWXdefdAES5:NK>7KVci7[qZTT`^L@9S]f@KW
PBO\CoPS8W1mkDZSle;CI5XnBI>CIG1R;A`Q;Zp;Gme:?p1i:g\^E`0F3OGPH4_M
hc_iOb\J4`:?p4]J[D9F:nO9Gj8d8`9Q81>06T<n:?Y=qBHYVg91TA0]XX29]Kn]
1Pj<iI<a;e?TpYn36dYD?:PiRHkTinQ3HG?kDN>TRJSOTBk`:fLqob\LJUH_@`B@
M3LmN>:kNMUTl4V@J[Oc6JqbO^5jQ8q1MiJ4?p1MaHkfk<UEJ@bPQI5MF5o<a1MU
?OaiaU<laPS>FVQ^CE<UjcFMHBFLZ`f=e]bG\?j3I8:67E4bQ;]9<?Eoo1PH6<CE
6TCXe?a8AeY609akm<3YE9h;BN34NMNZkp=majUD1kb9`d06=nbhq<d5nQU1VL88
O>?bG:9<SXNN;TJa9TV0n8_jI>4B7oNgQJE6k[X1Mm5:eV0j4nG8OEh<2JMg1?;S
P0i3IY:?j6JY8^`5<Vah6mlGEU8F255lB>h:Q=3oP`;hCi=Kp5fhZY]oU?mgcP_9
hhG\NZZm[FaeD>:XNJAFFYgS^cm<RjFIO<JM]=?NK:bfHnAc00LM[Lo]le95[;ZG
WIOO>FXIToOK><S@]3AUl;1PS>cTI>>>7jN9`^Pf;]c`qdbhcJnWZ`?jmTcnJTHE
PQhM2Ucm:k]o6O<;]^_lAdEB]>CJhI23^8FlgC;_8:HV5mN6TOg9gCe[8A5]Wk0=
S\MQaeE9HC8\9fbU9CCF^FPQGSSL=DIFeiEISfSLpUai?HU@Ie[3QB6ZiKYN=>IU
9C>QS3PF`XP28NgjPiloO3VXbA`7l3@EhCUL?7VFB@QDiBEDl1]S3:1ANlV2Fojj
2fT7Eq[O>KXiaAWNP=`XR7naB=jTVkJ6QK58`>XkKc12Y>HT_\9E6eL@<8cPQJe@
G?B9U`eRN=V2RmJ<6R:43=n\VFc7U`mmH92WQ96HWo>2f9nY=eIBM7KGBBUkjZpS
mWYaAjPL@<VnJaT?];]GK5dM4a0^K9W`a`kBN<`aJ[aYbTPB:IAgFReWQd40n7dj
BfehXh1\\>aa^LnkKoWDj]8b]b3d5NHZBJidNoTkC13c[<Mod?7PkG9q]1nN01Rj
3ImdUP\\JcMXU6nB\Y7mYOk:FjQ0LAS^>N;UinjHcOlVHFi3ZOLcO?b@JKo\OYJN
1A81VE_W[\CiP8nhWJpce>TT[B;iKA`aOnTiVVglBNUB8<edOM@?T5JdEbBbFjd=
D53EJ8<9R_Z4:>QZ[g2U6d@QYX6aGbSHNBSS4Ug?OFEQkL]\aa6D1b^PaXcQ;7@n
]^=WZf>l1HHe_4pJVd8[dM1YU00DT0=9l]OJKn2O[KUdM]MTm>IhgG^?ZVOD^1lG
Sm99TS7O4cgc:0Nc4oK<J;\ej4NCFf@RJO?0n7:Jl70@ddgMCPn9L\E=RYRl;nJ]
`O3nV;=of5qLCX6X2k6`f?ef7`S=old9S3o=>24Le[S3I=iUN8hD_8df1T<Lh]7p
1QmfXPd5ZBS54<Tb>28EnF3EF6KDa2a5M:fh_P4Zo7fLRKb_A?2\3n3\blhMLNPa
QhfgC5CBf01PB\bkJm?JEm33<1>g1finaZ=VXdB9\clYDh^afSQ[^OBE6P4pi32=
OOAnTloL`OPn^VBFDMSQ>F]X@O=jL<>eQLB3c=YB>8O:QX?803ENWbC[gdgBG1X4
L_nI9l[Ij6>537>>agj\ORMmUoLHLc?n7YWo`?b_ajPP0]Uo[]GnRObqnkf=?0]j
m9KGT8FQ2_YY[R3;Pi6RJbAL^<7?QGD4OO;j[ibCb7aY;?iRnWS5TmfcWF>=B=;D
S4?aW6NgeNK9ID5`h\?Zq`OMV?YW`2]hgf4<_:bn\=h2R>]fMBenMB]Gd1fn^`MQ
ogQBgKH@W5iT3mkkmJ3H665c[k0KXcCDj[J24kLkFQUoS>4<UO>>iZ;HS\fS=Y5`
lj>?OdcCUl10opnU5:<nm7XB<a4cQ]mN9Dkg0n1mJ41F8X@<167QM2l6dRlT419g
E=1<FPK>j_IiXQ[X<j[e2PdDfBBZYAAS_hF\OeYQ?l0HoX?cjNYQ9PSWom87\;d?
gZW`0Qqc=Y@8BJ`FcE;XfeFDH>h_0A^>ebUNFZMWhN574:og[H\@QRdIB_:9;CJ]
hGUAEiddP;TSR6a6QL<Zl0MZURLnmifQVp8ha9Ho]_PK6FMkAKZbHZCJI<_9R[FU
bY<_20FVJ7ZRHBY2Jh?kMhR2\ICddhSH<^89bA5\Se;hiR^D]CCEBe7LFNF@S8]B
bAZJWSSgKd^PMGgZZkP21pAKJL[OEUVT<^acC]3PF@ba[nMP<XYW<Fl7VLiFVf:9
1Fqm4kDLk^P6bHDC_fimZ5g2Lo1Rc_nPYTi2D;XkaeOYNOKYQ9HFiMh6]<TPhPeT
cM8mjM79?XhLdKam`AV7>d1Y1oAg:Y`VWT:7n\UebLJFT2[cbIJ7?Bp?\ZjTUi:G
46b[?lWSWInT17<HlR@YFiM[UlVZU2ejnaRWi>\U[]SHm`MaPACff2P?L6Q2J^c7
C^K;S0OL0NQ><GfXP9KUVibRg<QOnW6JJ3Om3:gkVHp9DK@TOYaQYDJejmk9Dh^Q
nd_<oXCRSULIm@5HN>aPanZ^XAW=NAP=`kQ>:N:hkZK9k=@VLTV9`8LNLonb5]69
d_S]5;k@0UYZ<KPSZ0lgU7NMn1IPgCpGN5d`6C2JHeD7aJgN`jnQDajMn@n>IlF3
IkViMP2=m?lbX]VCEX^;330;_Y;`[[`GPS>:P>iaSkEX@3bJT@aABpEE5O]R6JbS
RIEP>HGZlCnH[PoO_Q=EiEC@kD\AI@lL\O_5Z1NX8aD9S;F^LU:LWbeC>m^[Hlo0
oG43Lg^oLldg2[DnED2RmL]j]VnA]:=joN3JW_^J<C]jMiq6giI3a>M]b=HP@TjE
8gg2YN27OIlZCb46]Q`7SSBiC=jRN@Q_]=Iim^CP<f6cK2cHhNlP[:i7NVAc1IA@
Ef3HHJQCeQ_YjZX9OmR[S80H`lXeVLgZ7]NAFa0q1XjTT=h<UFDkK?gDGmJO`<3Y
h5JF[k4IK5E6<JcQd9D<aAgNM\nLBkDKH8[QQ[RbP38ciAD9_T\1E4@B_A\EHMAa
UBRph5hLi2p6h2IVX=XX16o7UI_eRTNpWTFjSLA$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FA1P(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;

//Function Block
`protected
IaiXJSQd5DT^<=?R<8:_@=4AAj9Rmnm\7DcDj6Eg2ZeP1G3iFULWZjo4GB<>9oqL
S7]`Q5EeOd[:[_4L5An?aGjQ[9ZaW:gM\WI<MNHA29=VR]qod4:CBhVR3KXTWEBJ
c:iB40:nU`ep19@XaDq[`IeH>JB:YBaFHU7dli[VM3YXek0eQp:L@KMeC>Z0fAmV
XAL8l\\:K\9;EVNeGpCa:oY01g1o45I_`2Jn8;A4JC\n^V>\XqHR?ikK?b6Ch_P7
]Fgdnc857@P`b:M8NfDaLfd`q9H\7]U7G:e6Kfd]XH4o1Q[^=jha6]`KT0Hq3V^9
3`SNLfOBe;9LHb[=Z:1a2EVUadmXKol<Blf1j9qYCF1PE_qSl4IF<qk:AnLBiFme
\7R5lhCUEM1NLBUf8:CeVETOil0\U]7ocNW@3cW\<=T\VCJFJGk>I9XE@M]NC5PN
lfWSWFJ;>Qn3d3ZnVW=Z@aYFaH=bGG[RAbGNldAM]E3K=I=k`qPJ_Gc1[]?iVH_I
alfX0D`HSRW[1Y<QY?O;DET2e<Eo7[JU`SkB>`\LWom_q3oS:KbBea6358SQoAOO
J6c1bWZ=__j8d1D\JRBmIDlAMZVIbbW=QYcB:;X2cO;9fBAARY7=]DbkCHo5PlK`
X3`5J9PEh[C`lgc`Sf7CXl4aK4672`@2MAn4_Ac3p6l1`104]?Y`U];4n2bLVd`K
_8T7G5V;`6JB[1KdlL[9kOAgINZi]24ZF^eF9dCi3afGGXaVICJRD6=96ae^3All
@KiZ1JMY@LO8PQT61=Q3d_l_0aJmAUEmf4bQpaHRLZSg4?Fod3O3BSi:ET8nBAbc
QkNE7:;E@UckZKS:<50S\X3Qm=<RBRfgRZT4^la?LG0?lb<E41b@KjcEj=@594^U
3eJ>^7>\>SBdYIZ8X8aV0V@OI\`[IK6HpmhMBS0MULZI2AEKOjSqA98`EmC_o2le
@GoV<7O;I88aB<MC5XJ=iVhmN\RE0I7XDCI=K@hNYdNK>EV[[j4?S1VcmHEO6WG[
;eEWk9E\7SUah5@>q[`aH[a0mI4^8o^Rob_KKnW_4>?00:5_OaBUlgS>jZVh3Mj`
i^n6GnH8B0a=;[AW93@DH4OmFcD68NGn?N8o47iA8PHIQ`>=GjmWQTSLGg_U_C`S
d@hoJmJbTpd]nGbb6J8_WG:g_oG6M5BV?\kBoC<bi@l8W6Qj?\_b1m?N\0nQ7aF;
RGile`2CLO5IR^DO`[ILMQ<Z\l1B<4AFAcn:;B\89;Ul]M5jNcZ4F`cVA=oM8:KU
9]pP01aX2^RoZZMkbCS6EJ5V1Ho=Q:FhGV38YKolZ>^KHb0OOCYBnP6]?gAO=[hU
3goEcP_1ZQak21R>ne]T50iJj3fe\qgc1ehbbY;GLRd8[a@71m0NR]gY\]fQZ150
4cL^P?jJ?<21i@_`LnnXP@b6<C4XUIdJbPXk1DgfS@\HD?UUGmbf2YkNKiTfHN?;
BT:V0JWOo^PB57\k4idIEkS^gqB<fHDV8o0UPCf>IUj8DNMO7cB7ebYojKKjbhma
ZUUIgU[hSil];AM>B8XH=X7W`eT]:mPe0HQlTPLYaB=V5dLeDZCE0V??>AU;JY:c
Tdn0^<1lJCSkMGHhNLiaYqGehfK_eH2c73fRjn3c@ZhK<<Y3Pko?aIXXUB2nJGQN
Lk1l]ba8GY4fN=6U03]AhbGLDW6MafnQ]SR`RWIGQEPKOf_[`NXV3kQeR\H4SfFh
=jd374Mm3BfOTNI2JpCMHA0]Wg?XoOaMh@_WXh68^aII>4Ga86T=0UnTh7e:GHaP
U^8>o^5gB5;`\8P;i_6UKlBL68hKO02=5Mk9;XZUC_]Ld1fCdPWUQRQL_fc>mIHe
j0O5[Xiah\BgbqCo^o4]igDLC0U?LaF[f2fnYfCh94gcO?2j^VO540JlXi>Pf<^C
iYSc:3H26JLKEAmgj;1Y066X95kmV82];87\Ci8]hCp^_Q6BbAJ4L5UgS75gJ[S=
;iZ<b9h[FelOQA<lM6bXR1pac7?QlOeC<67Ga\7OY<JRdS6dInH\@XSH?V=PQGb6
S;=NFIee73P@42cnJ6QMYhd;f2A3Mf7dLSE2j79<JO^?Wn:lL_RAc8ECYa5FQNbM
\B53@Q9fFLUU;<QqD[IMif6A]G;YG3LITbnZH\:hj0BFa8BbEHd;]31<e1m[<XWc
kYTZAjAVS3S9_e9V?6\j2`9Zc\f@N9CokC3:R5Sl=U6Nb3YW@4[Z43e=ii]^k830
H0Gj35]>pg<FlbiUl:3]SXCZ\a:PLni[>8[gnlgZ_1M9DC_R2g_Gd:5QWSE0ZLcM
@afjWYT_7^;BR<Y5I]B<8T\aCdBgg`XSNb=p7[RIZooFPBk6o[i@>Z5X:BP94o9o
b`S3;A0ZV=cj5g5M4m3i2M6aZcVeA8EDXN?WBhkGWiBSVLSETFW=kMFH8P71RY=@
G1bV1SXa>Cm^nZH?UOKOG5OO@4[p6>`O8hY=dY_8Z9_NHPF7lk3D>;::GI<Ei>;l
K^mm5NC3Be\m>K<nK@W:ic0F4?7>Vd\U0DHQVhLD9EPFhAY@@cOFEl2d:iAB]QdS
DlUOZ7M:E=9dZ3XURf:pHHhN2V?\THO_oM^400kL22\XReeWa7AekKDRhlTFk:]C
B4@c=?4^fVAj6IE@8\H;5KUXRMjNaJSKZg9gBK3_j6QBCLYI][Q5RUD>lZcjaHP3
:kTf=7E_LH7qG<8172j7CW^?m`9X<9I=N;FD_J?L<5E1n1R1m]Tb^IRnbgU?d?mL
ZO93M>QOn1=I\O1J<0H^n[e[DCD\ZSmL@FMCNN1HQ_IVB?RB19=[F[B2HVg8Z6hj
a_8pHg5E=>gOo1MU8FkaiBYel:4dbeo^OlRh2_MFF3ZcHJLNG=]jg4<PU_cW]1i]
K>Z5Zd:A_E]BbO]BMg]Gi\TL^Em4lbpYFLGjDD`V6l3mA^>`PFF;1?P_]Z<KYmi<
>L_@l?D7T9_IL;;E505?cQe@7XG=d9\X=Pi?JGPW8eQM\\gc?RhZMB2edO3mgV?P
mmQ@lEG]b2lN_VL6:KHmR2YpdAE[36]]j^mCO[TE`^BoHjF^ne=L[Yb9AKAW>Zeb
Za;pLWT:V?M6mPBkZ7PedDYARFe_E=3G23;_?oChZ<WjMY?@3M<eZZ_7W:=SlH[[
dIo>dl><nA>VkCggReW>WL6]@NkbZRHR;SO;KElAZ<H?b7j=^GFH3VBe;A8fqdXE
F<k]bG79KeZ02WiEH7Yi[VbBm[B5_R^WMNY0AhheDR>EQEZU`a92@XO@1BQf0T?T
5H^B:NiCEal=3:XM;WhA?Q]]p^CIhLIplRQ[ieg$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FA1S(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;

//Function Block
`protected
d<BKBSQ:5DT^<6h:^CeUo3ETS5[XVl=7bgCKaWkYcAL1Ub6DY6Fk`P5E?eW^UE@8
ekW>iD0E_eILp89C\XlA;>2`NLSkI;e@5UY><732J@gA50D16O52>R5o6SS@M3fP
3T@Q]b4h1ibJH_PAp1n:BL[17YgET7RJljL?b:J;el=`Yh5d6Y\P\kI>Go?7n_n1
TNQnM461S:WAk5L3O]GjQTE5plgA>\4p5iGkNmT1BiFlFFNYPlf9JC6B0=T>`nq2
RENckom8I@A_O@J8Ug3834>j\[6>:=qC>i35ZVTIV:<Z0=;7PB@8G;5KgJ1L0<pH
HFgol_9c8lbgK9Uadh=97U:dOjh35\dQ`MLPNNGdQ?Vb17b:<N0OfUiH\KXPQH[l
3Q1mPq`JD91_egheT0RmBo3IJRh0GlH:T?@l]2FkAd8?q?6k@GILBQG48;e]:WG\
`E<Xd3kY5XfFh\`qJC_lXm[qVRC[AmqnF]@AC3?9Db:kbTEi@PhB5[m4FOoj2G^\
3Z8onTJ0YaDA_kSC=B5QiRcPNK>fPE7J=1B4hh2H0ME7KGl<Ijfa9g[V]E5e@_do
KIhD;YC@>oBcQ46HhfOU;giYo^p2X9eAInD:I4JoBkXh[ZaU6LeU=Fgn6<_c3<eM
6ZE9jBg>AbKNDQBT:6lH`PfM7`>9g4Kac2><naQY7cZIW5PD6]V^^jb3nGZme<\c
mUCC1^li>0<]l]W5LlqG[@Kg;PB;B@Jgg[@:@2hYLZXAU<=_3WmWVPZoXMIb3L5@
Q6nUIVRQF5`@GipXJbfZGN\8\7QR4C8Q81oFLHL>FR70fN@dRTZ2\^ijT6>Gf0Mn
R=S23ZkgfkmJI6UjmjAb:oon9c:?j^?<;14[L[V5Z3`J:3ob^TETV72]M8aH;f1:
Xo5Cm^q9]]`6;KZ9[L2HgA;OP]\QTUB>`7K2T>UT9ZlI63ECiB0F3k6aZQJ4Rk_<
3^Z0IdoP`7j9B8c5Z2dmLN3SCI8cj6GJoFNe<G4Mn8B\L`QbIUC];>0GoNMJ[j7K
L8qT8WW>@4@4J0j_M\FS>P`o9bSDN7:cC;LHBO]:EnC;J2UoNIE\BOZXEkl:?c3o
MYN[k@3VVk1g64S<MGETQ5Q4PCe?87ipU3VR\fcad==ac;QUG[3>oDo[kfB_CY:1
KgU^e]9NEEen0I6g`0MdCkZABmi9KIQae0Pk\]@\NLJI1U8BWUQ^4=e6HfJi2IX_
\43Fo]d3:GUn@kAblJQo_G[npAaITJO^on1=;fiRX\MfA\0gJlfk>3@]TMY7ZHdK
a6@kKVPTH@1A>?3OoL_dioNh5TZo;]e\g2l\K^lD\j1`cGB\E_Kob54U0>PUQ<dk
Di^W[Pg\_G0jmEU3Epjb3;`Lfa]m;hk2VfHQ?FPFN<Y5L6Ci4chnO:;944=^eh3l
G\?H`FHHW[\mlFpd^WYICjJ`JLlfP;^f\FjQdaaXJjfiUC]mATV7_]Y7nM[kXO4Z
>P=mMVRmc0KHO4MI2iZ97IEVQ9<7KhM8UWfk]\7O8qndZQ4XTTJHnQ0I<dj;L<Zk
6VXC4QdoSTRRlJnj@Y?6k>R;nd4O3d8@EVoGgP7jDoZ2Z_>C2oH7bI;\TDnA]Qd8
:F=T2bAE>SV>lmFPTa@Ei_<59>;iAXo\ip8]EhHfY8f1Ta0`8;U@jj9XiX24oh^K
nklLaYVDPYC:G2F6BLLdGi[4CZa61cE[cQB9QdkUDNg;G3_o@ZeoShkW?o0_7HXT
66@mR1J_RWPjgmXfJ^Ga@<IA>FEAYp>Ma220\<Xm08hC<kgl4^n;CTZV6Gb8eHkX
k;\7GR_B1eiCjgm3XbmS0JJCdBLASIRd6:ZMcfm<e`NI4OGe8L^_W4`11C@hNZKP
do]B]fOP?UCY?A[mZH_LKK13:pNE0G36HWmNHT3EecKdGJK33n<S]DR4AAqZ6PgZ
>Xm71Bf2fMD\[heaDmPYJYgk2\V^d2Ti5cT^EEVKneYY43FhC1lZficn>Q;gZei4
j>P3SF]40QK>O6XmD=J\5md:6]CUV2bRWLCl]i`gl=kUjZH@gWqFH\;c;Xd>;M\3
;?\2<kIDS:@=HI0:ilm[b;XZ;VhiYlUnAj2jmO@nC6\U5H:TMZ^W?9C\f99;38U`
gLCQ^gm1kmFqTi^_j9nDlF_KKIK=2kJ>Qc3IB:@9>Lh0m]falRVOoibNnJZ07J<g
^FQH@<>[0[RG\G2\g5SUS3`mnJN]Un^oB6;9]HeLP0cQki4fORf[R`[3O^jfeRYc
`NPlpd9YAS762m^W1B79P3TV9a7S0ohl<I^k34mc]4Cl1UJj<9l]@6Ub3JQjHR\X
0KB=1hbk?U4^3g@\B5JELO3LPhg2WRIQN>>o]WAd27CQJRcE@klYjGc6aB^5Yp02
C^?X\Bb4F8j04=^@9JaHNeEDPWPa2I]VLV\@dG1]9A]>?g7V5B[2<4TJ9[_74[5X
=2L6Y^J4;[IiD[HNbUHP^f[hqEE6^HMa\JhKieJn9ZGHM[o2CCnM9Dh3Dk^`Y5:2
HE7>VNB=BkbfJELQlARVj2]2I@l39MnmD^XLcYHYL>^6=;baU=n09U5IaQ@Q8f0P
`OL:[J?SiNSZOklVbX?bqCVZn3S\ciblcGEi_Dm[J@bOKn_YZUooDOG:_eH5I:NW
BR:\5UK_\3>IK@k`lJZDF70Gh<G>PARL3\9NL021a?_B\O_WP3ER3AB6ZN>f67X`
n]BIDNKGo9V_Xi[7qlL3MF1I9HL`Oj[A_QLl0=hm>l`2G[;DA[U[PiICPLG]PCN`
_W57XD68eCCBXWLd3KHalTo_3iS4Vo0>[YcU:4Y=jQKnM?kBmjB[XO]VI7kSJC19
hPM;:A=8pFh:Sa@?Mf]kh11]O856jinmmAX[k?Q]QBRj8k\;Ei^BEm>h>SDm40:C
c=Kh\J>bNCP>P?EhLPAA1BHH=KG3AQm8[LAfJn]E4Sfj5fndL:2YcRL@<5Vd\CU3
p=STTU^fkdBF[Zj[XaY:TO:L49Ue`RG0gZmATq:5FmJI<]YZEgZ9iVDV;PK7nGVh
=H@D\44fXWjR;4;?YNP_`YN?<PQbd_g8HaliRfa0OoAcfDjlLo:l7iffd26FRbYH
q8lF>BZnG=kh_Q`[U=dOOga8AWU=2cgoA=d<=OIVIINSTUbkO:B:;C7Yg6T`LdmM
A<MB0LOKTo_jQ;jf4]8D4gCN:VC@0YK<V16Fn]IMEe@R5M43_0n37^Q2MpWe[V8J
UeISo6J9HICBIdTCY<mJEZ`khi_nf6>dC]WQoiS^;W9;FRkeHJAPi7LUWfDi04OS
ZUoF_e;D^Ui2`47e;=VFYB8C;O55Mc2dd<8XO6?F1F]E60F3jZpCSWT7LI28eJi1
CMXeZT06KeJNP7]jG?BRdD<V4bY8lfik9hQeLnf0bDIoilCQ[ETbe_BT9R6jZhBC
n>81`Uno1gi>K1p5J=KZ]p2o\UY:7$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FA1T(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;

//Function Block
`protected
7AAD:SQd5DT^<4DYVX0517dIB5Z1[=pV`^]:X^j?Kj>YNjb4J5KUThHVST?NfibW
1Lb@leW]2N6lQmB<AXFpk@5<P<NTXk7<gaW70NCS060oTKW?b0qUYGf;=p7e?KTM
I8l3Tk1GVYTLhJ=bb@edW6b:qL2JXjlSHKUWFi7S[dI16:<4j?>3nJ=GpW:8[XB8
lbTi[PH:Jc<dc^6QL@M^QGI3qRmL_KJf=9dBTfWUcag^U[[7UnB0EXXa:Pj@6Jop
YP[]KS8=]SFggGAgjV[hH:4;e\l;JAE]8jpQmJHFL5lmSgA4d6NQ;:c1:E7>OY?p
VLZPRD`pUL8?i1pY_7I`QJ86U_CeD\SWAjU_d0G5`2`iH]gF1`h6[RAcgJImWVhM
ho^25Bc2YhHABe02PWUBlk[R[9`K\`2d=lOQaml>_Rl>Q[RVdnf[RMcbc<ZgGVlZ
cKPPJCLIN;p?R<NSA[hJ[;Xo2CfiOWC<@[^Woa]KGHdcZ:aMhkgRmYTlj@@<ikF3
jkh:SX3ZCK>YHCMo0Q8GNAIb6d;MoA\oYc^oS=bI?JL3VE[V]PJ:554LW\VlGX[b
dBJmYlqmVToRN0i9EOa@BAFBi^5An9:CS2ej52j4UaBkJKaD1>PHXG;?X3GQfIIT
Z;OAQ@o\jg1VWOO1K5b\bV;F4i>^lWN@0df6<EBD:5OI\OAEdm`KUW8\Xed0@F20
>ipQn<2dgO@:dGiK_7U0IT9<K^]5P8<n4EG4SS2dHC5oF]mqL0J9@]e\NlQ\29]Q
QG\NjNTQ53A6dOLR2kE4eTj7Z8dJoCE`0BUPKgi>o:QaNc=`;o6FBd;P^Q6>1noD
WhAl9<d>^O^?jo3M6P?@m9`Db@X?J6]@OWCYJEV7>CLpDQ<::9_@`liH>V`43l0O
f`\jSI;R0U`^H_Y\>:NlQQHIZeI>c2JVTnn812fhPYU`BeHJlLmVkKffk9`<TK90
WQ=UC=>Pq5E^n<T^IW=4>EE1SlY;iX3M2oiXo3^i7K_]nkL[IjmOh9dF7J1XG^@B
U\;NlacAlVF@\]6HTak[GL5_lD?k@1_6P8i=_>BkBF8TKa_EWMHdbfnh4Q41c3><
Gc<`:qKKmgZkR\_DggF<`fDQRNf5`RffJ5RGD9kFlh`oNGnOnkGGEkhIlL6_BePk
2<<MdlXBW`S7aZM<DD\oRnL:N[g1e42f2IP^=A9S?eP\6:eZ=B`kSL=JY7Gng@AY
H[p^0K>Dio8@hQ819g_HdPVRVHl2gBi_U?GRVK:DR<Ldh<Y9nQeaoS:F[RWB[ClP
Z:?5;j:0^5hgM8S66USj74caBZXKeXi_6pbM5naTa1b^VOg3UJ23fnjOhodjO7:Z
F6:hK^C]90[63\]QRCXn@F6T4nim3b7\CoNQG<5DTEFZf6I[BZc8a\2KY7@FQYk^
2iDTlElcnKkn8h^]<03lFk[7[J?j3p<QT2G\8C62;A>Ca`9XRk\lH:N\>d`;aDpN
b=Z]UNIXom@Z>?_Y:<i9Y@k@5>c]IE5^<<J[GJ=gT?LR\3]P5AT<`7Z7;P3]@R:]
_97DU=:=gP\Elh^0klgCUEG=:8[5Ene7]o9P9ZGQR9m43Sh??]:n_O@F2\q3iTHF
@Wo;Di0J98cKXL`e2CZ]_3`GQo7iJQ4R@b^KV<\<MA>^oTSO3nKK9KZgT>:fB_\e
HdTlW?9><L4BV5JC``J_i025KFEf_AQL5X[AB@IOIoJNHB2JOCMH;Ip21ULaWZPH
cUV3mS<Kdb1nnnFAY84B8F0`79`P`j;B<RJE?^`OfSKYlATChI3O[b5Z0A0dhmHU
;TM5k1NNo3;@2[CaL^WY5V`189IFfTIdHjo:o:enAiRP@OBX77p89c<H5[SoXGm[
TX4X<ncWeo4Eo<6b>WMmJpcO9XmlXL;D7jN[oY@3nfH;^J;4mI0If0GThSgZm@QC
LbenS4i@jM<aZ@^9MLB0nFBEf9LN=X=Z:0G9C=Gmd7ic6k\9H_p_16WAKc[P4ea3
[62OFFZk648OS]@fbBVoN`GlMHLEa<Mkl95VbKB[@HXgl8D6:SihYeE_\T9Yba2k
1V=\5mSg4A1ES]\=e<]F0mg^DbGP4]i:?nGYa@7m3::7N\Sp5AIT:M`j89<aEL1e
kOMeI6kiKcTa6KadK][j03`VZc>HMe=68\;>E3QQ`fn];1anO^N]^OUaAbl=1X0<
3h[69We97cWCAR7ThR=iWET7c1V5[Gd4IYGn`XNZFJ]:p9SCO6@SO9g[Wf=B6Mgi
Xc^n\DmQ`17fm@A[fgjb]2ZDDRAVRJ@1W:FLe8U<<5^b^G6B<4HG[4=i\k4PO>km
J3M?fkWL_V4q3<^af5L[M^7S=E2MN3alceVbPbQ^ddH0HAW9nCHQnIh;\LJj^]hF
ZkPmM<[nF4OfkTS`_C41nNC12Ig`LSZKjVNdVb??bmAhS]lIXSND6]oakn3d:6N1
N?``hGUq_mT7f?K4U^[7UhemS_=`EoV3o`CPbDBfGjU5?PnfUHm;<F@Ne\gMH2Ui
OQ`[4X:1CDfbfgcSDb0AeeZh<GYI<DGYH`CIJXe^<XGePjE_>ZidYd5oA:H@J3`K
o@_qKG<cPQZNoc_@FP<RGM>XhS?\WG0;3YX`QNUUE=ahMh>;DLBd=iD4I@J9[dMD
Og2WhnFV@Dec2T<2<`VIeDUAXVmdf2Q;EfHbCNUHY>mB[hY?PoLHMIZK7L>q87IK
]Lm^j:dGhJD54egndS`nJ898SN3oddVZQ[`eZ:bcScf[[>lfRME6IUCQVk_O:UGQ
m`N1ZelBY389da2<gF@;KjTdlY@n;KV6GZm:kL0jX]OaAo4nJ`2qL;]]g`=I>FY7
K45TH1Z5?6i?12U_e]gXK8_kH[]Tg6n7NbBX\@8F5OO5QM?XU>TNJBT_i3e_@0Se
:6<cg4bUAXV>[\q^R^eE7H<AR5f?TJlCD:Z>_=dMEaZ4M4J>:39a03=KgQ]HYX?H
A>ARTCZ>FhU4Diqc;SoB`4AGAQ\G<jL>nEQ_G>EeDUkb4OXK8_?j7A4;2UGBM5cT
gdTX2QLBnd`WK;efmdMaHTNT\11m;@Cj=`6[EgIc7UfS\b5E^2@bYDJ1[Ud7I7TI
lQg395BFU;Kq62S@m8L\m<0n:^P0[T=@`ODQlmB;?jbQOFfc6SgI3kA?488VXDSg
D=EaThi_oI2C?=gNOF1`J8hL9FXK<ibNF?a6n;IGWeK9;6G<9R9lPmfLOH\M5Q80
I8Y8\oA6p@bLJ0TB?0:HIkH7ZdBl7dZFik5DYeA`OUTh^d^^;<<1FkaDbBHU2HO>
M9k`b4WeZGEYZA_agcWBS1bH:cAWPDWcBhEciBP9q\GM^bVp@7B<Yj_$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FA2(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;

//Function Block
`protected
nmAM1SQV5DT^<NKhmdd78l9JRAhJED84_QJHIdP5JfZqS:_\dKdh_bIb>gTcB]7S
>LRS:gW\[gk0:UmaomagR@CJX8kRo]:_nmg2MX6jg^Ipi8KCY;IY0MN^=MTC@PX:
Sc@kfCCN0K5FlBDk=2gZk4Za3?qm0f>>bqc4T1Kbph4R0LmL[AT=gZn5\2OZ2lXE
1J6>Hp@ZYYGXqN]]KFC_3[Y@\<;MNhB126nWb7K]^oP[qdL4I2]WEnZPI:l0Z;Xb
m^@HOjd^SBmN8p\@@Z0RjF_OgN1e<5^2`g4?Dfj8?ZU0ohcDq4ZOMn`Qm22WD02F
N5g0\QBcmLHGM_o5Gk8WDpa\D3j9HeJoj7;^[L;7]ZOjVE]8iKefXF6QaAdBo[UP
DRXCpjL9RVTO\?D9X2`cMEo9ciehiHRfe^@a\7:9:q??\aGn0qO`g4RcqGa4gTY^
Z_meH\6JASUS99_1dDQdcZ10g?jXMWfkKg@SnDjN;0oGi>U]=cR5e;cEaPa57@BP
k0=jZiGCZd]hKJNh8UCLZV]4hDXIHi3]]8NA1BFLXC1oj^kM>Ylgp1o`BlY6mGMf
Tb;]>\UA04`A8eHoS24>3N6=\L3AM;[4edIR1L0A^6Kl_dBbhWKDj0PgTB<7?ac`
iK8\UJ@<o;NEVD?Td7?2C45Y@nDm4hWi]PF[5djFS3eeNNQIpPkc>2JGj^\NnEE5
OG]O4@BYMMG1ifl0BilSJnCHKETR<R7LIo`2T1XCP]H6io_\RAkNah5o_?Zca@_P
J5=j?5D[k:P:DLAKi`hOWdmMC0mQPEGcncVk;dglT@I7pEKQKi[U7UC11Um`EePl
FLfkk6b1f`55lR<efjab^5o[7d=jL:Cg@j^8;TiI6AIfo@dUZd59o35]eZJiWNje
`AeUdj0`k6SV7DdmM4>e6o]A09AWm\GT3ENF:5cOq160lQliiCOQa`i;S<830aN?
Jp1JfZOR6Jn:Jj7]UZ6ck^ECSOI7fIWHnE<HabDEgd1_;mSbONPFjCHjcmAC;7TL
R5f_Tm^6aj4gnBg9LEEmI`RH8Q\H3SqG5cc:ScT?AYIBoP`5OnOcU643UUK`3^6O
0X0[OH^dGboB3f\_KHfOWK^497B8dkemGQiV^?:oe:BYfiL?5OcVX=^lU6QSX_mU
UNDLE=e>kbSZ52aWmf>9kjLlai;pFNNSaBKhZRI=i>jZ?daBTUIa:T8;6Pe=_Pob
?AXHWbM4mffK1IbdL8;mf_V7O[4UmmiFO:MRA@3ABN6\hYEW0gJ34T^;6?_O4T`Q
HdnWJWa_BOK^aB_68hi6S[9hqFMO`0R]W]B48PfnTaVTXOW>A61?f_?Kd5>jJZ]i
6mjS9n9EPZ;3L_k07Qe<NO8Zd5=7IfZ<8`g^`0P4TGH^oNLm4A7E?OSpVLFBP9Be
9\edheLfNe\3800PjhZS1abGooVjb6ml:H5RMF5WZbghA@B11J^aRccM=<U[`MHk
kiW2d3JG?3]U1M?B@L3@>nd;7?G6dZ7XR@:i^Qd]P`i`l0J3_c1p_@L3J4:K5^ES
7aKO:JQ^M<F6KV7A^STJWcNg_Vl]`BmaTFb9EKU`5[2AGF3KAe_gjQ0PPG[@g2`m
0ll0^;fa^:77<T5[b:dJVa`V`A^@6MSl]nL:WUQ8@;1cc9Iq^Q^`RV9ZZbniTIRb
C:DLR\G@H2NJjoJm4b;hA77Qe?KG9TioO4flPZen1aYd0GB8iDhK>NnVq>JI0a;F
bfQ2U@>3Ck?Z=[GB@J[j8Y66HmeMWS:hYW1m?:Iloo\HNl=89kaS@<Y7CiPZZ_kR
\AoHLXX1Hfi\WXQ?IVc66EU>Y85RD6JVXC:\SkNc5_:Dg=5c;SIgpV]Eo8F7B>[A
X<:@Vmocg5W5kDGLa`mQ8MGKX=?=95\O13[nkcPa`jQ:T4RRSmS9YS;@4=3T2Uj7
U4Vc7PC\aLb86Ak;V0QPD2_ANS90ONP1A^XfhkijT6cm3U:FpWQTQK>j_I7W`1VC
Q_;bX[9biV=__Rf6hGI87imC7_F2;:<gVUH9o1>Z7lT41B`EW2onC_KBN6oFIFXN
=[P>gM2WbKC`Eq8m9`15i@;d>TD7S_2Ak_T=Zn37`U[10c`MA6mDZb^n<W`N87J3
fml<fe3S=9@l6]@KFVo5FKh_gLo\2X4^OoSgiBkaTF:DcBXbU@T;THFjNGb24m_Z
@MTRn2pfF?kh@i9Pc7OEa[VF;4\Rmingl2CW4XmdUcCPg6_M<E8Mn?WlV`d;MJU8
C8=N?kILKHCZgef?5YM=[:i0IH:>D1Wel2C;CI5nT8UNK3RIdenI0EJD<BWL>6D3
`4gp0X?LA7ii[ndG^N?gA5]7ZDh^7Vl?ek25MH<J`Oa7OGHVZ`n8fEB2L\FjT5Wc
lK0OS<UhoX?U6kB[E:blX2cfo>eBmJEm32q:f@d=d]\R`WXf3jiaRe0B[0S2CP86
G3]R8HT\JJ^@6h:M1`iXkA8jT3CKgV91d;8:g:knAlC66d\Y2XO>g>DB;iEc2^ZA
]3^geDmX]VJ<70JTl@FLWjp\5@ImDJO0MW`GlWT4d[7[a3:^BJ809bliAh4Qm9WQ
c9OoZhokXc`CjO:1S;OeDg9\kDc_?]L9OUMZ:3Ic6fd0DjlTQdA15bgeao6>I:>M
\5XKhE55VjpKTj<RV>dnPGHYj1;]bj]Mf<M^PWIX\a@n?_SOlU`Rjd1MI^U\K5ge
LSNW8W2kU:SKd4FGOc]TCG>?YHJjm1d0[@[@]82PRaTXWaBH8IUEZo20GkTkc=p?
iCf<FOKURaA4@dPTg`@f>Od29kOqX5cTDJP6@K41S>9Q4ccGN_]TQmJYX3loi0ke
<CeGPK8Mo1]n<BJQJGYc[eihVPXIX4253h5[jgNf6@UjCC?bN;>V?LI_FIl;ih?1
C0QSZgW^FOY:gRXp=NNd<<h47EEf_@0E03@JEJ3;:0kYLAkHTe=jn6QKP1W6l8][
Q:P:RIQ>1e_VT07n=R`ZJnIZbEg3P:hj9;;ZlhqDZ=YgfniZRj<Q_[n?c[24mkS8
lF9`PI^DRb4ae;G`MYG374DPNNjeIJeR4^Y2V[WDCkg2EafQQhg<@2a[9ncD8L^U
:6h8`JUmRQ4fGe[D5[VaM>4a3K8pbkc_cCeF0Th3e=aA5D4^]R64?MFhLL0hB]>D
<RU]g`Dom2>80PD\G]CHOQaEX:m5b62P?385A3a_bSCIgfi`H2H>Zg]TZae0Q]TB
bJIf2f7Q3]BJM2JXqXHF0\VMJ0giZYi5kDG3hBm4]Ha:^>SgjA`Fl00iN5f^;T?m
P>SCD\4i^FWYO^k^CXB9lFQ68j[O>9>9>JC6k=\IqK?1@KQq@437F6=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FA2P(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;

//Function Block
`protected
ofU><SQ:5DT^<c[i8SBY8h1_R8U>km0UT0OX?lT6lJo^:4X=We<f4\;=q;lak57b
WJA1cImKDR=gQoToO<GECImHk`bCq7SVYbA3m1>n;nW;d5\7oKRmK=k^oD``<W\8
27L:Qa>NUbBl=`7a9A;kpXILLn>pOO0b\MqYnj<:Ig_SZ53[onUTD@X:aHELFAYp
XIR=IOp4C\h6bFE;gS_afKf@QkITVVoVR]L444VdRnqOZSo5QQTZUQ>VkDQ06ehA
<aU>5;l9BXqR^UBmkNT1F=b?P6AB46SihkL=^4JLPB4qdLXMhM3A3>56AME2KTMQ
nE]1^jRMl@0>=Jq4l^I[f2<OWeKCl3VggcW:@04Z?BQI^f;BKbhq^;JLZ4>6Fdb8
Y==SXT4H`YVoY=HFjR44[GM<pjG>^63?I;]gXXEf\TQ8\RDOkT;AF1AClkI;]`H5
bYl^f5Y9HVNTm0eR[Vno=ihKY1kqVLah<YGq8OF_cTqV2RZg`<DaG=eh1UhiPIk`
F8LZXOBhcmdb<5^<BJfE=8fYki[`QoGlJWLk\m2Sc:AYTEX3<n=e5AG<o[<W[ZZT
^foXh19UW=H85^cn11EiURS?S=m^XGgZ_P@leXq4HTifVj[A5S0;Q^LMHJQQK18D
_3MNn:OJbgV]l]n2@MRceUlR7GH;[m<W=4k10465ATC7Th4^?AdQ:LOC92hkPUJ=
a58A0f^V9hh56JOi`CnJ4kTToTTa<HJE;7p7bK7DRZ`FgOl`X`C7T<1LK><ZZ4k_
]21g<<dHQ79WZ\R`084e_c47ha<1F]ZGWiLcm@MhBWNHehcLk_YN4=_J2G0dXiP4
6T?_jBBHbK\LXZnTP?a^^aeN^4fO_5pAQi92`8HhACn=UP5bHB[iMWU?2m<3JdIg
OCdj^jeFTO<[bjI=1BE[]9??WlNS9Xfe>@\IgnB7A>>KQ[^UNm;GWXM0;XL7iMNa
LN>9Ab`dG>WZO7Mi<<NddHUFL`qn=oKC40AU<T^3^onV\GZIfXj=`Z@2GiKFn=5j
UBI9;_LAn9ImDk00c6b^`kE9_K0_JZ;l@a=1X9;>NRK>PfTjm65KKNnq3Yakj9Vd
k:BTVU0b0=d?UU4698h<`;hZAd[HemV5<H2gkS_Xo;Z:=X8J2UefHQBm`2:9MCcQ
g5i53lNElBka:h35J83c3>M;7X287bgc7:0\:d3MjGjce6PdT9ejpDOHMgKX7oIR
6L2FdPokFeK?h9LZ;PBk2ZZQb@3J<@XK8TjQT_R2:>;i6VK\L2IeAdMVL[443D]R
7[nn1CK]j<h[55LT;[i_>`kbScN^SFUl[k=;mbKeS\7HkYbLAqf<W?PVP2oYkYB@
\ILP?m]QZJCg2eB]\VJn3R1NhM=[feGONYWK;e9aDbQ;AqWQTQK4j[IPQl1VCQe;
bXQdbLV=g0Rf]^nI87im>5?F2<@<gVU37V1>a7lT419]En2AnC_KBN6on?ZXjXL8
1AWKf]7Zjc26pcW>:R0Oi^0h50X2aoTF]gdA<@5?6hkDI[cKAVbPQfHD96lBn1Wk
=O<\h8YEUc5R;mCB0gOY:`7fmbY2E11P?FIYcTTY8]<4XO8;[Dc=V0CjBY;VJn1;
LW?@^f`Aq@j8clG<Vo\KR0<FF6hmgjYK=\=nd@DPSglh2K6G]HTnC43NAB;U^ki@
6HbLhm;SR@HESmDhD>AoRSJL]DK0:Dl^71[BY4jb6TcC=EWd?TQZRJaflF5m>V:\
]2Soqkd>EJI9IoefY9J7AHEjVFaAkR8RILI=m04bKAL]N=DlihK=YTohS[8lJNWQ
\NYnAE`l2`^;=0geKe5A39@TM2;P35JLZCTfScTO3h2ld7P<f71ImP5OMfX8L<ab
qlB_f\dT;d5XZn^`flikJLmkNRM^Occ?gXMmbC0f7i@3YMXA9gWi0j5HW:]l8a79
]a^nNi2LZ>lo<^LG=d606=lLVeb9=1om4=lnjV?4eXm=>4h9>j5k\06m0MG3q2Kk
di8O:BG`D>o5iSigRHXOojGA_H]@\Vj;\`n8]U92I7fZbAVeldQTig@=oVQLa2CV
^e`VfX79gmT:@;lCPnWT=<EcVq[m1F75@ogF:5LXFYK5HS44:265<G:hESbO[h]A
@80hnCVFIQMma[`3INE`qElo0LlJEb`<KU6=7S?MV7RRb5J5Tn;_5;1\0Km8XbL3
]4mAMGN>Uf:Vdl2_nc68[WPeZG5cgaNfPKJSiNO[_?3W\mJ52`4ASYLhanFBNA83
NKD=[GG]dRnjh>f?jp3Vh`86;QEX\?k:bTGKWlAd@JK`Ed>`<XVP89>Ejfjh3009
C7`LXRVA:H6L:>ZIXO;I:ZcD=o=Z^a7`D=_LUgJncjY`6]NoFjNHXTVOf=bM30S3
9`?]\KOl7HkASZp@8RJI`c4a^iOZgl2EXZN1C:Y?WS8oefkH?ST8R??B4`J:hIZH
IXbnnC]IW\PDoDg4^knA9F0FHTiJN994nFR26@oI167_KpR3UKHR8>iA73Ed\HMT
bRAI=h^@K;Wh3TOI`APf[f?KKaDJ]5kaJXGW>a8UWM[aZ9RWMVF?>D0eQV]J^i^S
6GJS[W]:<a?K3nNgL\WR:7Jk2b2@FBYR>qX=XPmEoa2M^efmk343B`U0EjM<B0M>
Zd5GDIBlaQKXdXORQNGF@0Gc1X=l:g<ob0X0NiDZV`c:em3cbfom]3bc?>UFS[og
Z3lZLPPnn9UZkLc2<R;`jpc8>6dikVIQCKif7gaZWR1gA4elY1=C:jkPS7bfoVCH
Y8gngL9lbJ3LZgc0f75?U5]Fd=j_oQ5\Qj9c3bnH5UA0W6M29a2\Rnmb?93:UYb\
9F<H7HI;W^Fb]pC0C;SQ0^1J;gHBQSKR5mb1DHMCTdeK[TBSfX\:Bbpo6=m?41h5
6fj6kJ0fo1LKcWFEN2=Ma?4K9VGJ2m<RoFiRYYL2DlKRKh=d=ND[D8Kg6CQK_ljh
M04`@Jl9ADBLQHZhLId]goh6V6KWb=@S9Q4O2[Ba<XVJhip4Q^HD>[8U>S0ZcegC
egFQd<a:ag:XX4iB1SOaZ5VmgZEmV4aGQ37dHo671iA<ac_]6eo=]X2?PO]n2NF6
`5GIG<O@bp]E_m;42_T8lh434f`>VTJFcWEL>CCJNGQ[7^VP^<hk<FCcXd[DXjAE
01?l_9YA4O]:84@e?Ua\HH:0_\bRIVAalecX6dY6cFX[7B`4SkUgKN13dS`UQ<ql
J?O=F<cY4nJZdb?g4o^FT6i9NP7bhHVpmA@PW9@D6K:in]@VPfT_c6?e;nO1o]2]
8VB@H1@9=^lQV3=3\:3Ld5<VIYIoUES<mI<NbJOi]@agLQf2]R@MdC:S@m]3AJ63
7VBW<4@fMX_6[G5:D_anqJ8SWLBk0;GjTNS^ZhNF[2HX[8MVZ:D=RNm@4j?<BQg1
OAA6fkDDVjQK:hFXKPlR2JAIhD1>i5@e=fYSLBHDQj[UpeO39U7pPKjVR^c$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FA2S(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;

//Function Block
`protected
V]d`nSQ:5DT^<L0YKY<aOgo?n0h5nGGTj=XX09TcT<A=MTEbZVo5lPm1b<J]0<En
^a?^_AqE6@^fKGaMBHfSFZdc0qQ>2Si=oDbG[M5Pn?H10QC5;^WSXRP`@i]LE=cJ
;^PPFH8JJOG5^egZf;^MhY68UcTWq63kHbDpgF<;Fbp9VH:hJ?N1X]]`7@;FBNY5
TU]Ngd1pC7lf4YYKeJ@Tda_jWQYVq=GGL\1pnMb<OB7hd3^l6afhC<Y<9]DeNn8N
G=5pcZ[A`<jW0J:Nfga:HWY^mmPhYgh;Q578pYfH9lYX<l1lok87@ARL038`5BFF
=\;H7PJpX`[9SU7;j>Tj07]HI2`PcIV\H_BmTWeS]^2\q_T\;i_DJ7daVH0f6o1P
][ZCFMBWjad<J[?_:qbYOBd\Tq32NN6V=DM]aZ><NZ\VA>QbM:57K3m^6Oj=1Mnd
Vjgl:pamPC>CqC>N_SR^h=8i[YomU^c\CX3E^@_NSQoKD_\mCO_^;66l6A:MkCWm
8Z350Q3ljf>SOQ];lg6@=dJgiXB<k[gFY>IIOA3]Cn=\AR8<]1hYk6UP`^5_1R7S
LCNe8Nj^pbZ_A12JQ0JfO_DWAjCD>H4KeJAAFCYSJSLj\nG^:\V?PPCmHM:E475[
jJ8af[HaCAPOJc8D4o>C\?Tol_2a\b7m9Zao`87AXLEJ=JhnWb=P>?]BeQ3;`T9c
>KV`pg?>ZO_?W^RDAAh_ZUaULiVRFUAWRalU`iGj5HNH@VOd?3bYb6S;kLn_cS_U
4U7EZU\`^PI]]3<n0G01`lOe\i@DfdEe[Fc5N:cA12lk:B3h`n]\k4@i94bCbVNH
p<_PJFB\W;<^Wg0@dhm8<VPmp8gZ`fWGjciK5fOiAFd`Z6Dg:WGPRC^`B<]?LBRc
X;52:K>;_98[hOC_3=@WJb<A3gjEL1hD2g\<bdX;j4]A:J<I[hoD2XRMmSE_1]ce
8GSfC[1Hl5n3O5hRXJ@9pWVgQ4220Rj7G9PDRl\Ak6^WCnRMk[eZ7XmD\8S^;4:Y
6gPGj_flKO`lGO9]2@CVAn?CWc0=;I@_L3]fDG@DnSmU0MN@Dp?e`Qe^MA<ZWa>h
knISYiPXBbkaUGWTSiQQk49UTnK77m^ZaHG0o`]hQP>;;BcnmM`aFdLEle:O<2Zj
ljT5]bHjYF8abkP3b\1W;KhV7?Ge8ARPeeDkaEEME@1iQjqnmaWN1_VWOFIfgE1N
?od335U0_6R@PmSb=\Loj9>bd\XVn9EWM400]mi98<o?:Y@CdJ[P\RDFk?B5?T24
^UN6Ce\W_4^O:9;@R6^dR7?QZdn^FlDB@?Rg4fTJ0;lp042IE\e4mn1?3RJ5@1[n
Z``InUXO9o<TBV;8]k]h9B1MhdYB3=@0_oXhmo?1c>Pf3]6]3X:>5_<bfc0S_O`T
DXkZVALhMiphQPIG8nZX[7XnXVm>@_JNhb\2o:nIiSFRA`\G]A4H;Mqc77NAVge3
U2kS9H9YLNYS[KY;]@YmAR0mAALbI@=1J2Ob0H]3D`c[j8[IRkhDBnG2@WNC^[BA
7QdCB==<9J>jCCkPP\n77SMHYNXa?8;V0]39b]jo]fL]8M6T0ap=fH1\_BFa?RZJ
4GeTkm:NG9>KjfS94:@U;1>0[RGh6MHme3[>=kh@:0TOF66NJ8I`1gW`mUBUl[k@
>d]no`BWken]SY0fhTMD4P:8gCaM8A`jQMTA?hRHVWE:Kaq3cdP@[4^iV?3I>bgV
FdS4?PMl[gKN=Y[?JbZ6L7^k4Qj<P@mjMC3iNjdQ]JS\9YPQDZSKIGT7HU3QVO^2
T]N9RU[PTLkk::LgQc8oG6PdV?B3IX3bfK@OK:Rgj=pVUbLTaK>JE0UC_iI413nX
e6fmkYPDFUZ2MNZ@PH<XakBI619OUQWjG]P<GA[RX9L;<OQ`TE7cS_Y=k:UkXgWI
a<CW<B5:h8`dVX1g=hCZ]P`LObQ:a9X9k^FAQLqaWCOU:6QlBB1MBAEA8R6?OE^9
Z3JUD1>^:bNS:`<27h3i;<Y8F5joojk[bSF3:Wi`I9`]aPWUJQ1e8;=@=J9bS>RN
]]Zp5G4N<mn1g9FZ111Sk_P6A^4Lkc:CAm4iBUQMm8`VRl<IDXB@7^ekekIdiAKM
[;lolhC[TT0Nd8gfd[e5KEi_2DV`@BkjHAO:2G<eVT3eYBTU77ncHkFG13]_pNS=
RU4eUX@HSJ>R57M;e`ZTcV1HFmP0D8>[fiE9CSZMeWaj0T3oB^jTN=MM`[OF`cg[
l=AXcVH`UIQ:WfW_T8XYAD1NW3K5NUCHEEM`MICS05R6i9:ZoK7KkE4@5pMC=mDm
073[]HL>VU:f>:OeKbVhA^J_3HnCooNW7BSj>bfJBh3o9V3O^@S9YO9E3cS_e`LS
L_H`I_\XLT29E<^cmWKOTZ]=qHffe=k9fYNE7^kB@;8GOghffdV?;QaO93jH:=bD
S5HEPJWhfDM@<MMZhkBHGkk1SHWDOE3h2>=XafZ59Bekl^B7SbldSV;OPT0854HJ
M6Vn>g::OWfBq0j?7@3]DmXfEUlplo]WQHkB1Tck=?BmHUifFI6OS^IPW9JLBo>g
:U>MR_2K7I9BOC28D^TNISl5Xi?=lD;=f;QMLjj7GB0LLhjm55E9PS<mX`JP;fAl
OJh2BM33T=3Z6iHq;e>oM=2L6><Rk_4U_LOTam6OXO=\YL`cWb=2^SN>IL@GJ4BJ
JJ8\Y2G]9eOaL9?P;S?omJ]>]]dSZb7ejZ7S287`;]\ho6`XH3d38DGiak>[No=5
WLmp6<igmj5@=;Cm^`7862ZAD_N<GmkW?3i\m8cAbP[n[F3hHToOdUheMgR8HCUb
BhDe68JCKmE_2QAFTK<A`eDMkHNLiB\^`GimgNU`BN^8@L8?XJHJBkZp5QO`0VPZ
L5NR5O@54d]iiMAPIkB\DmWn4Vhk:eSi1aJ3\>E;8_e0aAH6Z^SGgaVe5nC@_Ca1
`:6Xf`aW`j@]BPpiQ9Fo^g]VifJPSXDQTgcjiQEi5A43P?ZkkU8D0b@Caca78nmf
`M2jUGmVcI>Y^k`i6GI[OLbX2RdK3jBA_n6Zolno7ZnYcNLTkJ`\9YLLVa:2Y9mI
mL@pENo5T[ZW=X]:B7U83L@5HbLhNVSRRGiRab=I0nBA0<FFg9m[;2<F1<lbjLUN
4^a9EZ^Yd_n;=fGG_5m[VEXk?oN@kf^TKL=0;bNh4<IOJ2oP99\8cMfMqhP1Qco_
N`6M`2eUUb_GZP0SpTo1OB6KG6bdcV2m4;Y:?^@8;YAP[M[BNZ_S2Q:J]o:\2<PT
;Eda@l9KB[TJaY2[:TBdFRGC7XF81m8da1kTek37qfljd`Wqb>?dQ_V$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FA3(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;

//Function Block
`protected
N8TaRSQd5DT^<WmHL^OdYVSDpb<YBaRB\mRMbZIh0q3?Aob]<Hkinj`6CWnmJS^I
JTiiHj=L1eHdZRn^Uq9YRo`WpSZnm]WpJW;55lElQZl;_R1OBhR;G33JL<0dC03p
^1SaU9HL>0Ra6k99R@omYHX;8XD<cY6Pqj:1oLi5DAOi_e=CTNbAgaVS\mgPPChh
=pe_6C7>\>Sn9ZPllN\hdeg@OB[j0iYDm6W>GqMR?EEVc_QdK9TWMYik]5HS37_h
GD]51JkZeBQ6pPhkeL?p^<^EFoF<9]a1=UG:PDLZfkO6MT@Qq\k_cRIm54J5Ko<4
^IXB4DRWLLJc@7=qf`7H3JBq4;]6k3qe?TUf7=d7<T33JA\FY=CEN@6RBY4:47nQ
OJ=o_T6;cgNmDa3B4M>Ihb4Wm[SHIWh7Mbn9OLPX[`T5Mi1U8Q>11@l5h?<Mk_Ja
jeLH>IXHEl9_JVST3DP3;\J=\=pi\B\BT=VMkoW_k;2AEiETTG;K]opB_<>TZo:<
FSHn2e=E?9kISZc1lUgS30>Mm1^On8:_Q7noR[]\2;^:R7QAJJ\fZJC0DeXKK9Kc
IkH?WRVJP13IEcb5V:OC6bTYPbe3>MZn3iZP_OXhSi4fF=TL=[pMPW\CmZ:F:n]Z
=dFdM5C6R0@9UaAnDSdYdb1?3_A\8LVdloGOE95i7Q^ODJHfYAQ\`<]2GJVO;]S^
LC[=IKTA4<fEE3\@AJ2S`7IhDd:iKZFlBWENU@``[m75a?pJ1RS3O\3=foE3R;0P
S@VaVo]9E:5;:=Cg52JRaQBE>m?jODgCb3XA]Kh3=Sk;>Q^5\FWLnASTU`QFAWD<
N?c8onGD[:4ESO3dDQ@I@iJnH\EiIT;\0EbnN<;^V1qn]G8YDkOPLQjWEKH`BQc?
Vc?cmdkql\07kOCh68kOc8KMjU83>Fg75>O>HTA7FAmD6Q9DJIOl8nhU\A2VCg:h
nnb9mU1@m<O>cggH`_CGeMI_DiGogcE\c>n5qM88jB5P]f]a0o9Y_7ggl>5XE7o9
>ho4<g?ddUhJbejSl[`Hj=K>HhkC`S9neKkIY02KIO4Jmh?aj]=8ihjlI>H=6bo9
>Q3Qhj87k5:VBNK02UFBIQ6[8HV`I1j[=qMOSa3hWY[_4:5[mDA2n7774BO0XmfR
i=c^X0<Lm2KdFhIQ^M\C0fE]?V?YmbGT@>\^6Y@7E58_E`6m9HPAkXe6Z1K0Amib
mXefhgW5aNCb<h]=04adIX[kkRXL3fqf6d1Kmf@L4ENC3Z2WgZneac2O344f9856
\0^cQoHKH75P;`G:2eJ@gLF<C803UgXV37UgG8]BfUG;`Gk_D>X[aMfoaP6lJqSL
HPc0RHH[3FQ@QoCY5LhDl=P=ZUK9EOeU^8YA^pn6iG6>3[`h<SlYT5Ra_Llhck_@
VM\=LMPj=>FjiiPVITRmA<cIhl<l5kI_]EdIY=Z?><6@2D1N0@[NN?>aW?VmU`JM
Ald>X8`:m08dE@YDUF\>\8nN1J9XdI6f9p7n40J=AHV9<RPNGY<Wb8Vdi_V8gARZ
aFK>lUmjOS8^IMDIXJm>:lEfQ2K1NjnWHgFMCn\P@gNSHAI4U6QUh4AXPM0NEWC=
V_V>XCQbdIdcoNR@AkBeCWHMZMYnip_WigAJ4T=FfT=6\Pc>Ma[1h::m^7ToLN=;
IVg`Z2De]I`[C^TKXa=iliHEMA6:1e1KaojK`bB6=^598]n9=l?NO_?9[OW;lmAf
`5F1To;O^C\l;i^J;c<:cQV_ZqmIeUJdHEg0RT92]mW?m\ni=A[dGFMG6hKQeeim
Zf5S=MWc^?=N]=mIg^QN38FN5`\K[M2Pf`DWo0Bm>nVgH4n4ShTUFHTT`^Zh8Zk@
9]@jonYKYYh;O6oldcB^hq6^7gXNFYS2b>fjGDd@hno5:>N;8P<AGJhJRn1GRo]_
5H5X0VA0WA^<>I`9^cVC_N^QXSHJB7YZ\Noh@]^:D<\\jOLXUUqo:A<1@Q[[J\N4
Zh>T`Q@gQPT6F;W2>:M4RfhV3fWa=_@J2c;R62nL]:h5c\?EEd:48W2Pflaf8IYC
@bf9N6Fh0`g0FNTJHfBg7hL6G_eDB?6I@Rb\oP3GM>T_nUap^3j;eT?<m9b=nAc8
2VM]?[R2@hM7\A7dFlPi^T<h_L\<NmhJ:YR>6SVTmGH3@KX;TRJ9cVEUCaK0h\nT
@b?11SgV?h_^R9gG[XILBlon;GGPEnd8S93NdQPhe@bhq^5n^7UaVg:L_2OkDcOF
J0hi<HlcX;MnQfDMg4N;@1dLN<3`ml=oILi5Ii\5W?@;SBmRfKG^ZLUhQ<HS>>7S
mEoE^4I`oV[qDXaHoHEgRm2;XK4q2hUh:3^RG=OZGnmk@Q\R:NNO7hJ3`YX_RC1Z
oZUa:KJN?II]6UMAK^klG:O]3b7G2Pk0DekSJLF5WVf]c>ZJMd=O\_JPakX2@jCo
ZCiWRWCbG`S;Gb0q6:dJ?PV3jiOB15NHN`CMZPkN3\nM8\jlAj;IL:E]jSWfiD0W
^KEX8mdWGQeGg[YE642dNX`?00c;2``V>1<bJX<R9iW`CRjlo49c8lTWR1:B;?jk
9[Wq3;6ReE3iR]aB4HJ=K_bc>04a>DPWPTE3^X1BAFeVenM<mWM`8SRd@hdY>efb
\Y9k3@F2ibY:D5WUaUOkZS\OnV`n>`K:9XE2KEC\mEjW_bRiD=oij[hqWD?=X?Vj
MK[7Wo0kUGek4^f4EiBdReL<=gmI_2bXOe>F0D_b`3gCL_4MA5CmP\K9WUMYTnl5
g_SkFc7f>IH18[NQV^KCliLL?MA\M]a6PRNJ>eZ_ea:pkN2]ZLW0YoIZGMPLX>?3
hZD?UF9mLB0`Z=M]n7T<e<0>=V;RV8_BbK[TTS52OS4Lkif[`\7T]3N?30Vd4\m7
l;qXeXk7e2QY7>aN?Va:\KJYM4:dUK_?9BJLK?5N0KV`n8TU=7M[B:];[94oUkKB
S:9X[6oX7;V4bFJSkKm7Dj]`b]\edgkG<NQLK5I0:b=a[h>J7__Z]<TpaoC?6BKG
AJ6P;mn4hXgB>ciBYWK\_n8>SoA3>a5e1XJKNkkTgUB74LQeoiL?7iooaCONDjh1
823@8C\83mJC9@kA^UBbE`?6^oANM1e9d>=^en\?;dO<q_>:HTX[h4A1XGYf=dbl
=K6l12JiBJg[j_2XQ4<[o]b`HXV8:Sm6oVk_Bf0::DT2pTW74k;`ISnM`]B;KReB
n2EK32O^6<]N1BYG4Q^QT]RN@D;:E]iU;JAQ\H4kBijBNTWEK;WidO]ElkK8JE?W
Q4SDq^4i`D2qPJ^S3NW$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FA3P(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;

//Function Block
`protected
NK8\NSQ:5DT^<^;`JoLUokX>SViS8VjL3FM]VPpRil8Tfl<R5Ec[SYRdDlH6m]??
lP:pjGQ9O7[lJZCA8KPYF^Xhg<9A]\;1]C3cX?VC_`N@8lEnRV23?7daN565>EnE
6TSq12^EHmqA^1^bDqC0@^OWNTbnV9eMX93dB`8_^=P?;9Z[\pg?aJkN1SZ8[nDO
k55CXOZ]eYb^2DLj\cpnZP3VKQfY7RLaL@Z]adhjlHa]SRDEll3p]=Q??WnNQDNR
3=fLf99B9oBkJ6G<>7^jJ:^q[YPQXQ_Y7S07cC7:K^:ED0on4c9\j25=\M085:qQ
CU9LYJf441?<7:]GhQ[h1aOm2W^38PnM=<WVF;9p0c4Xh7pLb_JX3F7aOnKN?13Q
LoTiGb\liYPpL85A5Z>qH\N;G6qY@[oWAPHoknEd0ESNU0:T`;31V9A^1d;41Goh
Lfdf_C02UARbnC^5g1Ni2_nVAi`INLR\k=SiC^gNh7fIVR<DBc2fSV0@9mk^L7X5
hPPQNBLC6Wec]b32ShDo28plPOX0E]m3ZH8`6LRI`ob:INoii]48Z;HGR<g<nZl]
bl2a`P[7a[fDZc\P==M58[V=[TeojCDf1goaL3C\XMfU=B7Zg]U<Tkghc8m=l\S2
_VeKc70H<FLh30H_8]pRWRDTH\eOH0iJgJHFi@j5[?Z0PTI?jLeT8AbL`J9J;bAe
IjKXg]dG:@I3gIMnVe?B?EF@@J]J6V4cZVHWNoE63NY5\L5Vn>CnU^kOa9Gf1cJ?
MkE:o^iSWMc7c5qUb3bmGiEkEJ5mcOpZj?Fod=[mG<EhPnI6la4Oj_RSEcgL95mB
X8o1h9NEgLc04ZlVIR:Rk8Al>n@L[DHlO_4j=X:SAmQ8S6gG0B=Q7dCnH@kRn6LV
Y2fW9>bNLiJ97U7RaOOL\d2k>1qSjgo[nLc1dGg:kTgWoSH0YV^R3PB?^F8[F7a6
EB]_JhN_dW<6XCkV1IZ=hkD\ZSKBLQk][U6F6l\oNOLA4E[aR4Rdk[Pp9j@7DF>1
F9cOhFAk27SknkSZ6JEN_:ZkF8Fg[27biRdZ_Ekc3A=ZK<@^L:VFV6f<KcaVM1HT
NO4Rh@AJDl`U56KNDJEN7jh_I3cWJc1oiBYL5Rll=@X<bbm;K:onp6V?;i47TSI4
oLhfiPD=Pk>9EZgT:d\4<bCG]6cLIg\Gb_C[Mo4]Idc]`1?9f2Y:>@TdfjhfjKaU
M[70idHhI;8>_5gB8d?i`l@cEB]Vj`e1PEm]lD]bE?P1N\_\mpCcb^e@23EFU>;R
\bdQ3\4`8fAhPVIV6Z;]YlMK37S]34alaUe?gY06BEP:3VBC\IiianMXAEm^mWQ:
XY7jCS\5E<kZJi9ApmEoFMD70ZoL:=2jMFFJd5ETIqfR5T^Cham3g]El2B^<Dk^8
G:@8E8La1H@VWhn\HJo]=DDd8B=MPN9QFEBUJScOQ8NhdOP7HJ]o<j[imN6K1FgA
6m=]Akjbh@;d@[F7n[=Vk3;Y]ob0I;aBYCB_Uq6jb]:>\:<XACc6em9hDC4Z;`?d
jCfO;f?mdD3MVPki2Qm]R8V@j7eSl2B]=GA6O1LNC8on3SXog]`Om1T==XY>PXPY
DEBQj^Tk`hnN1b;;[>Teh4;Yb<g]O>bY6q:8]jJdHcN8E^I`63CeV_1F`MDLiA\5
?lX_1dUbe=gK`2=>07QaI`^_nWHoXBZeFeAkVi4Df^7E;EJX4QSOZo1Z`jNGJF\]
bWMKP_WGI3QGKif_VIm3dYZPiKQ9TpBN?@CIB7X=1GaLC>RCQC5CPOHE^YDhJ>@9
j:ZF]3S;Gf7J9BJ>SL?k28Y]_f>>Q^\iJaFLiJD5:m>O7M2gH>0Jl^Fhi>bon`WY
O5?0HVhAf=k?<1;2aY3F`L50<pQa]XC[;XKXV9CP\4?N73IfY^@NT1826hH_F`me
m[>99OlQfk<aD?O23nC30m@eh;3lCfKJPHR`C]@?>Jo<NIe8^Zm<PSq`9f7cP:L^
V3[K8bWV`<O25CRki06Q<7Oa:6^218n0_d:A@HHjo`oUKVBW0TfDZf;Mn;c`Gf]l
EnakMk\1fE:]Y082iKf\lB4E<?l3`e[6DUU^1M7Lc`fc3On`19Fq^;4S3GjOLFVd
0FT<8><N_mTM6a8dOG>Xc_WOk09[`c0T=nFXc=3Y8CNeaNC13kF[Tk0l<VMBoUfm
BBfRAEU9lF9]7a7dABc:[Ai7Jj35J\C9a>:<5FaQ`LEXi\BHp\V?3b\ic2ObPBh\
LZ:hgfLVG<00Fg;lgRYM;fALiXhmldG_6UTAfAOK>3JS^TFg2j^4N<Tmi]>`QeoW
6MPD[]l91`YGC0Eqf<cY>C_1fI\l<kX<I;e8X1g6bodQiRj__?9[jgqe?GIBaFkZ
_AMJ3a]T8c`OPKGl;03kV0T;7eO;E^RAd0C]?CK^3?BgKo`1=MM@Rj<6kmSG5AjH
GDNm`d@[HMiR^O?InJDNBJVfe<ZW3ITC1;7`AN_OVCOBg>qP=NLn3`F7o[cL7m80
lYf8]7?]7ofH:FV]KmLcn^^n=\3j`?QDEe0Z;8dFHde^VR5jiKb2jj0S1J:1R?>g
8OLe^5@4onODiK<mZB]JI8B>?jW=WcK02>ejl:pfDe9Zn:JoFnc:SM5\JI5FokRO
E6?XWZHbI3ebnT]KMmS[g94XN=f2V6Z^63BYITWflaVTViH0e[`TVETA[n<RJcdg
G]^OnZVGXT=M_HjUQ3l1b4@VmTqDa1JlKQSj2^HIL;;Bc0Sf^9=gHI\O5^W345GG
<\W<FXhmA^>[KFO:LZT60ck`?3_UmXm@E>X@b[cNA<K5<SR^bob7E?i<2[2YT5Gj
TQaDNeU:;S]?N:R4lNpVdo79d=fehAIek1H5;5NaRclQ@gU`<hGhCS`2Q3X1XaR=
[3:D^mU:k@`AG711D`R[Hg[`c4e81_b1<_GO<9Gbe=43EpQ\SADf11?`[e_8A0`L
h7aW2PG_b67>oYUDk>W;BM7[oOfBN]`P=g^Mdl_nRUZ0Q]QJ[gVe\1?Fb3>N`7l3
h8YMTQ>nk[]jGd_DkNa8?[B:ZlYeS;Nbh]pheTbMY[LBe_f;>qoK@2R`HkL82OGa
O8>6Kmb]:<PI=Q2E7KUI4c:dSV`6_F7fQi=gG2=FGDeH7fjhU:oZT2RR_EGMdV9^
bI8\U_5Z^H:f_7HKc?ZI4k^NCHJdVFm6?RNLfUqch6[]fNml0b8E<JmjDJXX0cMP
oHb:h_iNPC:c52\7YlUiB@V_<QLkjPJfThD[EQdc46Ok77bBHG_79d9lGc>J@iq_
GBe?Rpn@BFSm]$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FA3S(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;

//Function Block
`protected
HHCe<SQH5DT^<<f:07[JDdanS?fmP_0>PPU_T^nLXmB<>YV;d4ipjnMN_M94A6mE
6i[@:QplYc]_DDNZY;^k0^E0=i5M8@CHaY5Y9OP;09eaEkj@@BJYMbP[[n<qUffk
Enp<cBcn4pB?QJ:ABdHO@]HFhRGDmG0=;NR[L>mY4p=f`9RJjC8?h6fl4MQ1L=a[
dgkePpg9]K_4lg^eIPm2BZXmJI9b78Ph=8Ai@1q?J36^>2VKYM^0S5n\6A\QI;QA
aCT6@^jq;]=?MifJ@bSjc@TW]ZSL;jZEc\H7khR9=8?pWgggbO@Wf0Z9mK@:<6OC
c4D=DOK9mBoRIH^Rgap;a[CnnpoPZ_GhVmNjF6^<Aa;GYURif?\oaQqOfZ6Jh8qC
kZBF`qNm<Z_PNPlilTQIeTQflhp_ceh_oa8NbP;mhM`CC<G=fC1>@2D:S\@^Go@a
5YIZa4FRcLm3Bg_EV0=XlNO=b:5W4Z:Oci_Z4D8jM@[dlbQ1NNdViF<=TX<GIPSa
P]HnEo_8TIlkVo^?gAnZLPqHo01eDdS1i]\Mf9L78JQkDJaA1aQUQ=]NDP2[CgH7
SBjE2VWLh8\EM5EL>67NB]Ln_MWIm]aNehk0ljda?0a[=kbSJ17;HPF<[X9J>dJ_
OiG`[<2A7:JcMY0K\hp[5XlgWTI4^45?cEONXl4B?i]bX@FdCk155AS5^INh:n;S
cgdCT0EBl0Le@ooQoUhIiOc83l7D[MRbj]gBfVWmFBH3W50WF2=AF7II6I?i^RYE
el1MgNHlX]80aiq3dnO6m^N5g1cSZ_6QQG];\IeGHelF9X4RON_lUY;@:Y8LOil;
E4KhNQOC9jUmR?8=COPB?XMB?5bd75FLnR5U:na^]F6L@NELUGCcVE0=S;l3BI9H
4hILXK4Qk2p31a85J@=kD<be:jhZB7VK=DQAgcc30Z5;`ZW\8HIMCVlGDoMnc<Uo
m[Y>MLHd6jXf9dUoT\9YHX9l0IKES__Ad`;mo4Jq8eTFX<^4J<CTg10RZ[oO]=^[
=HY[HcG5:m82Dnbf08RHHXE<<Q940Rh04jpO?WTBcOVKEZc[aMZ:l9^g\01k2\\n
5XfLkR15VCi:6WQ=OfVnTC@knK7OJdID>Do@knQg6DEa]SjRQP4XfEJoQW9B22Pn
_BikUCc2=mT=UHT792_k9\:D<5I[NCnqJWEciLJ3E29FgNEd\EdhmN?Th0XC@MAl
1SLY3Hb_YN3_6CEneL:g80CSn<;:F\TRel[AIR=:CA=F^I1WlBlNSd2IL0N_l5ZL
7fGk9hnbRglNOi86`coedM[WdnO`pbZOYFRJkjLbkk_5XROgan8kK2OXJE\Q<A^K
8X6<DWdbjgHREm@@MGF=fgB^foD_a8@S=DhP7XiN6=gcWLKbHXQ_5VKI8EYqZ5m9
^7^UDDWhO:21Li^GSE\9NlPFc:D>fc?YjW;YCgnl\TJE2WcgjAhm65L5>jSJX:JE
>EEfQZBTcLma]]QMjIb;lZcjaHP30glM=HEh7UJnmHjT5iWkHU1K1chq;n9h?mSO
`SM^aohAn?XYWjj>n]e1?O1k[UhX8^G>=GE:SneZbOo?o4XNQ4LSE<Z64LJLk@3L
ofTYW94U@17`C]<<;Q_gePLVgoNC[=8MnZCjO_6CjJ\=NTbRT=DpiP1Ig<Yd0S76
WF`9?Y2bKn?>?LE:jRd2giMOLIoYcofM]]11gi1c?TC_L]FbS4fOZ\8nH]ZXB<h_
52[CQ<jVC1GWLATN;RCjF`0:KaX<Y\b_L>SVVeZgeWW0E<5pAhZoZSm:42QYm_2L
_\JPf;;=L??<BHi7Eb8XVoD_:68m;UL2WS<SV0me<XaKX_`g3lYeYBX45Z:^3GRL
0XaBO<DNHKD6N7\T`HaJ1oRTC8A>81ANfTm]fWNbNHDp3C49TgdJn8WnZYI[5__]
G4@FdS8IMP\L<;H\FmZIm8S_GQJT8;bDaL3QPUS=\JL6TRURRF8]Mb\KlHN=8O8J
T7^<H:g:pVMb2M?e:l;DVD?885M\8Ykh2qnoCDnNSX=NmIO5?nK[2Z_C3?==R2Do
D9G2JW:KQ\KK[OcWZj:W^J[AEd;2Qd_2faCkobOGP@;QMY`c;S1_Y?BYeTB=_g<8
NQUoNhO;_E67\h7Q`Jd<?IM?2>\>6SpDHQJ^Y_PIKmUH<P=ogMnfk`H1[D>2YIB1
970WkH9MfgI@KN;Zc9iO2PhU8IkjK=kFVIB77J^N4b:Og7NMO00X58[;[l@MlZG^
65W2c;PPc7nW?k:571g3df6gXKDpB>K0`AJgmSlRlB4>8FVSBJ8m]U7K>k?_CS[W
m3Qo4T75bj[OECiB_g\FbO7BHRR_[4WD`>7TIlY=FFM1O\R80@3djY3=e>p<Y=SS
]CW2V[NP\`c]O;Ye_=iCd0dEWJK9lUPf[QCK`lgN]0Hd69kAi;DeTf93\H2<Y9^R
iGj0<eK24D_i4miHGnA1]OU_NJIVe5\W16SXlGDc]X4W\Bq88P2_KYVoo?1Oij6T
lLgAnJN63EF_jBBO?RaDANnO?g_hhif@CEZAT_PZUS_k_Uk8A4bfB5`E;e3YYS2g
P^6l_L<fU0`F<BPH]Cjl6X?=XR=?mk1IIPqC>i3aoecQo]`HGGlfVQIS\@:?OPA>
S;;3fnD`c]W>1l6Vnb4U2ChkEWgLGKb78h`Cm=ATf]O;B^@Fll3IcKAAVf[K_D7c
c;iE>BC3^P[<^24^S\<V^4pc9ikSl`oigS]P^G^J]i5lUW?0kd^6X[@U\dcjFOiW
Pg>jU50GFGP0@<hPREb`Ji5cdFYnL;^]cc9]23mj<?ai4Q0eDUg>>[K`2O^eiA<m
C<7X1;WKI=qGc8O_cn8;d4W>HhYmZF_WW4218J^mo82VQ4?;PVgL;Kgh5cO;cVdL
ScGfG]B7`\EG0WUP0``GeV9M2XNIX>XIRp^KMDa<=FO^;7Iamib?@NaMKE[f8\_5
JnYPX1C<]eamKCTQW2e@cl3D]U6b:484FW^nLDIV0@bFN1idKadJ^hL95mT7d6HE
<nWPe:d8^I`1<M]Ej\9b6Jq0CThZH=0369>:470EXP\NSP:i[NEMLlk1`0oZ@CRS
=qH[3KF8O6Ue8Qd_J5KmN`6U03<ahVh1I9ceeX>gNafRjnZm@b\BF]_o49H@l<_S
aHHT?7bQLG\kETYm3Yf9YK>K<HF4a0AF=OneehgJ:nLi;?\gPL34\;qmnaf2obgj
UO13_NE209loM^4@=kP]4TgHe^NL7>J:SCgRR^SX7i190lGBWL`UU[0mcYl:iDSc
KiVKPb9YOhMh:gqnP]3\hpoT7GYA=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FACS1(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;

//Function Block
`protected
=_]Y5SQH5DT^<?:l]HkF?DbRM<WS5`f[4Yhcm8BfVFmAf7b<R1ogY<nmRbMB7\Wa
pJU<Y8NXQL6TmJ>TdH<H4pcB9T@ocdGk=]MFFpLjkJKQpBImKK=p1?j>el[jYhRO
J`:3[HD1W34b]o9H?c3qa>YhoGQfYmYYe=I7cG0=VEVlMP@I<=:qGSPeHmq9<bE^
F]Pg]keUXlP5A[Bk7NoL:lZV5enh>\kYMY4CLnM?2_RiGn:?E<Gc>a5pe1kg6Qqj
:VK6nmm=;Zd0`Q:oS3k>_>QM>CCe[1lkabOR485Bdk_IQ2Sq9SS6<Y4LVPgTb^8F
3NcKB2Kd^AXcPBhqjG^]d`c@kfJVb7=i6j\HHGHFo[KWK<D0\:h9plkA1S;=J`cO
V6C0WC5h1N4S[B?4ALjlp;ABnC=pcdNKKC?PEoBNKZ\UQL3F_T<_oNRH59Sa1H2M
VlpCOMf`H8nI5Pb?:khM[iV>UmN`CDEB`g\KR[IqVOOnRUq`]1Ah:K9QIl>UhW;[
ed?BV8CVL`T03SmZS8_]Cp9n_d<InILQi10@I]>cS6[4mKEi8G<AlLc4>Kpa`kfV
`Emo?D6ej0fJUk1FV:A2BU8GNmI5M\0MRb9M;]U62CWjZeV6Tnn8EiE<=3J7G1pI
hbeEa2q2T0YOip`j7iHU0^ZbYhhF11D8;\Aa^D63hL;Fj]K83]:7V_VUd:EKgB@F
]jWMhdo26X;P^]KREN3;n`\lX2a6kXjbXE3<h8;nYa92P[U?51MY[3fM`^a4BEjU
ZXiVh9<;69Q248PeQ1`AG7YTenXRq`<d2Q79oIXo[nhcQ9X5kE:a>nbX111SQ<Og
4a]JIC7k7:o[CiRiTAkDUS3=7RUYGH?l8IA3jKF?BBhEUK]QP35IPe]QN:D^mf^c
EhNU24WAHhDdUSadWN_HDCP=H7f>l5mJChn\fX:F1`gqI1JXe>;OeSd=7d6Lj=h_
V:al6X8d8E>:dM<mB@GCV@;`99=J[7Z:FaKJ<bBQL>61Wh__LGZf;SA]k1O]=LFQ
M1]Rh:74ln]`ZKKIH:MG3Aa2UXeJP<CGO6LkI\BaYBFYUkTH?doR3UJWB`qmOaKc
b=AKfF\]Y\1O[fQ8>PB4jZ`NZ:53Rg;_n:fha[\^NoJJ`Ch5\>17@W7Ok9D<HnjY
<?IR7LAT[FXE`6=E>\PG_d?\3?[V]O>_i;]gXED>`cTOhW\h9JLi0W72E>AXeIlE
P>aWK6gHVqjF<58UNZ2Ra2CQ\ReO]5CBI9nR1MLSCMI8ERKbKHf6TGki_GP911RP
SjV;bRdmDAU_0WP7`^PCPjk@>b_1c9MAcc0_[;TUFi6QTKo@RK\<_BMC[S?en]>o
edV:b1d]6[6=RGM=R1DO`3Jmq3:@fjEkSZhdhL9fb\i;aTDW2fZ_PBdI_J@jQTO1
mG^4:LUNo1R^^jYfZLeX7S_mZ`AJW9Y8KUCL6\MDlFj6Ic2eS0ZWD;hY6XHYBgY:
<TdWC0H>a9^[S_T[QgZX^KT\=dkmoYL\I8IblN>pV]Fnjk<\04of7gDa2k9dPVCX
_6=9qm>S_I4;N=6L:R`j`:=maSiJh75_m]07ZKS=KbWVR3SYYLnOIGbg]1MLN^88
1`2TUSO05b^9C2_E^@iU]A3A0hOi>^5KbQ8llO0Tml6l[Y[P?eceSmj2E:;PJ^o8
Z`54gj307@hjDLNI@=Lp2GO[_1YJSWe_WbLZVP]a=Ri`Y<5l>1Y^H[_GPnYZTekG
7?WKl2AK@8B^kOV<G@<;INR?V>29TTD8?V4Gj4[a>4<Qc2c6W=m`[G>72R;a>?ml
aiXDk;907WF0bTVJ3DohoCh`BYf>VME@NMp]>ilZVDOOT<OZRHBE2JRbL1BcnKFG
E;n1MRk6hBLoZ@ZI6eI_\Z7EB9iCJI<d?RKFlXNW]FVSbQA;nc\g\olCa\M5oc6O
Ziq1=@b2[NMJ\@oQb=onLALok7bU]\cUYW1FXQPG_7N<]FAnl95nI0G]RN@VB:RI
5=DlDElG0XkOjH^T>TN7mP=kZRA1_:fPiW8LB`5JTPAjaN=3e5KEX]Bl<mYN__5Q
c4?SR<ag=3g_YW?jQU6a1iIb]kWJ2p\MKGMWT=12ab<b38^9Q`<Hn:ZDYEchBX:U
mKV>LThM2JT[09og8OeRSfDBTP^5WF9;OUN4afNNcjSMY13:Z1]o^Fj2Agf4T5Pa
m?dJ=L_oMCflFQVDCe2h;TQQgRf=n_AL_3<IYnZgnP=Lh]0:[mZ6WA3np8egXUJ:
^o[3SS]L2HX_6RCR386=E;lT7Z:OTFh>9m;_2?Wm3]V<C\87`8L`B[22IMaP^i>6
H=734cEQOE=Y9@:60?^d<RQ=n]YOlVj28E^<]OPOY\G7R3Nf[6cHXMJEV55A7Iai
bB:=:@I6kRSJnU]DYVbp@_1Z@6i^5[P1eA7l_hOE:VdcU\bRQQ=7D825L;_4G1<?
BSdd9eLh`GfDLm\b_0?aD@57a_UnqbVo7Tl2Mc_ESid5ZGn\?RU]di:\Xnf_TUcZ
cB^PS[Y5k9BLkTT;5aCN75o=J4Q@0k]aA@1<VE>H2MT9_a_AU<60A6A9aleC@X<Z
SZm2NT9KER]gWF;<1Z2G7Q\Kn`^DGE`TLEnQ^Cb8QC0]K:7ol[Ghm6`p9_ngmEa1
;Rl:inEEij^fhalYDcB@OEOZiYG>Jaga>HYdWejM:fbAe=lUnK4IGi@@UOCnD[[U
8;iK0G<nbW<>T:g6o:kEl[2U[79Iglbhe]kN^n\D:8FmaF3n<;k=_hKk9X>CkGA]
9K<JM0J>1QAlgOG5ISUCFVqY_59iZE7=Q=AiN;PLbVKn]59M>=1^gng8G7^?Lf=l
b74T_J[gNC:Nj1o9KC>Dj6loT@g7]1Vne`nSiV<]em@;:3D@<26M:>3jhA6cgDHa
ViBbjPl<WJiKCaTcPd8M^;mYF@b@5OlAmIM5fSOXgXJQiR@2kI^kiqA`I<JSW9]M
d8Ke=e4SbnUYTaGSLb:fj[A>>a09ENoWlo8@V25mT;OS9amAU3<>bOCK=n_:LXgd
K84A?En;calKbKc1mDJlCc]ObKJjKnaZaeQV8gFVmL?:UD@i:iPok8ARZ]F=3[0f
>8T\anHdo0ZfcBX]Cc>WqTn[1Sa7Pf?AnhOF7bRdD79LAEFeOXX`:>VFOd]W@YGM
72[=`ceZdA]TBP2Qn4\_LaM2[JmhiY<M@P2YM>WYA0H^1^ME\hGVLQMk8Koee[YJ
E@OITXUmQN_9<KJ_ndWIET74jIAUFFPP2RbY1Ggid]Gm\^KlTX4pWF;jZl7WfWF_
`ZLe\P=FZNZBW7?dT]]4\^8QE4iWGF93:FGM6md9;jdCHOCYga0leG1S^^XoN\=l
9nAT[e4kP7_g1Zj1>Q\Z50_[ARg@Tnkb14Z?3^]UF=UkVk7hSI7^BhS@[RjHgL];
Y:;fi44nd4EQ@_q9^YDFY<dPbSQbm\b2LiR5Y`dCH61Gm\@nXW6HCOHhT>nc\knQ
fLeKa0GF3:UTO7W3Doi\46ZDTk==Y<hj7TdXEK;?HJ:Nk>b2cWNHS1Z8=VKdK8d8
g:eV=OVbMdTeCBEFM`<JGHGH80X8G6^Y<RBgnDl9;p71K9ejSVGQnAM0M2::3an@
^728mHJi;Oq4`RTgR?oGDVecRU1IP`QE9NC<c[ffU1^<@Ui=e9>U2;db_IZdd\94
PFXeO\TPT_Z8m2lhamoJmQ6_VomFOaXj;B=Q[jKUDVh;hUi1\?A\SV<lRjP_OZiT
QInU4AQCiMSS8?Ve0C\?=LacfR4bQodZW3acYpDDd5_Pa6O]n<_;9_GX_C;C<>E4
DVV0mWcF4n]39]7cSI>Q08T`UNNiMcc\eVL]leYPS[nI<El6bE?@lOk^XYTdd4?j
Mb4cGLVCoYgdiVe;`ET65IHcm;UEi9M@O_UV_]e25;h25ea_`kEfPhBmcaniM7h^
qSXQQMAK@SoO8imG??B0AgNN0>KSUUWF_>0W3RYK>DEKh068PDXSVOO?GSY7aWcG
W8G\PUE<bf6VUfnfa=eaC\NlXL[@kYVSH=dWR96Gm];4[2QE4\[NMk5V?R8LQSgU
=Z`a=Q60ce1>SH874ceSN7AY0<OqoA2XGcSeaSgchY1`^F3]38AmgZhF2@7P@UPX
8LjN[@Vde8YWid]9p5BNnOcLaGJWkBdZ2`R8LJ^R[SWQKN0AV9J5XB9J?WG9c=5T
3cec087i88hj8:3RcXnn=f]lFXm2o_k?9?2[1M^2@TWVl\HBHmG5T0I>i`7bK=X7
iGHfR\j=YAM<Cjl1V3M6>W32@YjXFIGPX8dT;7;>DQXp\K@k]^SJjIa^P9d^Pc`O
_dojiCoT3;oin5?A]e^jfJ@PGi=l5CIj_lcGRMXL`b4TmMSQe40A`LnFk=cNP^A4
_dCJVlS12FB5D3?F2b[nb6?S9GgddbU]U2NbVS91kcjgS`8JfARP[jWKJ2k2<jC@
4VGhnBqHXOW8:3[a8_fAd:BBm=GDkRH7@8:;0f7`G@J4nIl9SM<ciQ>iK?<TUUJg
dcoGMQ_`4MQ5l_[hABOFMIh\jH=]k^5N@30bTNB=e@]Ho^KNQAgPZ:EMS:OZP1JH
;0k<C8Id21J0m2OH[fo`U_UHE4hbHRi1Rq]>LocMKhC_hg;FHmU=KAHffmQ4=bEV
h801\K0idEI8A\?aWbJVDW61LNR^AOf7gW8_P[1n:iX2Rig8SWVQ2JbfZeqXEAZo
b5]gD^Q9Zlgm7S;e5D]RAgbn\Z=o9nc45SpP590a4`L[:<Q>N9@i4A^4:^db7?Bc
IDgXcQ;cfSF^MWN>aje2D:W8Nie?6Fl3RKPKQT2c@mG<P^iE8=bUlm8g;Rh1_[[;
W^<\^?c>YC^_W`QMNWnBXB`AG;?;AO?_TW\PDWF1meY=AQ7B;62<6M=OR`ASj>eB
2qDh2e2;^mFBfEGi=liWI77F4S\JZ5V`acjD8<`SU<YgVebea5mM0c6J:kgDL7JI
7A37VS[d6gbZ:3cUoN=ZgWm0o7R_k`kMPah;:nekX`=\RSk7BH92l6RV=`VCSF2M
l?DCU>aZ5FC@@BlS3`mb]hQIanWSbckEp1aPGh@N2@OO4S:M3Dl75k5>2;7M3NK[
001`jBj;ccEJ`UWcW7MCnAbEkV8>K?oMQi^HK275VdbINBV>WZ;HPK7OE@I_NWBa
jkN@DM^\1EZ=9O`m54imol3MUeMTlZFD`1738S2G3nmZl\b0Z1k7Q5AQJ]G3mjMq
SjCL3i88oW:2HN?R8R22V:AKXEG36Dqgj:_<;<3So_kj04?9G1GS;<g8kl\foob8
Ji_A<e9^DcU:C4PYg;>T>R=8gmckFiX8B[DYXg_EaZ11l5WWdb2_80lWFRM>mmlO
k4A>YfX8oQT914cRHm]7HG4^A3\2;nlgd;fSZ0N05f0c8dgU\2fUfGEPmIibopf5
bEL3U60=6T>:=eCJiPTeSRDQVj1=V9Fi_P5k^Lc_4ZDFhKCE?F_?d=\3ocBl:oa1
JDPSUHDTl[`fomQ1<WemOGmlJ\SV`]:JC@D^IeC7gJj=naJW?aP28M_2XV2?jjf2
nG?55WZ86k<@OQhcCE8Gbk[\34h?po;QkL3NeKXYDSamO48e>K14_a?5_kU;[2A`
5]M_K5A\2EoWAS]5DNbDj:A2SeF]@md@GMho0VS2Sj_JU;jY2cK`K0bWg;AO5m`H
LZ2<PU9]D^;G`Kg3aJ4TP`IC9baC2o\8dJPCK;T`COI>GlTYOZ2gn9[EJ]=pcUCC
oaDXF0I=jb<7=QTiKQR5N@0XA5[h7e5YgGJ4jJ=mTFTjWkGLN3i;R;8>nP:GSHFm
0`79XGimZD@e^f;K@W5AaEgh\4FL]j^H\Lfc7fkVaOEZ42CgZ3dDY6LjDc1Mc1j1
3mOQic90\ZaYBVLe[XMRBOiiRWp`jl?D[7G8kefYicMRk8h1[1IOagI0D_Y[`6K0
X^Y2iY5THKfZP_L@bHo^M`MTWL>eRLJPO23I8b5Lk86kLRl:IcNc\01Yll[WVaL\
>@]bQGB=FQFTob:@9BP47MYeV]c`9QQ[?lgU0S?<0ocYH2^=Z=nITFQa^qjG_A>^
aHSYD:Dcm\LjEEcPK3cOQgfE6B\i>IFL=R`V2W65QQo:i9FWDZ^n^TDiORgWgdJL
L:;o:G:P816E7\B56<K0iYdW7QiKi8IcNWm:Ah]4Q`E4W9TjY^cBRl5ndCjnYT?U
60jlSXiQHk46G95jbMZ61_Jep`dj?[i<>d4732_5H<P>X1Y47g?@eIY_gNkD21Q2
W\5m^6aU@:Y9=3fRN5He<1Xm`U34cRL^Q54hX?eU6e;NMW3;VF^]9H]H=\:_>ODa
Phg8J5Rh]ne`^;CiTXoWCX:Yc`Tf;lCGF2WPPFOoC2>Rh]:S=Yi@;GHqnF<D\Bbj
ee5OJRYN48GHAJ0P77Xn@T3WT3;KSR8Tf?Z3VRonSAAkICXcOWH`;7Qqk\SCbB0j
Z_>^V79883;P:4WPfRN9k8_T@DObHa=?1Qm0Z6l`0TaQ>kN>lc0g_bCRRFdA58@U
AHLliWnX2kfVjCbTOOAe?lV0K1hP`:ofeO7Y@dEYRNlhCBIl0eRAZ=OQkZ5P;:4c
kXBP\RhI7BMPf;aEiJ>LlhpE3NI;IHO[dFcM5PRPT4<`k_IG1cD2@Jl_J>8T8`XQ
EKkX6>MCn`?i3Ao5Og3V6Q;M1^ACci<kcT5KOOJT4GI0d=<W8HeoMGbQ;f=GgnDa
^@1IM5MRoMUelkh;ZNhco4:E;BjV0WV]g>U]?1[o:\kWbbm<9cOY6p0l_ib;oiiA
L:X[b9c:aXeJa9]aKM@3gKFELW61D5QC[aRgTOa_V==_=coQM1ggPK>Od:YM9REk
oZZHPUN<I@aC><8]HOLhOAH9dlmog8UTGDchMDd><c[[DVe;]3nL3Y06nP^m6JG`
g]DAmoj:?]lR91L1g]DQp6<68idBDmCGe3^S<DjDH@L<KcKQ9JAS<BaViN^QTWN1
n^hc[3f5SCf4FXG>p_DN2[LMiI@BeRPMg_?@o<eUCRRJnCRUTAA\A]5lMLZP6>@O
LeQ`\X@[Wld@kYQ`a8?QlFj6Xkb\Bin^PWGJM>1[o=3aIYKAPTJLWHWZ::;8AL:Z
>a3K36>TijLdYZ<lk_26S9?lR>V>amcO@MO855mdiXfk4]4q<S7GfF[0NJnLnChA
cgcC[2jRbdW;@;Qg3:Afd^U60SHS3H2H5PnNd>ggX\=i;?VIIN^0j2K;UWfY>8Gl
O]TO3`IdfFZ:GAECV?_LYKlLlF2jBLO06KI8`Ckn^4N:k6=9<0;A374RE;9hkn]1
:RaASK1h`=6cO<pI^HKS2]>N7XHdC@Zm6dK\5@NTWC?YT4ml?46N?LRDdQQQVEF1
_a11FCbHM\m0e<:;^n5hR0dW600>WG\6BjYD=eiW_nENoBeGcXkQcLYa2?TYWY3o
V@cQ6GG:kUDmg;RI73J\FT7GiPi2NQUgSWnOmN[9WHb?opgJGWA\oP_UE^AdIn^f
EIUb<9Ld52BYPe^J>?;HbCnCCVNB>9YkUZR]11=jKDOETSW2Con8RihY:L1mMl^e
OiNgLG739Aqak;:G<7BX39D=V7dfPAL^4NL\N^V0607`W[@@7V=@G5nLZfak8gac
8T\ULF5B6?6GD=_K3@BKEQ=0@j20J6l90nE?3@F56LbH^e^ICa\nCcQ?8Dmi<RJ_
edSk<Fj=lCebm>f@RoABoiT37pY]Y<PBRdF8jio<R0RfCER;2>?]bY;a25LZmW=a
<3TBqH8cojL7CeO;J6lb;80XJGYh:>RhAVg>EoDdoAfSO\JMbK7d<j0;V74CDOgJ
b?GUV[3XNFP67]c0hN];eBSWZM`?3C?cgY_K0^@2cfUCDZM8In<1ABA\fBM16<>J
1_dN1Co7]`hn^HnVUomqB1C79DWdZLl@34j0Jg47i0kWM:hbRJKSf?7FYWMCF5JZ
\K=[S=joP5n9?[^5XD9WkGQjD3Y>kI8@jPakGP[aJi`Nim9O8;YSj4A2Ld=YPLke
^^c^]ZhY8`AhhH^50?odSGL7d<LLC>aUNlpZTEYI8R0QJNIGchlc@2D9^\D0;T39
787LDGQiJk:?fbc^@Xk87GQ5GkKM8VVZ[I2IQ`O[Hg[`c4e81_b1N95:@3YS5<oB
<D_02h2bTWnb`JGC;aJX>2gePGMb3V:Sl>WkCM:O==jJWMJ<TpjlDI\_OS=Qjhnk
:5k7^QILg;E9ke\V?kciI:pQLG2>Jm<QnhDM8JkPi;<4oV?B6hMF6d3P2lUX=fRF
a5lcgda^P3_b;m=dYefg_aECXL1:5Q@mlMm:;6\Nl8V^E`Y[1odL1H?IWPG9U=VH
ETNjLnCA_ekRM276Ce@2DShcb9XbXonlHaPJ>pJ:8E@>GCOSCC=XPhRA?]f0R[YW
oHK_BLm0H:N4naEO3cm<iCTOW15RW0PcPL7Q[Ta7G9HmC\?E9@KWlG6AEc=F96Qj
=eER[6=kCCa:_3ODaPhg8J5Rh]TQ>R:CP@7o3LH:XV<CGciL>hX2p]JGB1lla?FV
O1d>;D]bNO[=Q[Hd?kVWZ4IAlhfoRGf_6I`:;UF]ZWGV2N8:JCUmI3E<m5l`7oj?
E>VASo4J3bVC>;88WTEFUS9;ZCJLWHWZ::;8AL:Z>I7@WE>:l7jD]d<MjB:PnBj:
C``qEjMBQ_en]Hih\eRcD:=]18b]47>gNQ;J_0C@=UH9Lj]KdOEJ5[^?Ck_FHLNi
F8C:?Yf9Ni9P@j4hUc99T:41H7cBR>I3NESYPAmU@d=93K^>>He]=0g@MoSihbNj
F@hKhi4>EPmoSTR0YJpCJDCE2K9kYebX>=_k6YMcESK;?[2\LFQiJO7Q53M164Y@
S_[K_k\C0hNq78`=O>U6UMNEVbFfY7;oN@8D_c^B3km_9T94`L^hcF4eMKeCXaeW
?GMP_=>NiI075?T\Ug2>nIK_Z>1O:7?9\n8UI@fHlf=qYE8_nGan4ID7oBZVAh?[
`0PZR1:Dikk1_4LG]0Fk_j0i@1m5MVOMc88CPKe2_\T9Yb<MZY@:?\SDg4A1ES]\
=e<]F1FEd=kjhjhbkm=^^e_NVSH37o;;c7eC_SH?^Uk8LKGYZRV=e5m0g4A13bW?
oYpG;PY];MWVlGVf^UOj]RIK6@Pjh]Ud[XB[X>jmM<Z\ZU91DMWk4_RPXH4CF<KA
I99G5XeU3\`JKJg_dO1@EFIOZXk^hO4f;X=;4bQM?SVHGbKQ=mi6JO]PC_Ond???
nS0jP9O@Z:D8X=P_dO1@8Ob\KqbaM2^[kWMH@XfZ2_m@W68JX[ae^^L9Y<E0D2Ge
:YN5JbF1L>jfgJe1i<oZc]II1lbmB>Z@aE\3dQ\<[I^5oefBj:^2f@U5YjO2SF>F
ZQoo]5\ITYKl^5embd?oS<4Ge1T:M0:A;[0h8A\<[If4VFlbqbeSkkKJKF5TK\>e
?hGSd5[V`bXYBDboQC8NYhIZK\^:6YI::@jVO;aDf<7g7Rk[@blH=3MYMN@L0?Il
QS?<YAkX0IJSQ=Ro;:HRXhU@ikkU5J>k@AXiW;_^cKGH=RSbSO4H7cEcg2DId?Il
QNVY=UdqDJ>@20?d8Ylf5`]jMm3b88OaXQHJ]:lYX0BO<feKOhKC08[Wm\l^OUXX
jlKhIX32DAHkjC^JaSdZdHj\H4E6^mcgZEHETOlC7AT=<kcKf`QBZZRSDa5LO09f
g_lCkHUkh6Ki=XH`24eodHj\l3jb5hp\I\:eC^lj>Zne\^VbJcG]]_Q;9eXTU8I8
fcKKG9Kh0o`=IBMlASlZ8G82IPP2?:d\ZnAJ]H5hdH7Bk0[nUO0bjCRElCF^d82P
e^0QofFf3PNc\D^;Sg=Z8F`PliRf9VbU3UJInM:]C?ZBk0[:fHP:0p^ZLdjX8NEl
4IFFS\9;JeWVe\m7@dFOH;?Le]:3bPEk13Wbg@c@<76MkU8K:E:dlo^Fi4eB@cMY
WKM1do0hS6FPhHg7Yg3[HCE1b`gbPN]O7WJ2\DTjSf6bZZ<7Z:gHhEE4F4@n6S;P
IXM1do4X<l@6pCcn5m^>H]P8TZW`c`BQ:;A66Vom@8^EWY?EbYOG]`YBblKUJq;_
5DVfEm_`om;cU<UZf0N60`DAdQPna2_UO\VJQ9eZ02WRE>;E;AA\AeU3R8G4KK;T
MQ9S@JeP\7KCTMU=3Pm>jMJAdoDXaXELiBGCC0^lT[1hYTW5AGAfba=aJWZcWW2:
X>[XB1\5hBKCTM;ViYZmpaWX3bnQRiaGnH\kYf1iIGEi_kW[W26B7B_hT]o9AhOi
VcElf8Ann9i:Nd\j\7j\UaQQ`hSEJCc48ZS0PbQ=5V9qSEKKmG:iK@WFlNO@bM7j
Vg1Ke2@PST@CId8LCT6EIbd8fjQ3IS^6Ej67Kae6:V;mS3nKOYaR;8m4nY4hR`CQ
BYUKS7;W]Xb\eHCf9oT3CD9_?X_EZCVRd^1qmh8DiLZ>@:9^9e<Kk>Y:;Rc\SiCn
k@ZjGPWB?0>MmZOF3:\PfX[ZXZ7JFQR6ZDDi`nW;?RmSfNK^[>`hnFGG^mK=QRV=
I;Z8?gY_e`_bQ=1N:W0fUc=]Fgea\Y[p;eP`SfKknTl;nM=lo<[\@CU64N[9Dm7i
Y0]MjR^2K\JXSG5XJ@38V1>jmaj;iO5Y@BPk0=SNV^V_di_O2YQ=GUe_9cDpl:VH
dmH\\12clY;F1VbQ7Fm<OG3;c1Nn<LDY97:@95e;JkiQ3\7EZoa2]UGGGTbC4IXB
Gi8a_To82fJ:^E5]B[Q9=c_G_fNeS^;[giDIfC4BK<5K3gh3RBaKN]4ph4U[X`bK
n`BHMWI`^K\HGQQU9X<RlUj_n:cQ[Z[8O`DcWcGdThIPD>Y\GSbGN`kWNPD=Mh;q
Le1AT]KI?da9Ek13?gg@W;hZ`XgkKFaJ:Jh:I2E`PWNl`]\>6dnDKfiXfTLcGa[=
GT3JdDHjET^gkcjC_1[gT8BZhk97O^a37@P0^aAOjY7HMbJaPJE9HG6[TlepI@Oc
NMME0>\8TU^4Wa2K`f?<fT7\aWj]WS;0RhWaSSX>XHN44;OjGc^P=K?Im7U_nYCb
lENSi:B81AI[Y4V0FM08EZ<qSF2CZnohdal;7X0Z13]cDodgDagY6K?\1L725jYj
<h:]nMSAc5fT8SCY_n3Ifh2@SgYkJR08TU9GWajHI9^Eo?b2NQcN6K9;S>m`cjjo
N<1kkVZIKgNDTGnqbeSkkK;^F:TD\>e?AG<;5[V`bTYL`bo;C8NY]IlR\^:6Y@:m
gjV\;aQe<ag7Rk[@blO=GP:2NhXkC9;B?5;P?ZCZBYiiX:;4K38>Zh^LOWCLKZDO
ANi9=ZOpP13Uc2algo<?mVDJ3b5LRThicJQ@Z@RnDL7W^GlVT`M>e7<jY39@Kik[
LP?CaQ<OPR\b6QE<B6l2V^G\FM]GQ0P4dJp`0KdOjY@>Ig78X1R7M]3=5FQ5dRhM
\k0c5hS6M\DdjGF39YOlK6UN0DW[]RHIDfc3=3AdW:0HEP=MGVZUD=5K]Me8o47d
maQ>mml[^MO^1U3nCJ3TnHGLAo6OhKpChfJi\X<CWAjmnAGK`0n=Ia^WB85PMDX=
XdAR>e;B11SB2OWjG``6?c`\6hbG;T4CH1Jh>b1Z\1dK;F[eGTfTc]`SZn3dW2h^
Hc\4D<jQ2TQ5^3FX3fliD<qk58ML96Sb6>_8j`@E:UFMZPUN[XljCUeCaQQZ6<60
=3CaU18C<XcdF<hYKjIT>MBkgCM]5jT_<Y71`C:S891mm=pgj:_<h1QS0_Dj04?P
81Q:;<18kJLco7H8Ji_A<YDTD[P2G08>B>XF6g]djl4C^UBbaiX1F<OU?i6fJd9B
fJKJ;ULaNVehOKUkk4c>YfX8oQT914cflcfC^\@abQp=n_:\Cei=:>[IHk:aHbRL
YPVq`;1\fReB=:2QOY^:od@lIeCjVBOEk:fM5@gagM?FHg`\2>S:Y:h6IVh47=VV
8eb:eWInV2OBBR`fId=K_MRUIMi5f6C]^\ZMR^oHch<^<Dn002RU:]e5Lb<U=Icp
KdL5aONf=8YlNEnMM0A^2KMZ^HZf]bbVZ5<eXI`<f3gXFi940d6DCkgE9UNUG;L`
hGC92[cbhQBP1Xdck9:HU]0degCpb_G2PD1TS2d:8iCWN=`0\8_H7XE@=F6[2^P9
TO@ID9CJcoFooKf\?5eCBeE]5B\3b\>Wfh13CHo]k^oSNS86dBX]jAT5kA_1GGZS
\ihP]M`Lojl^lV5PcoXqCFKXUUZSQ^KQUZ=\j`:\mjna[Ke1UD52ZC]7PifHNH9P
6cYlllUP?4Y]7R=4=UJRS;>3Vi_pFFW>MG?Y=UMnjT7eM8T_8<@FGFWBRoMnU7fA
d1VUfYJOPc[L4[3E2KnZ\FBbeKTPFX1g3EeK4Xi3anm:m1]^K<U8U]aFJ`WX1^68
c4I1jL<DYF@27BM]nF9q<\ehV;T^IF65;L>0D[01dOWb]Nl\Jg=2HHQ[Sf1hg]8Q
j3oikeD6i2MA7GoYbXa[<>CV@<e1iG@@<Id7onND7^E6k7q\99Y:aq@iTG]2C$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FACS1P(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;

//Function Block
`protected
1>5?VSQ:5DT^<g`a1:hhbAUCRdDn^6F@QP\?;<ceLDRRb:JP[XI]VBE1TE2ebo6j
W`UbIMF8B;\kDhWq@8=@i0_^EWcEWcZMF\Gb^XClLAPfW4De;9_Nad[XHI_hLQ^:
MLO[moHl0Ihb\B[5Hn_>oE[Zq1`]_Kk=TdF4eV\WGX>kbmbRk_UamLIV8VOQ38[8
adBVcnT\pe_j_:?qUIHSHBqHdBLl?A6O=:hj5c[H[LZc?RK6[AIOBZpOQe5Uo\m4
Tc2n<:51MTgRCga5<hPRcFp@M6AZ6q]iU:j:DW4UD@SIHA_cIlR>B_m6<jh4L5QI
GoVaoEcn8SO?:VE>jTRk7Bn2LjpHT[DE=q6jb]\D]aSS8G^UZK[I?MFTX3SS=Dc3
lpcdJm:6M3g[gbAXZZ<OGmRJ;K;Z=pa`>m5e9Z>\jWk:WW2]4T;_gP\32F>]7TBP
aeqW?cUU4]o[lU:<C@oRjQWJM=06VD`6n3qE:677Xp;ZV\=U[kgmgA53lNAY`]A^
ghJIbMoff[:[FL4<pG]A2e@7LkdI_Q7_NQYZUbV7SGh5XhR;SRAD7qF[AfGgqYVG
c\FAZckO6;g]I`CbHa\?^IndOPkm[@2YFBhpMTbOlgAc_`0QU[54LZaN>U@^iWj;
^LFjgG?[pSgYW=iJp0mG=VFf2KHc;V^Vg2OZg@g[J=hKhIA3Nl[>eSn>@]5RVqPk
H1ESq^BN2X_?OcSOB<e8X7J=c6<?l:XBAQ4\Bbb@DjmI@f:m@TEH;hU]Wn0CKAVP
N1lDBO`eA7EZog6eB25[52iPCa@LhfHgen@BS?Paf8EIoOCXjF<kI<8IG6<;O>7P
Nm60RD;8L^WGe`=faP7p<4eHY9Co`Jcn>C8BV5SPOPACLja0`dcMoRZSSObD?DgX
j]^=jX5?PR_5Ook52D=JHW3:fcia<?W5FDb9R5]884c2V`YJ?Vk=bA<EnT^anKm?
dIfj;mgIZTK=HGk3?dLE15j_`?WcBePQECqc_Tggk9M]fZ]j`BXTB2AS3l9GPZlg
F`_\oR76gKT2mX\qE2b=e=ML65kalQ5\^`LTSg9P_g0UeD66Z=R><H@J<6GlcEC4
@0FE3?P0^X<I3B3YY6:a35ENI_^=Q4J@9g58Z_3AP@g;[:dFZMImnBP<nm?9k7<<
3]RQf6BRdo<loD_81kK8HGhNK]FQQ7pmYj_^DbEm?:Qoo6F>`8j?YOnZdF7foea>
72]`<IJhAWK<>gG42ES:KdfnSa5Kl=NiBNSTQHYWckA6VV20`a@f?TOf:e[fC9?K
bk@O3eQjYh?dG2^8@kAHgK8MOa1@QM_UYRg[eoJGFW;>Bq_OALnDAJ<ki50`V@dj
B>=cdo;Zec9TJkW9UlTEO]]IZ0\@m=kU]bid2X\lVV;]cgkg?]H]Z:>5]XI=f=_a
L91\07Slk?NQKA]n@9Q]TE6hKmAj_4Q6oWfi<enMVn=JL2J8JJ?8_Dj1C>?kpXg9
cCJO4?\]7<=H<2`b3a=H;5\<@n:nEo``hilf>N:M50Te5Ko;S1JkJ1hBNf`B^mlB
ci;L[eUN^;c46i`;E;Y6^OgH=B8D0oGI8dfSaKRXiU2539CWg9k01F:B=nO6=`H=
HFbkOS[QeXdpb8k4G>ohmDWVGgK7;1BoPim:ga]SKAQ85BngjR`lS9Dd]@B^PY=0
GU9=ACS:WC5V]8UPoI8FL7lc3KWdA8AZ7DVhQj]eKG\bdmj\m9iLCDoY[Tg:34W`
illo1SS25_T<HcSQ?9B@DPXc@Jq45?lVk1Fh54>G7dHfn5HPmT;Lb>9RIUS:BJ6j
NQ]FEYNH_fdCXN]S_6\OCD9_Jdh?UiWM`gM0FM>OT:U=n;H45TZG1UaRl1\2NUDi
lbV66TO_K?aZg<_e_SC[UD5`kED[OJ572IF3mfg51qd<4?YNVFPCa\ZYL@Xk9dYg
55P7VRFN@bfQN5=@dO]1:iKbDl6HA\NdORRL@>CEqIGB:ac]]D>Q6`1a^81]2TYT
bFhH3X:iEbCYZ[`WkXL[2FLQin4a1egDj`6XAh151:h\EP0^fEL77l6Q\E1n0[`Y
LT^?G23Rq^i=eiggF@`N5P9<=0S]9CDPI:\a;J[ddnh^R2=a0EdomZ89]8e[KlUd
OQ\ao@@QY@A=B3V[e;ceF9W0m3mU;dlT<V>TlCZg[5?iKVK@Fd97DnOHR2JFbKEl
AZ<H?b7j=^XQ>TQoTn[anLCKGO_^E_L`[c04k41pP;k3UkMUUA>jc8R9OKi4J5C^
:GN]`>j9Ra[gB;Q`nZ2;GZU@@mZU4PSh7GK2A0I_ImfgV=`@EQ:3UWD[F8CVFkTA
O_30]<KGlF0g>RmUDOdTH?f\OkR5nJ]I<n;oJ`J[PR[UK\Z\S4Bc@^A3<PJ^ij\N
PE[O1kqd?`ICLH4eg?S=f2Z9TH5dZkgnUmDD]dBMFf^92DG9Hc051CnRBhh?_XAJ
>Ge0aLY<b\nYOYZ[>C\PgQCUS7cZ^n3bgA?T@1`X_:]i[lATmSH:Hf469TcODRbW
WP;`H_:d@DZQW9WVi[1\Um5YHkb_fUHchPO3aqDM@3oP<jE?@ZgX?cHjok]RcHF8
;eP`>pT@dh\@jH1OEDV1MB1G^T6=2@2TU?eE@ODURR[6[J:L6L\fMSob8Tf2IIH1
bDl?V5\9JIHF0;c99:J4>9X?3ZUBU^aHLFThFJ1IO6Hg;\iBCRBSYLE9cK2h?EI7
g];OoDTOWBe;4VSCLOMKTIj]EW^KHe9SN]=npB5F[<=kO6H2:8bS3l2<4_>Jd8f0
]aD4cdA4^Q0@05IPSVKZdTQhR=`^:T0WT3XLheiUM_fO4@3VHID5]>o>L9JOS\3g
UcmG[kO>[4_b6F[M=E9d]EkPCkf\aD7^XEnC1BbI2o=^gKLmN?iQCY<V2SI;Y@93
LZAq<kLMe@5^Ida5DM@L[iiG7@g0;@^O=mjL^o7cbH>G;X@Y0bOm55f17Q=Dn3l:
im;YHGa@@<jm<\4<oMkn?jf9Ii8eK5Ld1eBj5bdhVmhQmT<@U5F2gbKf9`Q\gfI`
QG1K<CFFYRg9oEaedof4Va9L0@RSD5NEg1p52_Di:_^Jjk>Mm9F>fR6k_0AIi^Je
WXHB2bPMM7oeeF6j;?<N4?dZE6JA@G?MTX7_=7W5B=@`aVX`DkhCA^7ZU4CR]PDh
?JKX^F>;_=h?PATIQi8ed0bP7BnoCO;Dk7>51EZgY9MifnoN=TX@d2nUE2TdinI>
Jqg509PKXgYQY]e\KihYia3kSFF[:CDK<eWhCfZGI4<VS8N>aE<JF]]?I<PRZ_Mm
2F3?WQdcbQ@mb0d4ILHaBP78n`L7b\A7Ek_T:>6il1Z@9el;gIn>?JUgdh`fUBT7
gagIfS8`\MVaeli4h4FOnQED[m54jS;IpaWX3b0Q^iL@=jdZJ]DeKWkhXjE^[VL^
^d<Beb1cC4T@Z\WYD7>\T@bZ]gE5BIKB^20L93SKBCmb=ZG?dAdEe@9G8I?34oGB
gA1=U9ni_6jjWNYfQjgIW?f6k<8\N2j?CaS74]m]gb?lAZo0g7QRR\RTA^IlX?Cq
]Rcl:2DeYlKID][=f>EgcKb07GnV1\liED2eLAB2D:3<Bhhn>0U<QDh4M8Jk=9;l
9oVeceXT<AERPWWZ2K=G=lDQj8nnA_ekXfd7U\0Ia4MKQ^Sg3POmEH6UU[h8gonj
]FUGjAX?BX9UPQl?3_gOE]TmiiM[6mp9DPUINN=AC`leWeG7AWMjf`K\YDV@nP:W
]k2Ql?WM`iQl7;D]E_a;<KcL94TIfR^Tn4YVfkG3T2BQB1aam`U>;@[`:H_PFaNY
fMh>JlDFm>=K;D<I_29D?8KX\ljoO6191<3RYRNTJ[1nKm@nhDLc_DPQ[cgACpKN
NMjKcGKRfcY@bW`_KG^AkHS2Q4WB0YD>24ULj8E0O<Q@=D\e@HiGWO^^CSc>IOI4
>dlmAjMImJjg<:VOdf:1`W]6J:564<U1eVe6JBY8K?4QJjdR3_FlY?2AnBWZi;KI
V7KWn=jCnj:fN1kKi_C^6F7Lo0gKp[Pl3QZG;jf[_LoTb2eU[2j`YlRILehL8\L<
ab]PfMClVP<q`Zf]b_]8_K@e3GJIf`YUe0aJ14Idl:>@35G\L\]1@k]2[bfdZjek
\nhW9i>8[UEPSe4gjEFao5P\_4f=CG>K?b8mZ3WcL9DlEWZH`RLQ[;^``<^5c5kI
XdY_5R3NNfH5`6DK9AN71ldS9?6Hh`j1`Riag1T0L0pnSDU:XQ:1ASMflD@Hkggc
G5LGW9Jbml9SGn;\_E>9e6mKlh1fLn0GbL547i8W:T;oEjeg_nLH_jJ9VNH3i9a^
M5YV2ZT0P>3VIeGj@[bACojih3aQNl0jfaa3o`>bF>9nfjU0?LLXiAJ:5Hi`MbAi
1SMX<mmimpfR5T^g7gmFR]El2B1JD0[8Gh@82o1a=__VWhn\`EY]GoYd8P=3AN99
3aBUJSSYQ9^nd[P7HJ]o<j[imN6_1jgA6m=LA^jbh@ld@=F7n[=Fk3;Y]o2eC0Fg
<;7DSTOU2ef=1T\`bUZXeGgj]mkNdgV0]Y\Xh]FlqZ`U<U`cZYEmjIe]9SFk[aHk
L\hmL=gVcUL;c\XVB9cRAj<eb_eJ2OUASD:XPlQ41`PbVhV=jZ2SIHDM@egkYQeG
8>hi;WNfohXJ`F:E8IVM2DG5^JU_Ml6UE?;]UW^HhZd@Q0;M\FO=G=WoOg<0aTU`
?MoWb`epm;i?[PMW>9=fc:nKW`15oT]bG6><cmITDIZLLU?K[?n395M[o<hlPE2[
W]L9IRDN]:=gUBW=be\c28O6g[ONSZ;Y]a_1pK4N[KBkDc9QZSBQX?BKZF1`NYTW
TX=Nc;[_6g>Z2>8M6A[58?S8NeTMQ_DUHoiGM:lS15C@_@Q3N84Zi9DN50o\d020
i\JLa6kme;8Xo75Xi3k;Uf9<@mDLP4<RGl31RKa61cbLI^?Q@_Q[0CS?c5>RCo:;
0d7qd=?lhkB=\D<g<@N<j7R6E?deGA6neYLiLef1ba]hPCm8CN=7IGHQe]]nCmkR
e@PLjE_Yi6_XJTMG1IP=1B8PQ6]Ne8_1F_]W5G5LAUMH>=5D4]b<=cl[GHFB7LCN
:o@kdR`I\ZUBWA<@D8`XFFRQ^?aKJc4=XTqRm2hZL\eeNf:hWV^JoHVn]:T@cYD;
?NSIm;@b@X7kS3^3k0f5FG?B2:LLTe=g2LKJH28<K6XXPmYOPJg_nj5QX6Q0QMdi
=7S9fCYf41J]NIFIdXbiM3Aj_fOm?DMT1@7R16_LFFfAAdLVke6H\KW5FFV>RR^l
`q1n9:Dg<AjLjlF0ISj]7Z7E7<d:PGJl?52Bf[;_U=\@DCHD_0CEG\G4\VA^Zb[:
V4d0JNjgZ6_fI>gI5lM?nOfV;S<T0@??[kb]GX8F7>=><jL4=@E;@\ZT_P7K[^CW
X]1QIJG3Y0;6o70RagkObBD6kColf\M6pAJTNKP44\kcK2F1T0l^kL8JQA5>\bQD
[4Aq1UfgJ1Z6UXo?XnHjRiWNZ4IW?c\g?;M9V9:UI1=_o2c^2Xc`CkBM1i0WB<7j
L?`_nGRDSZPXNFII\99jnN7Gl@F>bO7\J>PV9hf>]QJUPQPod6XR>ONc@?Y_jOW0
1B;l1GT5hHdgk=k9CbgQVD5^<8kC0;7UMbp@4aBW><9b2]Qe6>=^SDWOh]i8@fY4
;\o:JL]8V^>BSI1WcQY_W[XQTmIcjg33CC36[a5ceUZ<KP1PJBL[NWBb1>mUDW\^
3M]66XR7\J0h6\3ajN7dm2eii08]iXHE6a3@Sl162;0:_`H2k=XmGAi75hmgl_c>
OpH;@bA@JelKn1XManhVDnH?SlfnV7ePdTThUFKi9Ua6fa`GLSm1?AMlob6T8A45
9RdM0HPLBdbLIHnS5=EZ@`R@fN\A2YOF<J@<F1VKRC0>IZ4hVReMETfQlBF:Un?I
FdHZKbC\;O>dVN3D287gAO5M<3gER_O7pHmEhn?6O]PS@XM8jUKkYdlMioR<?>_k
cY]DODF;f_5:j?YS=UbL@PeSTXJo6[NZna76FVo7V9SOWNNUkSZYPS443cZj0Pn8
5VNHeD:hnXi15FZH5ND]0n\j>kgiKI8eVHMi3_KGJAVF32;BQf7;GWcknD151k6q
j]TSbP98W=T9@UD;K4:f=j7jGK05lSkNMS6O8@E<<EbJ:\h?:K`QX5bj:O3AV7M:
\P[[KQl\\6DM9@8W9:><fWmJe2]l9_XcTP=SjDfQT3Pm1>P1c9bh[99B`Fi]6g6T
jD6[_AYK5X[[B@4DIo_0HBg_OCb[6Mq6fNke2PI4GNV@g<X2@0?cRbXQ?KA7W6:b
M[V1fH3k4;?J\P0gPVV]RpEE5O]T5UbakVEP>HhXl25?[koO5:bE9S;@kD\A2nXL
PQRbSDnaW9SE1VioiH<6IN]X;n?O44Z7iD833MOHSKH<\?h0EX1Q\ddO;Yn3X>1E
d\3;b7JN7NGB8Bhd>fj=C]ETnO2ZIA;CCff?=5ZgG_QHE]4ZhYO6qW;1OldV>UV_
Rm?F`m7Lc@176<Pc7UQ2=oY;1`BeUKkd>TYkdWYJNRKTPEVWWe>>5J]CFYBh3hBQ
YD=^nEb]P?Oo4BSXk\@=ZSlScdVEXh0EX1Q\dCm<`3<W[OOLA<1c9WlK]dVoP:mi
<dVG\CC\mEoIMmCDSl8q31POo`;Te4T;49h5Cn>_f6>m^i`EKgVddZG48?kR6HZ:
OD;K456hEe`VCAo2BQ<ANjV=h6;d6@6iULgUb`lhS`0\fUbYfj=fW6o3M^d2k0jR
Llf@5laFTWnYJ\dj;E9C3@S9aVbGYHKfB7M=QOH09bO58O1E9ap7[HUPSI^8RQQ8
?0H16B=70o4<C5Hn04_W@k93>CX:NMKWcU;Lnc]@LXf:4dDRP^12WIhLYR536f29
U>oH3Ra@nIAcWFBgH9^HZF^JZRB<c26TaHNACNS[13cBBd3NJSN73RUXd]GbL2UE
k56cE;;PWEgSaUA>9qn<OklN[2VOjZOShGOCph;AiAj`^SR@8G8;E9c6K7Z[dhlX
[GUOX3F_9a[^3aZA4:QTK>0TW><dN:P?NL]\U[[;e1MM1:NCi]Mi5bCMc:henBkb
8l;;8MVn1E;]_e=HLIi5K1N9lYc`lE:HQ:iM0h<<LXmR>SE^Yd0?8P>Hd_mRoK?I
CUQqlZED2dM\2HVjBb;d?V]ZWoOYKNH:[J8@cP^T04o4RWPk]LZK3A0\<jCAB2VT
TYm8enZDj92_i:H03mi8m5]lbUJF<Y3<4C_GG;;7bc[`MnS3X=@9fY0]K`[6LXWa
bHcCl7Xk^:VfVMdPK]nFL?OcCJE[7[LhSopl8J=oAK[Q\5VJ=CnIIgaVnjiScaa3
7JF=1gQ7P7GEG1lKdOCdTOMQOCZk9hQ7@n:_ci=oY<g336VLeUUTUIcL5WPTKoZ2
b_[F]6g\Zf=P1\N0CD_iBBc6YU1]D?3^V>9l=QJ1m]=kNL^>KSLAVE\59hfinKNR
dpZmNVQS;mT5o7_=be8Xdh=hZoQ;iGEQNaGL_7?Nk9l`5fHi2DU1fl7eWJW6T>i4
UQ?mE`dAN4d_f<J9@D\RQMIPB[98kcqDOUfT42FJ:UHJXVmNYS[RkC>IMfZUoVUT
`SGR_B1Q6NH02=c_HKgb<8iNTPiblmn`G:c8ncNYaca=`I73j\I4?bdC9I>624_B
iVZdLa6N4a56ghc:=23mOTPajPQbYENLRoGMfikm3Qgi[qNj1@L5G[MC4Vb2:JQX
IEdlIc_<aqn6AJR^FQ[`EJ`Z@SO43cOHbl=C=TJQT_17:CT41aE7B7BhPIZcdKo9
YRLmgRgOYe9Jj6\njclSM`R7]H>SO_i77e]_m:ZG;Dc2jYXK_hmDDIiZWZ5jW2fd
G<M<gAg7>f@E2nm7N:XWHSggq>0MXR:4;R5WI]EE35Gi6JT@KNMP5a<D0M;A<iE;
7FSLD1X6UAgo[]jITi\>JA9?55@Xc\WS6W=gcfcX`Kj8@S`>]_<KF=]iSj0>KmA9
PCF9U[bK<^dWK@LGI][>X>dgNC3A8l1loGcW`h^qOd8766oH<b^Z`o>H6kDX91\4
ED@7@ckRf[G8fZik8IQW`GA=XZc[M]JHMVU:gQZ_i_bQ6kL;lM?:G[DYMSjC>RNj
>iX08Ab@U82bZ8BoGLXQ;6>nM4[Bkc2eYlUQg\J[_[kYLVPBBP[cX`p4M4kAh?<B
o[U_8l3UCFHBbUdNR>e]m5hZh3JW2WB>kEWX\ZGfeN287:dGo7mQjEE=;NTEl4Z8
nVJZB<Bf;lLT:bK;4fN@9<e;ga=>?a9gdnMfU357gHhbd?Y?\7=F>]SOh?K9k0TA
[cnXdpX`VVaZ62:dO6AgZk;K0b?m^CeIP\a?F[k<JkCfN7[cb0LM5=JY0g\KG\07
B_hINE>m6Y<Hfm]ENhMF]8gSJe\:QTICcK^m@CRf>=7WjjHKi>b[[loYP>?dI01e
BU=LW]G6eE]V5b=@oQJVq^C?c>I9<DUjC_bC;=_M;4`T7CKp@5PLHkXOnHC]IW\P
WoDf=^knkHTcV0TAgL9<oC<Qk0kNGhZ7[en3A]B7QBn3I3Tm:KJIZ^ib]=6l>j_^
<OgjD417>A?<U:=NOmKKT5PZn9@YBN]0`3NddTS9m]n4f4X2@dhTLkYFX8fGf]q<
5D5FS1:@T;J_Bf3^lHBba`>:o>?_26V[CJkkiTN=ibjcNm1^oAia`gAf2oF?oiDF
4TG8=5V5Pl>fmGAOgn:RU?gbl^Fmc]T;R@U1Y]AIP4[jABZnFcnU:?f8:oNeIeFj
b:dd>4Rb_Ak;oqdEmPabJW<[?C4=]B=@n6>=LVLh^4gWL1aW\W6bOoF[=bQPFMWM
Ho05K7cWX;P]gI`eA]NUJSgEPOA>bHK`eJYVZal<J^MZZp3@H<C7adOcoc^<Z7K3
`BH7Ee^Q[7gPQVlZ:Wef;;1E_m<@R3]SJb<?lAm1mO\QJJ1;VCEng@\>d<4aKjjK
aA4KbaInaKA8iaD?YlVF7N1hAf:onVf7c;E=`=RI;o:__\V]EW`JL<J:amT\SAjK
aA2L=5ZXpJ3kY\U2MOkM@?4Z1A9PT>bd_@b\;i4IM`h6``k_ZTH019Ho6M5cmTBc
J>n6i5;mIlS1:[oJn79K3^<\`H^I@FFa@n6PZPX3mI<CKi6Im]`^j[0:7obnO1W@
4G<<FOh0;G\I:jS^A]ZPk7Zf\H^I@QAW3n4qIlZf3dhR_SjBIJG:nIaL_6MIko9Z
mZmhj1IbRfIWmfRh[?oo[fFVE??gbEEA6TCGWL1bNg=boe3[:Le7Rnle<>ZEMR<=
OafNW6I9_M;XBC=VKdBmRjaIQ?b3bBGO;j>89=MQ>n]mH6gm][ZoRnleUA[GeRp0
A7NeP^9`7[\LSZ<OT^O]NFh`D3;U>^H3C2gmXgd;enl6eRGYn6hQ;JYSXeYfeUne
ALQ1CZUg<l?a\EWKA_;?6Z5ONZH]?Pca<2nG955XTmG`]km[C[PjC3JSR]@E:^KL
XlVIHVB?9ZWn0HEKA_;\7^AHWqe;ZaKDDdkHLe972MY]EYX0SoAk^=@[8m?J\?gG
TGSIUqcKED5knU92JLoNU`GQLfG5:If66WoaMISk`bl?P5Y>PlAV4982:N8]h7V6
m4S=;DRKLQN08[F0MHHB@bUWFhdi<aUUo1LShU=B`n\nDcFEk5lI8Q\W<@k^iGVG
]V[\320=oj;dG6R7_l]Yf5UWFhIX<GOhqSX015P047c\0fg[HT<XfYiS_0nD4N^9
Z\iXKeR718XE4]Y`PS4BPnPDcMT78CV_\eHdTlW?9><L4B>P\]GAk]_@[:j^D2MQ
5J^XVZcZO?loPWUi=HXOCOf9GMJgg39hh]\I^H1gMKl4Xh?k7]GAkke?lfaqGYCi
TYRaL;h2FTZ[[fSZD:l<kh1Ijl=k4LFL\66J[Fo@1RoT_CgnABQ7kPm^3c[Noe\S
`H=hGc7ER?o^dn11RI]I]F5kD2bkZ9?IkLQS@gV@m_>Hj:jCSUi=N8f@3O6WiEb`
omO<<igf]C8hdn11k?G?HSpRjPY>FWPmY9?YM9c1PRBjoc^H:G]3D>2ff?gQ5BD]
eLCV1eOV_Ibk]=L_8I5g>UL0\:BQ1PXUARMeOMhoiK?BNoff`[KkkXWCVg^Ecg1]
OTm]F1[o;dN@]:Ha>OTn2lOV\U?T7]UEa@oHGbYoiK?IMU=kWq19DGIZALQP:6mM
8qB^b;h];^P0PIc_QgjTcgnM=lY_[I=he\RN[gDm7iY0EN8_T;_ORfSG5X;[3IVY
`UY9FJGaJfiBhP0FPJi?3IJhS=`Mqk5K\lk;Z3Hk^3j8L8XKG]Qhe@<6Fl\m8F;Z
bC>GTXh<e74AVIVBSjKl^ZF:6]\hBg84[8hJDZZ3d@f9Uihb=gPDGUacS2R5fnYH
^I[XEa5_CcBiHXbTe[F[MkES^i^fpHbNJE?6o0i284<Mk>hbSbf^kmBkEUGo8mGF
KP?OlCV5OKhm;8_1YX163D17K7^254BM09IQ4R1gdJ@`LUj;]UKeigm``A=cJIW9
`MbNYL7PVV9JE;gOm:oV_IVY7d02pMLX5Mh6^j]]e^0T1MlB0OdE1;og@\XNY=@]
2Q2OjI\eG<kAcdEC0V_FkLjVjFk@hkmZHdMiYJ9O`nRUj3`76hD0Eg7B;O@[pIM@
n_QhSa94M<a?196cVUJk5@d2P6IAK?QnV<nJ2REkH0m<bSnJQmSW6B79PHOV9C7S
N2I>_>n?Sd0Em7VXH1?UCkW]@=E\;T9^;716IDAaGe]mRU>:VW@2U7\lGaM0p?4;
OMHWh7m[jJ8afhBa1>PO[CmgTGZb<=JG<VF?;emcZm`gf9U80?]IkL:EEZ;7eFQk
@_Qj@T[?b:He_WA`cmN4@9Q32aT0i_Tgc]daiWhd[Z7oY87AX]\bGJVn[0T4q6cC
W?kl;;kL@Ali:YL90`lIZ_[F\iDIS><U;]odCAm=SAhPPj6k\UG0[XSEDAK95e4X
ReW9FP0SV\fmbY`3A@Bl?B43AmbKp76HUgO3LLnZ<8Uib]<SD8jVMBLm55LKeje_
C21AaZ`AeVdYPj>LF=6>a51pabY6_4cn??=kW0O1>dn=\LQ`e<>9[>A61Vfm<5D2
M25oURoSjTfD`Cc@K;3L9UJQa0HM80E\LZB;_7NYUmQM^DW\o4O1fPFDm_?MAgM^
:=n3ZJhDb7@g47PpJY00@mR5blH\`PcGjInNE^aM[Tj=DWQ:E=m>2dm=R?1P_i3g
J<j8FW[:\:EmHcS?Jg0:[NJ0J1h4>Fe:jT_lCZheT6aT]44KhnX?fA7=7P459cJ:
kLc50:>q<ZjT<FXZ`kDBfHXd^6Zg1B]SHERQn5h=UjjP4DNPmI_odD6lC5CSi^Jk
Rb<WFT@N<cDTBF2ii^Win^Q]G0SJ7^nhUXqJJA\LGj=7[=XVeAo^?CWcG9cCQ6=_
diZN`XP@DNHZ\BRXS[nRGZ;;N4DV0=^1h3fO6\a_V7mZ?=2TmYn5O\8o3LA3WR^A
VEajDaETcW7P>SbMReTXGSU1L^_B?^TmhLq<mogb?5H5<h5fMWUN7dZ<P60Yb:T0
Sj6;@4dFO>2j_]K5Pg=6SVHV]\b9AjSHJ>i^2\KT`okZ2h4?^@SAWhCFHlm\3?KN
H;T>gD?05TBmUK89Q^?f4@MBfC<JX9hhUJqH3a\FNO2eN\V`C<;ljGlh:Y]Q6p=T
Y7iJDBYQf;17nkJ?;S_j6G<Bc5kDCd?P8KES71S?ji]3?K^dTOEdBC;Jcd5U?NPn
27Cl[GH`fY2cJ@0_?@lMH:7ASCmeaq=WP=:Z^0P^4aEF;T?3;T[?bc1oc=Q9\^1X
CoiT]D^0`N>THP0MRYIF26c>jljFR[DEHDZ9lH4l4>]df@`<UT]]46oPhdb@C=3T
\Z0jc];HOLKUX\]Em@d<1E`g`7UU>pSmWk9`Akg<GY111fe5e[;_h^gA>h^?iG_H
2nASlS2C2J_M=E:gko:gR7:fiKkBC]?NEKOH4:i9Go@WcH`Jf1L1cZ8^3]i2PeHP
o@[SP0QFD=>b5e?]QAenAT[N@`NS`q\8N>:l;DdQ0c[OZD]lAKd?1iAA5Y^PfnJP
M;;T_mKkYT>\CW\FMVOeRD6LX?jJ`c8UT1A1OG7h0Oa04bmdlih1dm9OY>c3IqS]
DNHA`XF838TESW5@?hnK005[P^0?P[=9jDO6hV0XUcAPanb<GiB;da[_M<<dB7SW
gi@KNB82J2<eTWkQ^cJl_PKJlbnn9JJoP5;[PP`>=l3^3j0nD;M44qcYbk9YRIF3
1D3lTRX\K8fO3^_3b[6B^8ZOZ1eJAnm;IZ^QDaV4ABVm1R]<Z;kn\GcAcbSM53OQ
6IWYlNb0VGe?oYLGU5CZRME44ajmoE<ZF17oNAlJQF_1Tpa1VSS0K]jLcm>49bBa
QD;f36AkOV]b0aEm78jcTj]87QH[HKNX43Nhl`0Y6m1Saja56]9]^?JY[W8Th?N6
5F0Yc[[7q=_<@5Vk;LJd\T7qm1e8ZmpJma`J:i$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FACS1S(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;

//Function Block
`protected
<[Rh_SQH5DT^<8]HNJUI:TCi>UlQR?V0qOEJSae?;\ij1aBojX7eo;cOUPfNLR\_
[6:Yb8K8FcThFVfh>iYj:3QYe2?@PnjU3_mep>clgM\8eLbDEnlKCc@5KY_8[AD\
_8HAWeP77CJ=Rfe;a2RRp^]C?i2qL80aEnq_3T?@hAGe^lnLF0_3AOo^T1Ejh\X@
7:q2BfS@bBCYT]K6;:=mcnhNEAhifWfNXCpZ_ZW:7pZ54F0Gj7j89<bllZFmj0L8
]n074FdZTXIR;^A0bPmDXI3a=[FJGH>]`ABn4hqOXRe_dpX0Z_Ebn\eESQ]F:WoE
FO^SPYB3=aMBhq3GS5_7k[JZZnl:V=Zk:Nf3n4eAY7MUJHa`hEq;0nCD7`gk5>N4
?dabjMdD>RSh;gAncH7a0eQ:X:fM>F0n_HMSdN26eK32OJ8p>mTI]61LhA:m5iRe
M:gc9C0d5U3IUB<p[TVR?7q06ABP=^=dVABOe[`YjeBTPdEeX;^AE5So;@b@`qoK
IMJI4<WYBQFE_M]\6_M;e_eH98bMTc5GHoplM;AaJh[:aOPnWg6MmbpSYjMH1qNA
d3P6a4JQa`QhUk6M7D_<>dWb6Fl6[[B[WQXNp<Y=SEPUV=B8FBF9DWS_5g<l;;2M
n45EH`A51p;ZTWC;>p`PRbYaq?SfJK]FjPOFhYfg31F6FGGQm6IbB3IHL]XXSM3m
bFd>dKUDGf@ga[J0f1n0EU>a\=^7@H^1>]aJ3Qgk@@F2T6]^ZEcm:3LedhEZUPZ2
<S80_A=:_UeN?<AR`bM01O5lZYaO2:4D7gEaJ@6pVRY\K?Wd[L8\<O:_@e1P1GfL
jfIUQc1>_5CaUV?ek00a7]]=[Cl23EKaZKfj]QG8YS4]DJCdgX>nM7?F7\0med8K
cW7ck>]MOh^KN0K38jf3[5>Of=Bjg:iHilfj@9<e;gKEcaPWa;6KOHqHg8?1HRME
:dZEeQGb<TG9AM3^T_aRkfQL>i]1@oH5Hf<[f8\?i1IQ5BE;=g3Og8;V@=C3G5bR
HmhXEalT<nbmK2EmA\gKEhiT<ZNTU;58I`4V]g^M]6_c_EeDjgiTiWD_k75QMU?4
i]1EQqD8kMW4:alQg4WNT:KDS1o?C6f2TRCHa?Zkc3HHXXoe_<GB6@24:UH8IW1C
>geXP[]XPKGVbDH>Q1C<dTORE7^H:_gJ0`D`QRLUQbCNE;FAnbPgG>^]3NBgj33f
>IeBLCL\SSFU=P:[JJU<q>S16^`M<<<jlZ1E9:=6@FNPLoJQ;\b9O\eERVIRbfBn
b[l2p[D6o8VWioj7JomkkcH9`\AC5S_MBl7PT7NTV4>>M:bb]g7kNfgJXa8C2;Ze
GkDBE_\BeZTCLM2HTl2:GXbf5c3EcdciihF22deXQSg;nB=UHUM>Nj>8o[IUUdge
RIDJ3DS4XldVmIVXR^Xqh`G^gH6]YO_fd@@17ClgSB^`U?84lLED3MSXY<nkE@k`
cXH1[E0R?3@7bdZm4>a<ZiO=b>mNi0V7NmVXM@UM<n7W;HY@l=9EBf[TNZlf;CP@
0A^aKKW73VQ>^[Z94?n@1m6UN@]SneK6k?qFbEk4B75ncHKo7SR@<Bn?g8>O:WL`
MTDC<`KibB9<iYfKE5A?TOe5GP7SDCOcZHHUBiR<LAZ]1O@P^ne?ghf0Pb0XbN_H
bXmFln=NLWMn7\4>0VfKckBg8e2EEC6fZDLk?;Nnb4>[HPf@6q1[X\>73R>MXfnU
45>RRSEgAS[`d5aeU<5cm;]13>_?U;5>6U5eka0eb2S[RoZ`o:16Q5]Nkmd7>?Dn
j33`Fjh\gFMbnTD=4Zi5dVK[14HmUOf:^JULH>@7InKaR?>CUCi1Nl0R\6V4@gM:
pfU52NGHa[KDkZU6kaoYbCfdWIRB]N;Ing;Bo40Z\gAk[9l0D8A5FP0Mf;YR[FP<
NQ:\k1Rmm<f<fP^aX4mQZ>:nndeCiPjGqadRd9>?IK9:4g0<4T^NY7M=lS8^<b0L
WdUC9U6>EhdMblkgO9V06F;51XQ;IaXKCIh[L<N;3[_3MPIQW8c0RFPRL4VcjM?U
i1jlS]iQ_i46<2[PGiKImN@KLcAWQH<;aOSHg?]JR1I<:1h6djMD1T[bPO<q35;9
2Ag;[b7b4HCZACe9i4ehPAG;YRE8\f_CgM?D`W[:48B50HaQIXf2j2WIR>ENT?JB
G04^30AGNJk=jU:IXU52Z[iGVZh@Cn_nmPKjOU_4i0_nbOFoO<XU5D1h<=:T^n^R
6SCJZVM3B]WnKnac;YS;G0p:EM1ilD`cbCIZiU^S6deo9I?Efl9Fmip__kcc3<ON
^d0dK2@nj`]<nQS4i9j>FZ]lH1Z?k9WPm?nOCG<]1i49?Oni>S<laDXGAcTIkSQN
BHF_]HlOX]@a\JkRJ^?T\5>XW1Vib@h_KIQlTXY=RHniRNMjScPf]]mIk656[Aei
61^?_]QW5;NC1D]3dqHYZm@RDiYWUCS_eTKLW?nHdDoe>T1U[If^h8<:^aYRAY5N
=eo8ZELl`cP<FiJ]lXj6_;ambZE[WnBlIHPe7]oKWJ@U]CFa5hA9][Co0`??>AS6
ld[O<M@bgA3NCaRcf>:fNS[;=67K@=YoMiQJ9Gg@Xd:CqO^ZFFmAI8J@aMnn5U:?
XY2TV_f^J3RERna9bf0n@:@GPfDAQQPZT_E4J;6b]CLgkblf5jCZBkoifH>l8i\S
C@[L6Y\aR2K<em^F<C\;KQYo<E9DL?9T=0Y3K^9]FZ==m[3Q\^>M:MQ;FI=N5>FG
[O`oCjYq1Z;BWg@NSIcfnPOQMg2E\G7kOaISWU`OBRZ9Vn22RG]in1F7>Z^BI3XZ
DOPG0[ZBcNO9nQC7mnTbl@\=W727^SQ[SNk6b8fI0k;RN^eNA>NIGU0]3lRU58S>
f8GMDN2LZ\>?cEHnGbNUmWnRRYj<Q]\nbRqE8_fo;jB1^=UOlde]E8Pbe3[]J5=G
eAeKJbb6URR3Eh7:E]9Zh3ePUQ`QTXZH;PWlkPn5MPP_3TSRX@3iVFhKkkD3\15U
QI5Z^F4Y]YgS?9W[JKh>kdj2TfjiSKO=m`n@ocH6IJV_<lIJZ^2f[HN@`>KKdqSY
5DN^6iIN4MUQQ4meGIo51mjmqH6E<i;\48hd_>R8J\I=kTlf_8aCAHm=@IQCSJh[
B[mFgDOOc>jBZPNm>W?i3X\>odRYF::>N5N>caY0i`2aO`64XkQAh=?4N74bioc0
d6YoegK94TG1MNBGfj00cQRQee?Q_U4B6^:SAdVaC1A?QW1eU1=qm?KE6eD]hW_c
\5E_TLDQ;SH[J_jEnJDB5DkE^==Zg?3DR5Xk[05=Q=h]ckONbhL^Hhl:XgWh]BP8
mGZB[iaiSFmMGJ0]9=:?8]ngNTWDZ<2^FcnhMPBOSM5oCHZ2^a]cjA1SS\7TQa9a
nA_WG@?[01kEJBp51<K5XWo4]>eE<lYf<e6<F`k4=;`GTdoZRoUglNgD3KOVV:bn
H8lmeFPH[C[TL`1OJ8\blHKcWnl@UX^@I0bf4XfKjf]Y1gDUWoUA3NngbRHS36H9
m7mTGTaaj`;0045m2FJfFX1bCQSS^U:VWGJd>aUL6qUaN]ifF;R]AP`fHP7]lncR
5Mj[OqOHE]Lo3BebP`5eM6U=7eebJmUYSb69^kiI9M@3HD9]PLgGhi3SnnO;JVWA
LYP^`iKokWnSm1T8gc8dkNgN^f5:dPKnW8o>Gj<i9b_b`fe=JJHi=>?a9EW5m33c
\b_dLiA`J1k6bY[Z?[9TQ0eCTXm<kV87q5emWI`J;4g9SHBQBT]HmEhJ02LA^?\F
UL@`JL81<YRLPF5Ao@moSaC23?JQ7RlC<HXOe_jV@TYm0Xa`Tmi^eKf:5kMNVB<F
F`CHn\F@NR8Z<YkTgZ_P^b\S>=d16h=S7?i8bC5>ia7kGgXY]]W[gd7L\l=qVDmM
jiNUAmoTF84D9c?kD7a1:FB;hgA>Mbj:1aNOj@2A<8_aDfl8?`Z_aB8F^4GJG@WA
1P25cHXMSO6BJCmC<78g7jX_CATnVZj@GNL3Wf]lS838>`Y:0bO3dg@^eVAj=]ah
HEPfOWO[i]QAK24F7Ao\:5pD[SdmmKo6?fDcoZ[6U^BAa6?0L^:<C[0O4hR8D2\o
M[n?IhXLb1LW_@4EkJOB6kAPId1@Q=fY\=57ET]<Ng0Oa04a<e3`J<k<Rh3Ff>;^
X?`_A3:Kj3c?[o2h2?M2ff]FFd^AjBRYK40m\eG\=IZ<ZQI4Ep<GHak@T@P[>b@c
?IKdZUNeME<mkoZb:aSJ8p`^cWbZ]i4n@g4FBX;?8U:QBPO>dCSkKUFR^BBEfWXl
5dmjc=0W9B<69kAleZgCM2f^CdSZ_@Z[\E3Yj`=G@DDQP1do8hUIJ?2n^c^I4kJa
6nbiOB\@>_LS9nNI5EN36I<_F;iGUWeffOZ[bKFRa@`@L27]qfe[YoQN>Vf]8\D1
8P1>?N?Sn2liTT2mNM]OU3M@J4e_kTEWRDWGF8XGl?9`QQf]IHZ[e^]emanVd<mn
IcoDIR?QIF?[f7Nd:SAO:ZJYGc3a4lhR>D5=gKKh6l^G20l;CPNk[G\Wmcj=?dWi
=PZkf]bK;P5p1gXNlY<X?N=kBA_1>b<dO>ZOFdb1;kD<71_[j6]ae;ahZl;eaH3C
CM<^g0;K6mDhW9;JYI[g]Va`HJ]]<DERU8;aqmQjULc]aoEU:35SL?Cl]IlcC<mO
[VDMB;9^`XoRBU^h<Ilfe^?kYMWB[L@Z?X1_bI=4`SBaD0AAUX2IX:2lLbo2OXmo
TKb^^]CI@?VS=M>XPbm:b:gXGah^\WZYEO4O5mP=DJa4hNJWP^Qe?1nn]<P\hMFk
QJSpE=VY4^[m>0`3MnSf6THH2EoQSJq6Q2NQN5ZQ2Vc2:X@MH[b6l^OV;lc?JMb<
?ET4HMgW;6;fDD7>2JmdJK]emLcODKMI=XaAj04Xc@G[oQ>HGQR9HJD[mBK]0H3Y
iQJ3U7P31ViAS1UQcGJcCko0elID>_^6cJ43UE=e17S@G6DI9adjG:;`alcdPqWC
Q@5P[E<GXjWECVGb]N]L\f4SPhPe54l2<McfT9g2i2V50T3]X:lnQR:nR9o2=5fD
8KJ3a8\RF_B=ikW43cQ?Q;baWF[NXVSATiHT9Ji^>]WD9AGXUO^[^o86Hn]\0aWE
]R3O3l;`?KL3=J^NUBoQAWo][d7NqZ8Y^7m[DF>^jZQb>Tfjg<_7BU^l@noWMfPa
3ZaMX`0`?mf4hIFUkWk`I_nEm<91_5A=9Zf19UQ9DhYdNW5mc`S73Y4oEg8oYV8E
X5F]fJG>bGeVhiNj=RNoYRPjdYm@`Z5TPbkBU_I;8D6=LWofTG<o8NfAhmgpm7Z>
ZTTWHY[SQfmH?0I]7Lc<9n]cOHC1;40YXa`OhIGBY60_YWbmhIa547\8nXZTd>XX
657XYmN^di\F8SePnc8m36_bfK\ET?jUbQ`5OZNTn1hDTUa;Ia1J8H2o^[<km_0G
`_@_=37@WV_?S0h3B@4f`Y6@??p1m_]W@kYRKTPEVWWjA>>J]CF:b>lhDECe5G[K
gMW9VX7=0<m`fY`;;hdCo2=DMDCT2c4HjOVnh:9\jk33JW_^J1Klbfjh_^f88dNE
`MU]6F6ZConfJRVIgbMdBQ@0Zf114@5UikHA<2hg=T=@1@9bU4?gB>OWJp^AaDY0
Xd0Un>C>EiMWCXBY[B=jbTYMZZRk;:PXi4Z?XAY3_hSk<WlmP2c9TfO1IeGTA[7^
dOS;S8E97P:<Zlc\:Ljoo_[A=eX;26?;En\m:LY=YI\5KMlO`\\YT3oUEA^lV2=V
hlYe\PhZXiJOK_<<`26YNI7Sp_UEFc@R4filX4Cl688FeN0O:[WB1A6M6kCX_Jc@
>[h^ceNWHcNC;;L0j``j?jBP?a1l2RYa`TONmG<HeSiQgL[PFm=C9EC5dDh2>82H
^:K7oGn8dj_Egi`bLZKIJJRgj_^CP[enci7aMl_lF1NDX`?L]eHdb\=pkH1kj^LL
>ddUH;bf^\?8;KXe8JYVdKeP=1Gm_:P:71MVZiNTPk0chOiMo<L3cJTC7SWa=^I]
iZ7S]2D^:e0fP?=i]o;X5GHXHdfDn90UVBlk5aleJIf\3Vcm]QRm>\O7kKKHm1`L
>^O8gBaZ\klH@:QPoo5H@6q`eHb781;<R14kB:`jYhb_lD?Zl=^?DEjSI21>FCh@
dnCdW>8QoJ`]d3;ZOSaUWc:Y;VETd^PDmd:`KKYFYcPK0nhJ@M6J<`[dG:omPIYV
6meJV]\2UeE:@NkKDOcGWH2`P4f5lf@RTmRhj2fd0YMXO5;hB=ng1p<bYBhY1S5Z
7hF?1fKfh2kd4H0KHm_P7FjOWfYg`p?IlLD=EA7ijjbhaP<_3KXS5PHVd?3B3QQ4
f9:0e^:F_9o`90ceEaM>AZ_l2VXLF3mkKA0Y?6AF894V2]jZRPk?V076CVAQS2l@
ITiEbjjM@l@oWTh3<YIVSUfo3Xn^lS?DkABPBKVa:RRZl]g58dP\^C<<V@ahqSQ5
GgW<jY][Li3EATLeS4?;He88lWQcobY=db;@]XoCMF6Y>@8EJ7ZAg7L\mHbcXRg6
?m@;[7E`B\I]Sg8<]T]lfO[V9YKc0Vb5V@QBAj3MRb_O=S[^RUA_JK;\FM4[FSm;
Lc3F[5]aA=@leXFXgAUYn952eU7pb>5?9E2lf60W6VkN2I@h?;?36diQ^CXS@`40
>QU5Co<81X^UK:BIa<Kj8SQoaOO7RR1a`<9V[QPmXk3PfPDM2aYBhLDNboh4Sj8h
\:;BNC<\3:Ieh4:fYNdm`=jaSb05b6<=kYik`ak:C5\?HPnj3AeF2Z`[omp@G`5G
Cc^OfF<6[LYQ^R?f72J0]b?<jgRIL:2MmSRio<GgSMjJ:n:ihjj=2em3IhR=7:mG
:g79CY;`9?6]GCWiKnjgTcBPA]eSVlWbU;3]JKD1`A@gYKj=80cNSn>j<EC@Lobn
h8a8U1?6>fXMflk5je=9L5\VXqXJPCGj4H7<NXW9WP<hG\@jdVNB2MKX_n_;:=ZV
Ze8V3<:aJ4GKoe8B8M0Uo\`]kSPfd9OhPUl7:6E\g55h5faI6;dB`o`TA0AHnEGk
5f\SPVZfJ:U7j_c1jgd=U@AMaAXh4W2ULjIfXS@jjU3Se`oWIClG3@ShqMIjX@f=
Gl;X5HD0aRNJA=S0`6=5WNL<>XBkm3hQZbiE>[a_XDbB5\O>4L9fP:EWlmR__2gZ
3^R1HiW]oiRN6<8kV;@bdFCG?<feM00fIWjLAaZeFcW:hS2Yi]35@[;j3MaGoRNX
=ijD^4?7Re<7[L@E`4`?>KYqLm[fgYb?_6fE]V5<kZ3GIS2EdGjI[@Em74iS>]iI
>UNY@iK9^?HHYI\cMMQ?7Yn_iY;Nb3L>SU:<l=8GPXoUVCHGWSgUp1VFJ<m;U2o=
=c[A`_=Y<[UdPP<N\0NiTePWTkZV>K_o:on>7>f1gc5[HFj;h`F`faBVUWVAEPS8
m[RA][7T=T9S0IZmOdjhPR[]1J9YYS6e;YNZ[5@e^Jf;?CN;enV[5aZ1PjZn<?JJ
MdOqn>cB;Oa1kWmAEWbMd<B[`N7TM=<n\Y3Cm]Z7AC<oPe83D=fZknYa;NZLAnUa
4j]NYMFk9iIXBeM]@:RF969OQO0X<bWAF`HlWd@5hQW21Vi3R\U[ZYH[1_^LhPU@
fhF0GLb[ZP^1d?b7OWqRU\;HLGFhJc:Mb5Ql<Wi[\^le7I45a32DQKORUZE:c<i>
PqBXLIX;DJEh<1I[?0XcWYWIZ?l5OjEBcd`=EP^L=i>m8^<7gdK[U\<S6IOV85MU
e_cUN>jN>fNHEVD;YCKFGe0B@^3GWWRmPCaWg]LjR2^oI68[fH3EiA>>JQdK8YMk
fND?n4]VJIT7Cf`hqWMRN5K]^DBj=[0J]6:iGlEZ710TJg7]5l61a]PkHMmOZNac
cF9M1eEgmI[38kMego`TDTn03JD]\nW72Kd864YUm<`ULU]9D2l<X:4?XA1IfJZ]
Q9?\>j@Nf9c3U^5fmcKEoWZ=LAPoQbDp]cBOTP:\0]Kjj\SJia@Man9<A5[L9cnX
<F6:Nod9>_nZa9@n<P6ih:ibA_Y0hVcLNHaSiBdJ?Xh\Dcj;KH0G6:nRZ[67l_Cg
?CXD5eB_j9L^D:jfaD`kEgO_LfYbhU>i@McMIX5cML5n2=p\D7bbZ3>9ff8^6:J;
AgLLd1[F@U`1_UciHDSMU1OC`0So;hG8LP0>`VJRLPfEZOF3_jcLYDY2MHJJoRmP
bVY1bOhfa6f9WMI?ekMbW_1]>ShQ=?kLM?53oUPNaPFFbg;`jgVAf1A:\c0L:q6F
cKf<\_`lN7;996JFU0?O@[k;T^GS<F]\DN8QfC`GR]ac?`<Yja8JK79=<jQU5J<M
IQl6T:27QjTeL2:_QOom4T_f1i<H6J7aX96L5d4U?F;gSBB6^h`XB<QF<n@;_XDM
:D<fnXLQTUThp4?E;^Q0_Nf35cWBVEoTeeW3e1=@PVZkQIgj3BI1UhDJB6hU^88G
<H6Rk70Op4fhaJDXVIR=1@@UiCJUIZM4MS>ZQLc0`:36BSoi4D7]UDP6l2A0Qg1F
^;5?SDCbajTlR[9<T:S>Fc0]R<`DLSQkR>XZ^Ij;[D;`G9iIFFIl;i>?1C0QS;g]
baC?3nf0=ZS]XaL]Q<PmdKhpcooO4;d:D@?U1gA4[3Y1ZS0LJPbcdfjoCH9o59?H
RmC=?6iDVVbXb]F20l:MaDFY5oC3kn:?PPIe?aa8bDmYO6gXmB?BG@3pjSHbAHnJ
\VC?;acM1Limn>Q6KcWYPHUS<gT`6KdGJ>GP@8KIM>27<4h@UDHNY]fejH3@N[^j
Y:>W@5@]<`dkZ;ZOWcXUKUU:TheMCcjR<TG>>GcaOZ0m<4DCTgfMoon;d9Q>IBh:
:CnP@5@]m4`Sh5pc=M<SBKK:@CPd2?4a>FF:a9P5^TY:E_jP[lQ2`9m2glI<F4Y5
<g9Uo_]UH[HgPm^c^bH_PhQkESmlkSdlUK4dF<hN^?T2Z_lE]i0XlAC]\>60moj:
IhOUodkd0X8mC0fGDiZmR>FP30]lkSd7f@K31p4a^l[iMP2FS4g7XiV0C2SBQXZY
K<OARnBTfTH=0jQeUd=mOYcheVOkJ30;6[CDTa4[=bT3g\K]_[S_L?J0MkE4\=9B
1KiGRA::NgX8LlOoLF@S_Ih_8<O22Ffl03:L\^mfUL2D\Oc7cWS_L?1?hDQhpYj1
\miQ__4edE=FkG30OOILOH;VoGj;CiKfb7QVA@MaDQS@9=<864`_Hf3`bKeV4YCC
9;V?C@a^eYVH6RPd5<EiGZW5?>K;LG0<XS\o;9[YjnGk?3=cJ4D`Unl3[\Cg=WeP
;?b@bj1nIYVH64SST`EqNT\F9nTEIkh0l7Bjf@LnG8hB4WF0=Fd6Lj7@Q6[AcViK
XJ16DJo8`MXE6G>jMSH;NY`:6>ILOZDR^\^RLWOSf4`V2W?O7bd\\0RUW^TRFHOZ
cWg@\jK3`]HCC]O`H<9aTC3PQc7DHcCM^\^R4<Oc8Jq^YV0<6gKT5ZPP=;1Y^0HP
LOY4n>iccdnaWS9n:Yqdb0lDEFDgolhSVcBM[0elc2gYe5AW49gRA5UkP17R19PT
^[51cAANT3[CSn31F^ddXNSSP1d`2WBiKeLRcfSk7Q@:GKfY>9jibfa:gK[9jKXj
9d1EY`MN>]A\ce\@JC:lJMCmnj[:SNQiKeLWQj5fop=7CS23PeHVUFD\[9eWm6P=
=MFQ[5DX`;4L]CV08:`6LRaJobJoYCZ4Y=lUjkg^g7=8NSlPi7KAKGTkWeX?A2gn
0>fQe]BY`I8j9OcC;T1LSl6>MgVZd1Zg]U<Tkg7K<J]\SCTk0fBQLBTkWeoEdRB7
p@5;3G4\A<@l:AhoJa=L[E<_S6nD:gRX52M:7CL3;m`Th5dD7o:gnGGTUfSb4aRL
=@?G\C5eN@7CJ3E4JT3M^Te0[7n1gCOXj6RMWibIObDb?=ILZNiZHGTXTCk6Jld:
B]\dW21lc^5_G3E4JEcEREkqW8En^ZbZ`iglHl=1_nm4cN3koR2n^F^0idIHCkJL
mbg8A?oLTBNk5j9i[LJIn@3FW^@1R8IK<8GSD9o2b^C>klq_a`TN@L<hMJ1gV4le
=_HUF>8TKEmYU`K:O9i^E@B?@]8b0=4UCD?A1I_]6EHTKVB_gb2;Q4FR7P>6804\
bKPG6[?_=SZb_eVncjFfEOQReAhSUj?ieDYGgDpgmU?Y9JZ;HJ\5Dc>XVDZlBMP;
QkZ^ZP2<EG0GRC;bYUWU3<d0W7b7cBj2^]i=SBRg[f^e=X0ebc2X=NSdSN?IgDBK
@P7cA1C=;5C`o;On62:T5MQ^l`H6PKpIbhAFYjm;T7Yo:Zb]G6H[6c:_i<Pggf_h
0Ugak9K9lXB>L2JSTDdajcVnci^?:S8IiomYKX=N9PP_ImPR:Pj9Whpe?KRFkJOP
]\1U<M;FPko5AfY^dAV[[BRKX0nXS[[Gffp\cKK=lf0Qh1EPTUV?fO?1a6W6P3Oj
HDCMU=cP`nam]=l:1O:R<nQL^:?ME4GfjY;\n^R:Fe@aG563fYJf0dEZnh79M02A
W^fb]m:Qe[@d5LJ>2lB;oUj>bhp:7ajdbEKm8>WBn@3<4e4VS@ZS1Dm;BK2j@fRX
FXciBRVoJJ8KjA\9hSZB5[2fQVm:Y>ZSXb[<BB2iP[@BPE;8\0W\0E^T1^YDbNnf
oXj@:a\Ro[j8NE<B]0pTo1OBKK[6GdcV2SL;YAR^@8;NAP>m[BcZ_T1j:VTo:\2N
kTNoda@lN^@[UJ:Y2[:TBi>87MOgPHb:8da1kTe_3`p_^@FfeN01]AmJP934Hm;c
HblMnQg7a`>gY4hJbTP?ghdB?B7]0`l;A0k2C[nWCdC_FPJ:V[f<6U19T?nBi@D=
LmOYI=WJ7P[\O0^QLg7_mUeKYKcDno_e?^q`0M;W4@f^^aeIg0_R41Y428KHhWRN
i<ql1C\5]mkXlF;^CgAo@YkX\>ml?VoaH^jU;bJg\F8nkP3AaMMgJFF>1:H?BMRS
<nWlYTLVaJ5[o@Of^g2NOOf=g0>3iI_AZmkM\7E2B3?k<0]GI]OGg;ZTdbqP>WPF
O3PiLC0Qh4@\^cH9PDR>\AnK^C1bRMk`e\<NblB\@;EcXDg16\Q\]\DlhfPPCjhZ
2ZUW:]1Xc3<?\\gX]DJk5p0l_ibAfjiFIE7BHd49MNl[m^PiKAI\O:h^Km4ijd2^
6WR;29Ck^M3U6CT6ZKjL;c0FMG_o:2EQS^MfgWNKVB`G9nK1KB;kNE\BL?5=NQYj
XD:Ung_PbC273qZ>485fV8iDZ[5L0VF0L>;e[@lISj=VQS>E=2@L;Tkm=II_dS1n
H1K^[K6ibUIZ>@Z^lFI`^g@bCbKijgI]K[FRBO`fLF@_lMFnA[0cBbPhj6aPk@f>
G_=5lpTF33TlI10F0o^dPPLn5Bag<GYLcL>h5K4jJ=c3T7UYo1PoPDc;C_jP[=VZ
J3ACWPT_4DIKTnT\YSB3;?[?OhfX>peXA_CM;hO6PH]=AS``<7ikJaDP[41X:YgH
FSTcLhlk\o5Rj^cQ]XYC6odP^]ah?7e[Dd3[gTY[mCWDBM_E?VmD4ZEfG\B3kW0>
XOiO2HFijbJ\M=5XhNdlHq2nm]iP?QkHAhQKdO6j5W]K:>mQON<\[Lk7HP^:Wf@4
=06<0[5gOS9E?WLZZEHoRn2K55gLETQBZ;oe^WecDfmB@QaSc`^AZ<7abZIb?1o_
TlW6U2K6ImJBJq][N@^e4278\EcD^hgj_mSB7b_Yoai>ULf1cWn5kTiMXfXNRAUc
=Y>HbCY@C9WB<P]2AgGNIhToYoM^<J^je3J2Dp^=QN9m?g94E2cmCmg5S0o4=_fQ
;cogL^39\a^DUE@oLe:0]]jk^[83QIl=U;?Vn:aI`3QcTepWFl3Bnei;KLM1CJbN
3B3WG3lR2_ljBHI=;@BhJ8JAYEX1Dm`ZOFBHF`GmHkD7jg7WUa6AjM8G]4NVBaJ9
XZ:=XTFoo?E1gO@jJo70_GBTnWC@A6jj14ciE2qNc815KW=g`IMEU;M?\VG[b?^K
?CQ[NP:R>7fUg?ecfIJYd>]HhTdP_;b_jCfJKWSNEDYVN5NBFYK8bAEYV]hnIjAh
aPRAVY4^bj9\GB8jASX542\TSm;Q_9qSW4_c5\V7EMe9M`N29?cmKMgeRS5GEndc
j^liYNj5<hGRj_k0?;Ve1`iO3dQL_2DS`\?0ZdhVVQ2em?:BN>j]RkehPpZXIZ:a
pXk;WIF7$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FACS2(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;

//Function Block
`protected
AHQJ:SQd5DT^<43:TQ1_L>JD3Un6<o6i]P\FmC\FTS3j;Ipg:cTg5?goeYXl\Y4S
?8SE9E@bdlMTiQ3=4]]ZRL[_^<VgPdfl]NZLSRYpg=OICKFhkgk4RTk[ahH^i4nF
[^U_TVJWLWm9a^8]OPW4]BS7klPJee6cpHW;a2TpE8B2?>p_LSnW3:Jc8B8;Mbj^
k7O<N:Y1oDeHX[ig7c=:LoVm=Og6Ycf34l:m]kg0jp2gD9=@q05E:5PLPMo\2\ME
ohLG6U=@PL811c\`q@M6GM[Ph4kgHJ93M`bKjKB8Q2h`e_oKLL]OSp]Uo71?kGGj
Ef1BZX22JDlSeoFX]lGF:p=>mHX1q7kWfGeZZY51D9e48Q8cZ>6p:o:6Kg]O5j?k
Z8EnmEGS1QA<FiI?a:J]B394qC7fW]_A=MgkCejOaF<Q?kl@S@a5]BoMBT?`lKmp
VML[LBpCcnULL<RPg9B[Bo88kiS>V=@Jh`Gk0:n6`oDWokJa9WkNO@phL_C6VYaH
<3Z^f2VceB6T05OK@T02Lib;Z6\qM]5G\m\X6?SUoSdgD]3Q<2M>`4<0:@kmAmgI
UXq[7iMFaqG@\Kk;RUVE7KfA5LOAJn4GAKX>4V:VeC25mUp3:3deSo[lJ7ijkaPH
YH0]>cGNmDC:ZWqQ^Zc6n2g=gJh[?FJVbhFl90eWgi51;mq=U]WB[Jq5]:5Y4qaI
aj02JJK56fP_YDQ0j:cd4Ma1W;]26Xo>gJ62@Nj^2XT3OQM1MOhYG8XRMBYCHLfP
A@J=oPo<MA:XgJjnRi53ElZ?ddOV2VoY2i4bm^>fPeFGMC^aO132K:4:Me<RaKNT
LW_:K8:nJOgMp\n;<LBd8=YOH8OYmX\GH3Eo2bCHXagjS1X\ln;fclVO9l1a:Z;I
;?Boi\5=kG=DQ>HT1XW9e`VKFMPMC\gdhcL6[_9YOd:hX[c3@KMiE[^Z^@:<;L@2
`ClXXZc=c09W7_>iN:kOU1SXSjWqTkkY`W=9be1jB`BZC_6065Egj0@2n1aS?KIS
T4\;YFB8d7]5>?gMM<[nhaA?HLSY25Gh=b?>Hh4\V5Rm@Sd_B\Fc:nfI5gTG>FZI
i;Q;iF9YWgM<X?P;99hcBPA\G@:SALLcFQbFR;;?8kqE_?k4M\NA35ZcUnA2L2T<
m9Dkh_jnZ7==`bN46?TRUaoh4kET>2Z?dbf9O@E:CNOn:UJSjDPj65GeG00JgK<`
9X=;d0K?6cg<1447FA=b5FMN89EnJchJ]F2U:@jI@kT6[oT_5l;Q:2PETqhV_ki0
IQ`UMngLm[ik7A``[OFobOJFZb6?Wk]aAF_ikd_gePWibdA;ikEMX`3]XYce6EC<
DSYZi]K]<3l]IWGZ]B?i1N62NPiBU]5g<4Q_UO<=nYDh2F31H;;6X:GG00JC:6N5
iX;j_8OMq6_?kEakCK0SniCcJdE2c0nCDcE97MAmM6IT0i>hi_i29VZid?L7afdG
d?Y\[SEpF3P:;OBc`@M;[f25IkRagGEB83O<eK4]5L2hWj23GWbm6kIDD[dG^>n2
\DKJQBFGFXicGfB@\_Oib@ce<nfiW6PmJ`?US:bO9KMk5Ma4bJbO:J2Ph@j\`\[6
kDKh=lImg?EeE]jeHIM@k1qU@e9h;iQJ2U_0C7cDnNlgFN45llU1<WR[^:?@3f;W
?E4V\]EZ6bbdEdZk@a8?8:=Hg]^<lcTSGZ1jE[ZmhkF>I`l^lfQb55INBDM1Kb8=
^K1^bMO?5>jjII_5>adh;\OGI>WE68ZZF<i\Jp=>e4kE^:OWA>aL20Gm50llFPj6
MU30nSEYS\>=WcCFIe;?_c5CkAl1gG41A^QR\K=mD^[XlK_BP]EnmAf8310DOPQE
=Q9D>R`Ud_nKHfeOIAEO<>SgK7nfjA3jA6Y]Yd>7[gMAeY>PoFj9pfVdOmX_nNaM
YbWGkHB0PAY74BmeOhaeamS1enhd_JOWV67[^1ST?`1bB@e`LSe@NLNl<Q9Q12Nd
Sc;I=5:IVmA^c`K4R[YKpGa6aR5mAhc_NgR?VN<iomG?[1kUOGMmlk2X[IegRO\m
Za;[=__d9YP6216fa=aB2KCX75T4Ynl;L2FE^]=:P8=L]_46A:d;7dCXb9AXn4@`
Z]Sl>0D2gN6:OSA2KN4Ok1dKf7\8QB1DSJmZK;fK61i1dNDqaLY4?3DBlXgS9WU6
9g>eeU0?IcP9C=Hn0SGISEbdd]518C?<H>6P5LTM65<UmKbU9Jm]78MC@l^`=VBE
Xh1V6On:Z:aWm]XZ4iffAcHL2HcZ[Z73okU4ck]2SlJ2aIKVjVQRP=fZTdZ9TJ^h
dFBnLdEefBq6=@LaOQ[H705gGiDfODDUF]@?nWA5=aVc8[KiTXKnn9i8REEiD`@9
IKod6jJfHJg3ESK5EaQYAnG5AoNXodG70S54UakR\0RYY7gL5:PXa=a=XD_??cQ1
1[H1]UPMZ9acLPOi`[<VcGLk3AQ4jc\LM`L4Yq4nVK3L_4DENWN8G4\;];@H0=7a
W0FicgkGA8OcP7mAd?BXM?@G`07hPFmVOngXaZnKK6J9J@a0JECiR6:ZQH_WbKCR
?AnS?ji2Aa5XTni<_l:<m6kj6L=Dkm?N5jbLlP25>B\N2BPoflX?YB[6GZ9H_`GH
q6fGa;WPjZ]lO^lVj0==dZNI6cLn?NPT5CDYeXJc7n8TBh4a^?<h;q316AjROAM7
mNb:MhTa:55_9D8;:1eD\LDkE6Z7Q7Pk?QRJ[dAGdAZQ6i;D7:7KkB4gY[QLUHdi
k]XLeF>D4L`_UFlBI71>07d8EIW@H]cTE4T>[`Y=ZSfZXP08Ydn]T5>BV5M`EU[G
O@?I_<4kkFnk:YSnqTL^V5I`I8bm42[HeGL:kA_<EjO4dEZlg;2^oL2C98Djn8=C
j5ACk@\PXeZ`iQ1fF5V[BNCm<lWajN_BBFXNc@_:VV^gg1hiMd1^4o<m;^WVc;Zf
JiVW_6T4=fiXBS540\0?nI>F7jZlD1dA8;eL3BSEZH1p27?B5B[JhmLT;lUKfCQO
6JI?d=IYdLbM56P\51B0Ccl0_Y:oiH:XmQ8J;1m0o\4:^SM8PWFlK3VSJiWRgNC]
MJbI0bVP_PYB4gPOJmIfo[92NTI]4mN4<W^`]Wf\dRU3LZl];2bV0>E9Cjcf8E=o
7Cn09op>_;=TXQ55bU\P88`XdemROli8SELSg0`_`F@VP50H5Po1_>X5X?6kefA;
6:km4CcabOV^kBR4`SWlSMMd=4P\ObOVnBl?iSIk`FC8Q90?9AlD0\caD\U>[=P:
Ra;dLcL3Pc;;EkTWn]eFFS`Lj;Em]XeZ1pED@``mWH6gfhHJeRU:R6NmS9I8L^lC
PkaLOPe\kUkHGonH7ZTNEhORJm>ICUC8NM>;=5cYjL0NCKCFM<N7bdFD>kK;D<[V
\@<lO_m8jLOE[WMXg`XfZ63KmF3BoSa062kYDnU[bUU>aN8V2:b1l@867ik5pUf:
OGcSg2c@OQU>N\H;giW[YCSM50[VL9VBOL8g\BgU<lEIBmX48AD^KI5_g]Mg=hgU
G;BUeODBTMdYCg\_DBg<>3_=:@[I<Bb3QUR`FF0KcUgP8C[HRUGMT3OP7?\WN\jO
EDA3VJRhP9o;WY?bdfj22mVqfUQ3[iTAifLCaAmGT[;Y:h:YZ8N795@2:TcOR_Eo
[oJ07NT6m@ePiKSEX;:FX9dS0>COfR9WFOT90k_2M7P]D8<IgK6h1[d:JbamRL;@
UZSRJiPaNK8U3[fBU5LiDP>lliKL2a;0bKFTSUL`6OZlW@9I;RqgBhAiXBnPR`A_
;?SNm3KWZXCQS6e>hX8nla6MmVi4GbQgYLZd4k^<iKCBLe]Ak0J?@]=L[G1RI=EN
63g^^_ODU=CoOfec?73lAaTBo3Fd58ClFeX]HWg:Jam^4`EOVWo4?PCmnc?EFD]2
>c6V\FaKG`lh5q6nUQHmA4dmhoiC?7T5\36Y[@Pc>E_j=ED45<TIZEUA;Gkk38ag
K5ZCcG\K4Pn^m3RE^Ee0OE5Xn[7SB]KNPLi^bd><LDF1T2?EO2_BC8;1S7Zh3kDc
fLo11NGM5kIPH^6<>RaWL9E<WO6RAgbYZ;KKQE4\FcGjpjoc>DYMHXCE=3G;al`>
0Y2WNRW5D@SG@AFlJR68Q]\KoZ1p^3J[kYLWn0b1^?@fJfdkV9I[S4S@mZlCAl29
<cQ^nO7=f]HWl9@T1JQdC7bTK@nN9Y80e6On<aE8n25]UT@E`86E5WA0_L1Ji_PR
GlECT@5LY8le5;H74c21g^5hRCDT^i=8L^o0;JGGb844h;bh>E]1DR<_b?q[i]M>
VD[3nRBkhc2W?h5jGL4_j@>=cRTAEF:I>VOl8Y?RQV4>R^8a3=jWSm[hm<[k2^li
hK`e7[FWmMNf35Pg<S\lm\hh2XDUTjJT1O3ISKQL7LZQhYjjNU0cj^X]@b4[EH]B
@58SSP<=L>cg5<YB=R[E8H@kRp\o1H@4<WK<boPS=k\M?_mVooMU_KgEb`BbY<AB
ih@OBFb<H\mMEBT6=c37SHNIGYATEDPZ0WNdbllJdmlA30VE09XEd20lP`BgM;gi
Fo]J58A10_1j]\3QU8Ff5oJ;bM\0G=?jC[aPaTS9oUK[MhIRC4\=[CGlpY1WFl>]
B]^G;0l1QinAOQX_[N=W0590f9l>RhRd1lT:QS`<jk@jLee6Vb^Nk>=S]nYd=G2N
l?UVf3bJk76:2foll:^_Dq:ggRP2AObDMPik52kniM=14Ym3Nh1N=Jh]K`7gZ>WQ
>?E5b5Vmq^DSLkW0B?@Y9amHc>Ll^eVocD0g_Yh3R7a?[0LhWI\bP>ZO`Ia5dig5
_=a@SLk:=h`o_Cjn4G\mI2mEGFWKD^HX8nWQU?2A\Bj_L>5VkINHJ]000i_?8lHL
:DNT_SEj9^<BDT2Ai2O0gkn8G^=7aHBEJYf8i>kp@98V^FVj]bYLCX_JUZ=V7@=@
X`Ek\VEgMKI[Qj2:5Ub^>?XjOZjTWlHk2F7FYaj_]VYUHNUQTX>Gg1TEh?=H\YYc
C5egZ:6fHjCRBZO4^FR>QLS_VeZZPmR`>`K>l17U@N9YGLgU0nf7RF1mY=;GW?`l
OgXGWoq\Xd2=Y\i`4n3SgmFbP[7:>KE3gjI]_Cm@YNUfEMc4jhQhN_CgO2oj643`
;01M<Cok<7KnFSdeUTlm4U3fd\Bd:S]HI9[2Yh68SQCS<hY@Ij@7D;X=9i]`FIb4
i>H^C01\6FjVQC1ghi5DeSl7__L8VP4VXiS9Iq`F1VXC`E4[]5b7AYMbi29>:af[
XlKkQh=cDTWP_C2DnK`eA=i9UR2OIRNKMl50LY]_T=3RSlcC?[g@L:MlTbbXSW]4
D72l_7Ab@>7g]>d0P8;`H2>S3ZOiPT588JhA`O`FDN4_0WWBQDSe9IWoZhG46OIo
_<QdqnnbjBhbMoOnRb6QacDA4W39`1[J]BFWk\=?WkYS=PC;W44B<IXRNaniAZgl
2aGZe?C:8E13@`=5de>BR>`;[<KBj;[f8\SY`UgTR5JD:4OD>@1?dLoi6CN7Lo6K
iSnjRn5KFNA;1KJeFcLSYB]j4oTXAodUB6^p_J_h\U:J0_nVBFaeOgR[M0mW>jn>
LLCBG7Oa0N;LUOBO;7lVO=8h<?SMgG<jqmBHR^IV\hf4Iak<T]ChTPSHmR^`Be9@
;K4h[i3XRVE7B73E[hCibf5jET5OF?AV80Na0e8=jOa\eGF1m5NX\D7nomZLZ20m
_JQ;oAcb`7dKDo08nM<4EWY>QBX;b0YYOmifn5fHbTM1P=<RQ7Q4X@nT1@gfFknq
PMTbg8>Y8M`MYW0D^TQfVXnGULjFJ?4]neD0RL=X`d``KTe]MR3[SE4@HKZT_knC
[UnVMORVlWTYQ8A4ccVm\]GFR7f8OQ3iCL6N>>?<iUe@<\2^ggAA_15KT8A\GhM7
P`:m[Hj1NLoHHL9NA>Zihnmgo^0kN[qcC@oZjSW1GgUBiO@N5d?fMK:7WljOTK^]
ZdH38Ob;F8jSiNg8k=eDD1_olObPIn6f5IH1i7BNJ<0F;Q^8]@\L=\H6NIaIY6^R
0ICG47h?3GMKjW[fKJD\]kCJ`1HG7Sbc@o;OSO;GMUYZ90[mm@CV82\5D;`nRqma
Z[<aCXCb:abLZnVgEo0J6bDOKFEYm>I3\dpI4O[fY\O:NIcK]`P]V8083kC:6_=N
c579h\i_iViY;8TLMYea6jl3h^9mMHe9T9i9QB4J1ojZ`U2lA=f8SGD[o66Aeej5
Q3AalAa`WY@C3Ko;H<GchkiFPYIeX@nd4n\I9ZmBBoTi>Ti`2P4na5KP]H<9_3VO
?pKk`HD5`kj5WWV=R0S7iOFW=@D<6n4\DoMj[1=2X8g\@FVJ16<Q@3=5Fa?`dRL]
m>W^cW[PL<QQnEoOmI`mVQ^Og@YklGZjTG7H;AI>b[K723AkgHj[2O2^GLZ<JX>Y
WjKhQGL@k>P86946UQDCg\gnBjM=R06[pVhEieI4HIRQ\UN^c5:UgTfkEjgAnKLO
mI<d<@Oa;^`;d1=9i\a2YoFMhTkH:<lMdT\U]g`iG7g:hbONm1<W;[D4j3h]4O6g
giZ;MagG^jl_MMTofY_NfXjfN5`3]P7mMV3_4A<jlGB3LciTRH:I_7]3;V:3Ll;q
5ij[:O7bUJ3b`mm<d:Y=N10KeE]Q2[lMmnn:VgA2@nL5`d4DF:GSVmaqo[]90^<Z
93^dfCD?KP0NR?@ScZlTIQR:aH]2Q6lTF=Vh[omZghi>USB2Oc`l:32n`Ffo0:Pf
AeY9JKlH`P5_O>`o_OCO>j8ZjB?kIK_R487RFJC`mDFINdo^jlDoO5e_o_d]7]8k
YGARWF1TO9]:FYI?nIX1nnqhD@UnLX@Vg4diW[YjkMd^19`<VOWO8@P<gKH765NR
5nYc`6^56lVoWkaH:<8dh78Pa@P8o42R95Z4jlW38^`M8\ePmZo3:f0TMC9VTh`k
:IGUSl0FZ>VUNR7U=FUGAlmh085oG@V7\H?mbM7G_X9^?VeCoW_eIq<oNYC1o\J\
MlMN22C@27m>B=Sjo\iYWGD\h^\>[3MVM9b_n:`UBlY5]fSo3A;8<M_LB<f>1<SB
cicXiPhVmC6Z44Nb43=;Bm3BMP3l41e1nEoAbi;l]^=la8a2fM0G3e<VAe1D=RUM
OjggPC4H]IO_0QDS:cKmpfJ7Xd876oQj<hYn;\>W^Fh8ak@g5debnAlNo]SMU_Ff
QKDfoNbA6XT9Y<5B7dkfcUBoAOGV:hjc7e]B;DW9Wf`U1iP1WLgN5nU@^UMQfPU0
5g41=f_LZiRkD1Hh<b05NfCN1aE\@N5KfeJI?O?5O_[jQRW6G_JqdBaQORembPSa
6WWMQAa1G9f4hS]g14?5KjYj78S<S;KJm7QE6g_ENUV<pOMhjT_^6D6Kkf;YaR9o
MY]HUR5gJh7Y[<]2MQoT91f:bZCQJbZ_:QYV0`<YXM9@ZCUV1XTGXHC\^<ZD95g:
6IKC=@bfGjYn3N2:R<KiXf\92^L0:0kU]j3^6:0YBW0;3OhIBCJHXQ]834\l4U[f
d82@P3@ieQ9pk3ZQgC:1PCk84PI\UPTg@jGR3?PVljjVBj>[CJ3EG7?QleaokUQc
\SEJ8H\0NmNMAD`6>]jZGIf_jdHmgCD9@6o^n[PSqLmG5R`:l]>MUoD=C[V<ZY?l
WETnA8439RgI::QkQNT6JK4nVmHRo[_1_gT]]78DfaL38;OMRWZiR=^cEeFCG]mS
06HFbeMY``]GXCHIkf9`K^3]<]DG7^K]_@N]:j[]5\X;Wbjhlj\n1=2pOEYjSWXX
XjibP]=1?BX4?h0?3SQLk6P9Ri0q1C_JJOTSQTCHIXVn;GC0:_7Zkcd7RCXh0ceb
eDm_:`79Q^]><L\UYim?ZNfQ@i^i[<HAT^Eo7>NNR;BNLBfMNU\hh6mP9Y`MH9S;
Uh^YU3YL]9<[ml_5eL\P80f2@Z5]cPVaRcbn5C:S<mpZRcFIX6hDXN_hgJT4]1aE
Mj<cg6A;g?Fh]6==bo9e@U3KWMD3ER0bVEAPjb8Q7YPFJY\FC3D8Q\T`dlhKj5W4
95omPU_o6OTGn;JTMhSDn9aIW`GbmHToO24jCb4X85DmYFK3?=9]3>=ACqc5TKd3
^ZlZo1Y4mAiE\Wn9McA;9FOWRci>m1AU13nNRY9=DT5Qm9>PaUbU8_eV5jbYQNE[
[fH35^X15Ea36kmEhQ4IN[><SCSHZkj\Xj>k9EQZbcLEOW[oL2V388e8XNlAoNM0
b^M[Yll<pj0iLRZJ<5Z^K>;aZU[i^M_gh@W\F<A8ejE6PX?0Tin;BKShm;9UfdOC
OJ^?N>`cofIhH=eYb9HcHfHaXM4m=][\AQN>:S\oYOA3h5^lh9TCa3LQ_DnjY@K]
7<l?DO^G0K?mmcVjR3^VPWXqlF;0YfVk_LS@X\<]L=Z_7k;Dklp4oNCcUY5X;`46
58_SGgCOBiLl;RY2C7U`D7FUVnLIc_LWgNR4^A9g<TN76jf8<BP9i>lkDld9^Fa>
@nIZK8f1n25<<eDH]>@`LXCbDEWBWV`7U<O[97]G0GH7WjIoP:C4MoOHPi\gO<JK
6q6Xl4^?MVOdT;1?H8QWlQ9E5;Z`Da5d8akNCjZ]S\kEY?TfZjhTUi[hN[RFe6JN
mQG56RR8WPP?c5EXbhXFXA;BB<QXGi5EneNS;kBSl66SJ?UdF9^jeVJ<V[1Ce9B<
ncM61;[E@NiDAi8Op>_;=TNC`5627P88`^`eTE=l=8Shc`gBL4`F[VPL0b5b]kaL
D@fCIFWF[aFj<K>kVZ2M4cEPTo@oSeFYg`5D<:hl0VN@72LSCGk99DjhY?@Ah]R@
V>b43iidC2RjHFY7K^bG?2]d]L`Ed\dqJjMY6fKbiW^M<Z]V9O8GXX4YZdq^R\K3
KL?7X[d8JO5<LgnK\OYHE>>>SnIEN:0JD[U6fHQ[E4VDWQD>G8Q2Z=j6QAJBI<Xg
J4dgTC;:72`OT7S7ig0i7c[go?qTcJF?FHmM69T5lRfToSo1jcV1dB8foeAVTEkB
LjacFTUMhfCDD:;9<SAC5lglhC[TThUEHdm4WE[KEi_2DV`@BkjHGQkYIeDL`nGR
RcbnRUB]C_N1T?C9C_\lnmdUgn^5e5j>`gi^[e6KEi_eSLT0>paBVW0KB9Fh[;<8
Ca^\[>9LkB=ZKX<QjTNNgLiYOfKLFiDF75nB631210fUlKQPQja[RkXfTCS@@Gcd
Dc:]^kfK68oH2>DkjS0N?Ii<;A6g^P=`3]>m4I1W1JGeAZY:\MKGNb`U35UT?7cd
DcL[hiP`qgOZUU6h1Od[>MFJE7O\RCG@k9WY8^7BL\0KENd>j\LQ`4b>RK>E5Y;D
mfk=mCgdeg2emBi83=n[FklRF=f2D1LJCmW4Z_BBDI]DTeFQM;TW3\>^DfRAPYl?
=AC?3\Znd>e1o4K@a14i1klRF;UUmHHqJ2J3PjXXH^:LHbZH=Q>ma61cEAc6W73H
Ph`VXBhN0`8;A@jQ<[b=0PnU[GM8^hkKJeXCjEDHXc\e>bShj7C=O`C_MA4L=j3n
IUL^HF?0Zo]K=kSmiL:e0M7:XT66[[aMkU05_a8<j@=o>bShhN7dk`q6ho^?hgG_
O5QU7G?NjoZkGjm1XkVXnF][]j[@a?Jjl8V7W\NgRQpTaR91VJi:A642C6o6ig7V
hZ8j19=BdDdV4_jLlcjk9hQ9Gn8nbD_oEH9QfE\be_BT9h055SC<DK[`D_0Ic]dB
7k2C1jPANDkhoN]bZQ^>X6ee>7dleS2oE=]3_De2FSj8V;jehhB2nCI`D_0a9W>f
Bq]b6ed=\NS=?0\_g[OEH4lgiEDTWThHV?TTN1k30adgDhFQ9dnkb<K0?3]>;;KS
2o]bDP@Gc9`]3JcP:H]VGI<Nf4ZT]]>OV6A1I2\13HIML98k^P0gLUKH^WGOj@b>
Cd8Io;>Q3mkjQFcP:HiN=CN=qhhd6VehAFDU`KLRSh8BB^JPPa2a<^F[I@OWTDjG
YcG20hj>k5k81S7njm8hWbQNJhcI6TkI;8ZPDFX4G3YXFjg3BnhECA`[JKM@YD2o
[ceKHO\7Hm6DYS`_LSDa8W=kJQk7MN_a3gFd8FX4Gl`WH:^qDZR]8LRPI:=o^:LC
N:Y3jV8MLJIi>gWIRcEOBRZP23Vn^;jS9>oO??<IPKiXP<1^D5TWR8AQ0EojU;n3
JU\jTid=jQhgEdW\hbfV4lXJicY5<L5fT=TO?<^@kXW7kXl1ZobkVA`;1@7iU;n3
Zh5MYhpaZCNbPMMgo=@5e78f[7:h\RYfEB@NTcOFm[7cQGR>lm4doAUV3CQeCKj9
FEclNTDaW8nJnRNM=>>GI]aiH9X@hq<QXeC>WMZP6ThYF8m=GAJ<S5C@cOVFGLIh
6Ail7lJ\IofnILkRYN]hRd_^9Fg`baQBAN\5PMl_TJ<]_ioBBK\O[:cAakb9>6m1
7d>UIGd>VD:Yf4^B@8DH@3E34;@V^q5\9:@?ke^\Rk4[9pcTg<X7abEMdCM^8fUC
9bVU40\bW6gijiQjGX5B;\]6bQh_hGH=AA674L201iM4T_e\WkhNjF7>dh^AKfc;
j`2d]1`fWGXK?MeL;`Hn?SLd9J1kZGGE8DF]TM1IE7CnPqjg84CVaF93<Z:OH8>j
:8Pe9e1VD:nENT1dkoJCWToQT_17=SEVeX0j8n_gKalZAN8KA0@<\h1KiG1XCYc@
N_UZX;]FjAlF8qNKYTQhUQAkBkH5a4HLgg6I981JA3S7]:A<kEn\W\>B:<5:=`=Z
0Eh5X8RKgk>QJ<VD`lGG:l<@?6_67K971AT4A9;I>OKb?YaS?B\Q1nk5^9afk\J0
JIE?9[B1YIX\TpC_53EFj9RE:dk46fF=DXl?NLWV>[[3eDF97QCLOe1MR3b\eTMC
740@OHZbI\b<_XLZMF19ObQSf?GB^^_HJE0^PDZUK5fN6KGUGEBAA@KRXLKMYJ5R
f42WTP0iY:FOTpS8`fKbJ\`E1V=NG8IJ=Q48ci;d4mJO;9cSPXCJ8`RQT2dIXA<Q
S13:_>gkc`6WC1d0cHb8\Zch2^KP7X6U0QGOS=hP0>oekpHXOW8?ASa8?]]8:R]_
iN;P=aA_WKI4i?m>@n6Pa>XdGVYXj9X7`_i_1<[2><;44MH55YYfJ?73f\2;7THE
4higM>JI8Ka7NZ=e@]H0^>NQAg6i=Wnf9S;3dpKo^3@m518[;:QL7^oVTQF>KL9a
OEONiC?B@5DTMgP1Q\Z8jLPG01GUnW5f8\B5X6K50Rn8bcAO>:<;a3SOFjNJDOI<
ighI2Ec`CoGPWnjFQdfUgc;8R3ZH2pD]FFU`mW=6?eEhE10A^O0YfEJ_ICP66\n`
LkOF=g=FK6gSNLeQReD6ejmG[`X5eiD7LCXM41f94:bnkf`;6nb7=];Aq:GX9\F1
b^Q8dII4n5ohBKOInIj>7cH[\dR6VhM42fHc1^UPSJbSRdHoXoPMTnm9\2o7lVaC
KTa8j2@SjnRFE0L1I``:cWD]j_gh6Oh0eY\aL2V>KcK_X88MInWcSRkVp^E5_OAd
kA`GX9Fnc=dfeO^Mqe^VC=R;PG_L;gXeR9>8<i0JKgJO:CFRGd\d^PH>S_lma>5o
K`3S5dKGMNa=jZcFb1E:@a\XE^?LTZ4GQCA`X[\Jh6l[V44gN?Q_jSJ_n[@P45JZ
I;mW0NK[2S;Qi`WHq3:@fjd<WZ1dhL9fbZ4;7iDW8fZcU?d7[J@jQTOLcG^4:LUN
o1:^EjYfZLeX7\_m1`AJW9Y8KUCdebZ_IFEo892e[0oBk0^2pG_A9F3fIoBK;0JK
[Pb<]N_2cm6480M]LmW?;2B1V7^I7XS:7HRWIUH^Ngfo51_Whc;L]`mHYB=KafRf
hkC15<2;78iVdek=Afn<FHO@CHXVgJ3^hB`1NR8f6B6ldeC8qCFPMHonend`@\8_
H?XEjOnfOh^P3EO@dGG`M_3HPKn=@n]=VUB:VlB:?ZM502UBo[2d:kn8iRc`1GOV
o:O7Wk<]eG4?9A?5<SJoogj@dld5P?Uh9DS_I:\Q]bTV2AIJqC^9dK];T=]ViUYW
M2Gg7Le8a8cdbf:5_KW36Q\L5?2IJm5Wl;nOZk20oa[fJOohq117bDWL1WnKmaJL
[;85FU]a9Gn[j0YM[lMWSKILgbG:@XDkXefHBLh9W1LHQ\0@@8n?3W6mk9YKigDl
8aAedPPn:N[TBY^Bq\lH4\V0n813KL5RQUO>=7P00G]_YT`<iNEJ6MUldRObNWkl
c9M?0BkoZHP[_bXYJ\I>DlXjonlb`6ZXgOBe^MFlc[:]dkMNkP5d^g8F<fic_aKK
0dYP_L\PpAPRDG]TcgdgVDB6^L3^NeWei:7Q=YID=RW4ImUV]?Cd<l2kBH@PJ0T3
WcKiYO:MRA@IA>hTFONFNRDfBQkL@C^BXkLE>Qdn1J\bk281Ua@?;7Pk8SDg\Wob
qTRbccUl@?>ScH;LDW?:Z<KCTnPI0RmES7WYfRcKI;5JmgfZ[D`fbB]cnCCh<lHI
LTnVL01XNV3h:FSVGJ5WgKWD\nPqc]?\K<paL2nQ:J$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FACS2P(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;

//Function Block
`protected
gS^7WSQH5DT^<cMRZAUV<>2XT`OXk89KE^IX`?TLM0[a5dVK@Bf\CZJ9F^9pRX@d
>j6=0gc8YKcR_jkU>=[W_ZEKC\HEC04^CXU?2icpHV=@nX5DT]><X2;SVKRSN0L3
ZodT2a_^Z:<\LAn3d\KCE>\fI8p2bVBJTq]ImI2TqDf1Ba0^eJ=nZ@HN1lIJQa>\
=gSCQeZ6TWn2BQAJdfjcc]9kA:e5@cNCXL1p\c5LZ8F[16lYllm@7]?367>VTQ4N
OjbXa0QSX_`OeCSPcHCMb36Q@HO`jd=V10RjpmL7Dd^q1K<hJ<11Sj]1nOoFMPF_
fUOPYWW>c7AqKJ?M9^A\XTMJNMQ?og75k81iP3jVhG@\4;Ybqh>c2LhAP:k1@UC_
X6n@4oeg]acf@a<7q=bo1@8d7H2ZJQdU?_OFIFW0Nim01Z13hHUH5h[CN\mqX@4c
6:q2UDR[Z7OokI?SJALQ1>?Y?]g95LE@=bVICGSpFH_1?\La4CM>b`:7KGodbohk
5nb7Rg?m7@G]1JqUfg6Zb21I8:=T1p[l1GXlq5k=Clk=aF[VHZKkk807;T0>S?]8
B<b`B\7R9q058n9YJ@8F7Snl90om?b0TEMH2C?^LNW56RDK^q\86D4bF<35o5KJ_
pNAIb6XqPN5m>TIg[a6l?;CV;`3Cji7G=AGbZZopbl6SW`^O=:>VdV3GALgg9RiQ
b30k2o1p^oBhf5YpPC<NKVqYc3nP1:]<g4S]7fD93?BTD>95LlM<2@5Ya0IE1`Tg
a29W:HPT1kdGa97qE1CgQ[=KG]PTE>NfQ@>[fCWUOR1mMi8Rb``UP>[7M`O:OhUP
]LjR9nWKVKK3g5MHoZXULBCdAO70_fGOVlm0B7l301J0OTN5aPXXPJ\ZL>n;7db0
A_QJa7enPPK8NX<g[Z_SdI162@Fg`XpXcQccYbg?<Ajmb<dcmeWWJ;:7Ah7^AfHO
S\N>eVTRL\NH2jTNh]7C@D8S`Zg4?94TSQZ2>Wnm8EQ^;gSdmheK;C:[[:84_>j3
bhO]eN?1b6Bi?niK52eON`oeeZhEid4BFgTF:J597?;>9p6WAEUoc@`j0n5PO9[_
=keVkAUNl`JUPe2SEY7<j5:FTaULBGJo`dHlnalXn^PD5EhjOho@R=9PmIcl]>1@
l2F9<WSVF8[<AC?7^lUWm04>mX^Ja_kDj4_:::lln6e9c7HkDl4N=JC_E^07qhHP
jMU=8Tic5eICoJ2NH?3f6O8kJ<kgOCakIP0>[4_@51ifiFaWdjhUMQOjCOiOWXHW
N821n_WQJ6?>If2nG?5:[DT6k<@OQhcHUdlVjOO1JgGd0]G_jHOIF5jja^_nk2Nb
8P<MWN5`GDcpV@?3mAcLW0OYCnm4;GP8\84ZKjgo43S;HU:=j5fofi`Xl6O[=Q1N
7F_E0V;DiQ1e3<;jMFMA?0I_?DA3oG1JliI<2Rf94NZODZLWDjb4E<8L[]1A2IKg
;IUkoQ;9<CQT[FW6ZNZ?BPFiQJpYF=GgQ78Anb@Ll^5\C]GfkdAR2T8NE=^Q9Zln
QUWfiaiQ]ifa?R<Q;3CBe;?;__SU]e3P[^Kf^CmAc<;@CiW];YCPicJ=gEEGCO9b
_>XCgJUad@R_BiA4b6Ia;;mR:;mN5]Q]?IA];^9@3qO7iQee]L;a=108Y\2ZHKlP
PCSkKaf8kjfHYl;l5Hin25H6EQ41NNOPZeYPbDdo=L\U[a?Fnm5^kN@75Y8Z>VX6
oSg\MKj?bc8D4HBjKWU<l=f@^BBK?kgceh29bj8[H_:MecGdRb\QGce9qj6PIK9P
lG[a`OOb1:e[3Lg9j2bgU7c<PG\5VW1V172P2NMHaUb<FqR1F@d_Ll1ah2c=Z5d^
E^V;e[3;TAmnYjki86NO7>kKGWc7Xj<3M`HN<bEAZ=>mOjnicUiiI;6iR?@7VD=^
nN=dK^_AhOmn43IbF26P>AfmMEU12X2g`SY>[><KZZbXkVNgekg^O`^Ck4<<q8Gb
;Aceeke?g;[>9f;7EE`U]BP:R9NRNDd5\:TZ@Q<FaYn2QKfU]bISbk1lnV[3AbMm
o^3FO1:EN5PIDI;fdR\l58J>R<Ocq]TmJT_lVeFDIk:S5:M\O=fMGJP1<kgMDPAM
ABO`9]e<Go?j42O3]^Bl6Yo=<<dDO=FAm4No73`[PREc`AaHF@;X[2cAl0R1nD@o
]6C`aMi:WXG?R]eA5O9@<2gIj1aL<]Nlgo<E;K4\Fm6`;R>^mT1EoICZW[?pBm5S
N<5kJd>OdUPC2DgU>915=3bTK^9JdM\4I4]R2W[F_EGXaHSVDBD2OHCng2UmlS3Z
jmU4C?o3h@o2d2R@c\5CJlfdSFjSDX53bP1S`Q;=^[N=RHK=`P=^]:;_I]koB;WI
M`>3<>cQY_K0^@a8UW^?M]65e0q@<XT3GOG4JGh`B<=YQRkYMGjem0`=ZJ>;d=Nk
2<@fJdU:WYf2M3453TAjgNhR[<Y9A142J>cK7CD[lGMi:nKA>`DA[BhK]o9DE:K4
nTcU58_[7_k6\2oQ_;BEAlM52OO@a\2;2WJlYi^JG:Roa:e_H9K=iXHL9qoX5\?f
JTRYU_9Mo\eaMUG_^k=ciLfEj0`;cV1eVWobA\UY6_L\iWCi9<oUh@TKn891\P2Q
9QFU1m8I0DH1aAPLZdT][T]C2_P>@RP;<6\52YOF<JEWHA]61i^2fM;=ITo?VVmc
n:A@8b4jn8QX4X68;]4dLjWnqDoKL8n]W\F_ZfaTJHF94OETNaJE2dT=hQ<O;M_Y
V0@Z;L7`Y7l[JUNlk>lZCc738`]lO:@o3p^gAeKo`<@Y4Yi`J>5=cADTO9H4faMY
F8WZ8SUJD=OR]TG7k5cjI6ONM<b<^j\0CNeBYeFVbY6dOT<iZBSDLN5V^Q5]0`ZF
l:Z=BRi=Lc@D:mV^ggfj>`A=`TS2:FG8@S^1`bJNjP26fC^GLEcU0D[B?M1>c=LV
pT>e:mKJFnV;1WM56QQgX_`jSIj6ad2>@PVPO02O;4lmDhbIb\69\AblMRL2>dc8
Il3:OKh1@e1g57XIROK^V<`_EjbL69^bH@4]:HNC\MDJYYIlMn4WP[CdFXT;S\d\
<TmBAlnn6_FV\;j849Y0iQIL>4FN3VjqKF5?SbYkk024Y;H\dKMnW7\dSUjiK?7J
;SXAY=;<i=JiZb1PS>5jHQGKP40\oV0o<dk@Z=J\PZ]3ngOO^Y=TMd340dIJO6X[
2e>U6;47_:Tfh\aBJH^^@Nnjc3PD5fOXKlNT2HP1<7CY=jh1Yb<VYU_^fVF4;mpE
2^]S3Z^KZ9`^n6ih\n@l1Ob>?O3L64_Ql`\FUmf?EE7DV5YAXDh^GFe9O4Z;?VSZ
2_C6IjaOULMHfJhW2A=e6J468lBkaRXeRK?=Qdd1\hAk`ke@gO2iC]2EQOEdUd9E
_6fDLOIVSMM\MYLBE@E3YY1[_OhV6qY52_T>2?QRgd5:WL\bm;VEEX6Bd82U0J6D
PDVnY5N9nZHH[kdWVSEN12PMa]\NheK<iCfPh>4n^k>l0JMjiin`BM_>S3]gihNT
O;K[@_`1]Z=P?T5;m44KBjNUk6Q[9JYbbeHMfAYEk[j1Q[k0HXWhH8aSbYJ6qKll
70OlWao]lnG7A@L7]47_D2EkJdBDDV=ICCmRag6TF=coiaJgFYOa780LXeXCXcO4
0d0Wb2WHCj[IkH3?iX?fDoECQ]VQmoFFYIAji0bKbjm\SRP?TmIOK68iDPlOHKIB
J>6nA9^\_<TQn09lWaCmUlW2]@6p0OiQjOKPU?_F542Ka^>Ve_c5JcHQ31R:kUZD
M>[dR=egWHiO<l[Q6nihUcg3EenC2VaQ4lLal[<0J3A5HJZVZo@lMAOg2^fS`:bQ
PALh2nN@5hG32L1\D9VGSM67j=GV0FVS;0m<PoaDPlhAbDJgRi?\H_Ail=qc^V`V
19:3LOHoFF3[HcGY=P>@1q3PUlk;b\F9_R^VFLfeXb@X4V6QE[PJU03UJZjjUJnA
Z6UVMi4b\74ndK5m23j`lZ8aJGD7UjeBnWAgSZc`cO]de\6ESVkaN;Q>m1[4UKLT
2docKE^jjBgK[=ecA1RS2a3Q=7PY]U8N\2;WF41e=io352HYWlJ`q0QZ0`_Z`@WT
g]5:21UY@`AD6c^fH\7@6I80=b`dPY>ERB\LHUnaJ>5BaYG>RRKQDcmME;BJSnPl
\Y1D9KJo?dP_UlI8Pe^H@Y=RK6UA<IAT1_eUl`Q\_XQiLG\L?m8>k0Z09MLNQ]OJ
i08[Xf8Jdb7ACkHR?2jqJ1AMM]fm]>TcIb^@:h@<KkHNPDR_i5a07Og6de_7>53A
U5OoGAl[jVX06[An4]UX`86QP0ZFCM@\[ZOCf[F]7iA[lhhDiYAnYTV0i`_l0OD:
X[d=38^V]N7^bIYQgKHLJdEWAgfbk?GLLTGFZH9O:U?QBD3fUYp?Da_H1aV:4?I\
S]@Cm=@n5]ZoTNUkFgKN\4:3^9oWf[jE]Qna_8^k:i0c`=G1FV\Gm;Eg8SL9Efn=
KMfW6kNQRJ7NZR69FLjgdQ12EZWY`U?Ig]G?Pe_O?KjT>njVTeh?8]5@U;Wak=c9
7Y8cG7^_PHda\C0cYpf7j<[EkP^kQUVd9oYUZJK^bOR?MbFW<E22HTKl:31bmeki
0EP;Z79hb<b6Um7GEIU;>IkChn;4XZ:BIlV8hVDJ;;_InY`4LLPm@==R?`N8@AaC
]__^9F9lCD8\SO[BBmf5loT:iKilfj@9<e;gKEcaPWa;4ISQpMTAaZS4KT?I=mA5
iaoKF9G1J<S2n9[\;_20qmMB@iMV1];DS?l3IUAY7JWD0nAMkJ0]59C2K4mBaH;d
E\in;WC_[NMaQZDch?jE\giYH8gd^F=de`^;^3_BZSK^ljGFHp;:9VK4BRGj2oSU
YGoRRPb]:d>2:F?aAl4IoH4B45:a2oS72jC]3XC:XS\1o@?;S:5mCH^ZEUjWaO4\
^Pi0n`I=cNAcbb6^PK^egO5TkHA]^HCm]=55\U;WF>gU?OKemK;\TL42M>ZSBVFH
5i<4SUf@>:2UL<n1p9_cb5I1VjbWE?4hW=6Xl8enHRNI8X8EkVQCW7^Wi4D6<WHj
cBV[@Ul1JeBl6kVh^EmB?mChl9MSgDQFif6]=J_jkfJ@@J[6Zh1T:DYUVC;9H0RY
;[=l>\5cfXib]O0RR9Qh0Xia0f@M\VN[TP5eJ_cfRMLOL2=pK7O^6TW3?B0WX3T`
_fl\[M3V<OK\lQYEJ]Tl6@7g0ER<5V2o]4WVHk5C9aY3klVIb9_i2D?Y\d\^CQT6
OWLh[@AZ[k:F2:IMK]_LPj<K=6FhOEnb__S]9KS@Tf7cB2[6KTQ^M7i1haOigDP:
1APSO_5>ZDkWkOqY5^j_PomfN1b@Xi3i0KomZQOa[0@_J4PXS^eSlQl6]MaX\F<7
K:T5;FjS=EYF[A628[4dcDbcS<oN`nYXB6Z8DAY1SMSTlMU8L<\\dFR;2A4\Wf3j
daCn?Rj@7GR83>1Y[Y2]1SIk93lnGO[ccO>ZDa=RVIn<lq:Oo[jCJ^6ghScZP9qg
=H2MckEkS6^mH`a7G:0CaC15J4Y:ZdE6KJ8J3LeON`hZKFB4V9X:RD0?h\3QjN][
FoI\R\[haJ1WEJBcS>e_G_m8\3R^V]AEP@]LDFXV^8iH9mFZ^7FNEkoHlJP5m45g
jN^nAK2@Kaf\WSjQ[OThQg:3TeTJhqLn_M?MXN3C8l`^WYh<g8^Me>dR=TKZ[2YR
OEao@oKOR_]?8I=PKhn?JH1_]dW2@HYe3BLF3gnHi1WCAT?dmhA^L6:O@L4`[ohS
mN323>m>fD@fcnbIC4MKKfL2\Y5_aLL=njR10H`CECPJojW@;FgCZG?IUE1Xp==O
8HJI_4=>^mA:;k_7HaNBUHk]3>EkLCA=C?I]Q@]9m\6:kke\<X<^dAFcQ9Y5IVfS
KLXPWb[V7;f[B4hIJgJRFXM1[k7Ej@>\93O?42I5nF0nbD6SjaliA8H;^_4Mk=O4
TTL5m;Q?7S2ECng<H0hA^W9S9Acp^aaMZ^aBD<G`YknoeFoVElIcWPS\f;b_>R[q
53aOECOB_k\MbO7BH=Ro\4WbC;b2\R\_UTMfSLX9T8dNH2^2:_A\OegmbaWoP<SM
U6MF`0gJ=]0@ZEQ8PTfc@NKB``G?IK1<ToVn6c=B?93c9:j2PYQke_eJ23=3`eeT
5o_J=GaYW4SKeA`?Le:V`d:>1>>nH7pNWkfDZ[`B9A`=KZ9WeI]D9PCb2SKdDj;E
;BG1IPGhE:6Q`BX\`GjEiiRmGF\PAdN^QREFXFa;;>=WlGXo`iMj=LhoRm;^WVcO
X5CVXjWWM1bhXLE5<<0[VASN4=<gW]@N`1AUXLNiSCFo>ggKUU=A8^^[11anCqWW
h:1\:Bd5Kb>96iHHdlG\NGZA1DAMNZb65n:RC2knEmd^W8PT?1`f<MVD_l^69I=2
Uni8ng`F9]GEef9Q52gY06>UQ3n^;^13FTTb0ZhSUSHfF2cX>ZHUR:T5VVhEYoWi
<24B^MnXKL8FMlP8d8f\8E9[F87SpAPRDGbAIglTI]KkZ5OnC`j2MOJ>f7Sj;Teb
hQP6\]lNeim_fR^9>9@IN:2>2=BkQ18kfHeXPOd>90N;Rn\hHc?`<QkKBQXD@;d5
NU5@j1Q5d10S_P[Uab1f]F2B^T:BlAfWhBN6\;Yd]j?J0YdBd?Gi1PLI<KSp9ikM
I7f<7FM;Ac;[27L1Scej1JiE[9N]VP[Mbg;Vp1ggk?\9gYK9KIF<glfLeWlJ=o[]
3Vjf:GcW<>PL;FM2jimZ6X]:0G]OK38G6d0<[BgZ[6Be?1Zmm`i:Ve?U^lP:8]87
C^hWP4fTAMJRBCFk0a\=2l5:@R5G2ojnaCVSn1P?9b2gEg8cVM0l3<G9m]X6MeZ[
KmAplDlP^>nbaWnmf2oFXgibhjT?f`Ro4KX56:UNnYl9^[W6MKYN?_Jk@eLD71Dk
=cI5co>hfmli=iXFP:aC?ZJWLbD:FGen5]FYl5JaOPLcWn2ib;c3m4dT\R_n_iFc
ad;0lAa9Z_c\YAna=OgX5g\6`8iNA=iQ8`q@3Z:?8mEANe19`E^@M<O\_1Fj?=kU
aNG1RIRR0Sc]PXXC?Oki=SXlVWh`LTX3dP7_[A<1_gbm0gKX10jRfAN<K?X>Nb]T
3e:NDj^B;FP01M:i=7Sn\6oBd_d_JX=I[h`@^KaWSbCGXee<hli_kEddOF<nAl]J
Xq?YEZUfQ422BTVQ6[HU_A=U46jQlf:WB?AdEZN01Nn8f>MSl4iC8_<5@k2_TJ_J
Sbih:OGOB<VoDcm<E3e4<efoG<@m6hUD;]PUL7UL=h@8ETnO1Aa:9=0foZD5mMMi
UE?:>_mLmghD]6Sb2cBe6M<g7]bc>7AWqTMo_6dgN8V>VD[kHAI5ii43GB<KD6Tk
8Of6eTgg9AJV?<O_mT]6U?SdlEk13?2g@NehUPBjl<R<N9dQ[^6h]CBGFdXP7[Fd
0Gbg20VB837RdLKHN^HHeW8omk=;\SJL?Tf8Bg79e:^4E:PhKk4ifel6;PPhZXMq
9hK_h81iAjgh\3Me6e5ZQeMLp`X9UEJl6j8]B2SBJE2G0g19B5n?O8e[l_nHW50^
ekX0bBKAJhKJ:QhBVP?2322TAj<1jflcFncMIU?VWSlG[:a?hW71cpE2b=e>Ck6j
kolQ5\B?Lb\g9j_gcdSDP;Z=R><H^Nd6BANEC4@7>73RNJ^X<IQ73SP4:c35ENI_
^=Q4J@9<5SZ_3AP@g;[:dFZM;VnBP<nm?9k7<<3]RQf6BRdo<loD_81kK8HGhNK]
hQ0`qNjOgDZY2PQE<<aUgC\l[hUZMO[`_PaWXaEf;iUNVJ>naQ2KNh;hWMJ^E[f\
2eGVZeWeXIWnK1O7DgX3HaG@4fHV4i5Pb4:C9Zm8Wc8NK87=`@:j9W=kc?^GKV4\
:0d]IJ8o:Ail0c?V971pheYhUEWFkBDmWRTnhnaDM4Z`7h6eiFSQA[MEcg@SHnRK
LiQ56NN4ER`nehHOj=fP`GTk=UDNc_C:kFb91TKQ54;Ej>JDIQ?hI]6[YaM\IGn]
1iO0Ff3>9DVfT_H9k4O9B2MA7c37E]SQS\q2gGQMYZnaIDCoj8Y?SGSJYaM6;SG0
dE0K9H__`g;6]o4mE;BUEpdnTnfnW3;32aWDc9?ccVgP9N_RZBcICm2P]SciUUm2
:MfPDDXao;m[m;JVEb<cV41FDn`KM\oX?TVG8>B;o::VmSjdcoJ;UAXg=YEeQL[6
[J8b`mM43G^H1idnELQBW[XKK0_b2iCeb8GAq>G2glMAO\LIg_Z=1Xo<1<1Rk8HD
jOTSYiZg\O8DkS[JhS@[PoC98O6AI4kKg1Y66LcBOV?fU1kZfJ]e<MH9PcL\[5E[
fVcGLk3EIoN]Q4SQ?9IR2LOaVi=7`JcKb4M=\b7AU?iE7_0WFiEq4KW@6SC3TMl2
fgVfF916aR?02]o\=m^[i=ZHTATeDlUaFG^>mZ6KS=D9c^mHN=E2IgBggG^1]0Ho
Yi8TPK29jYYCmK_mfZA0O@`lmnQ\F?5KPb:B2[kI[2[Y>YmHKCe@CdU3;7ADThWc
G6q:Kk2k@[4OnKKOQbmZ<L=X68AL6Njd05MH2J\cJdGReQWK[nlgNTADA;2AiL\]
O1ZbOaYTGW8lN1<JToHIY]T[_HQG0B]X>V1JLI`6]5o>NDKU85TdAXgYl^fN[LKJ
gW=K1RPgj=7hS1VL9qXf82\bo[KUZanho6A49Pi[CO_6lgLJ;Z0=RHYU@]<DQU^f
TK1RI\Dchn7TjK``e=Rl`?Y8XIfVekCN7k9Af_0JRh;Re\X`fC3bKT\EUFgAR;jJ
9XULWbEn0Ua;j>7^DZe;WBC3AXd\:XNlq?Egc5IUh>?6:VO2Y[9K<:iZjIb=kSjN
GoaY=50KB`?QQ5obYe2b45E9Uk4?@l]38ADV;I0=33KD5\;mEGh>AaF>D\S96j26
pI?H>?lc8>=h8AEU0g@GJ<KF035\hiR:9EPI_8PT5W7jKC=^Qm=`_F@\`^0c6P]V
q1AG4Q357mNg`[cWK<:IRX2iDF^LS=0_3F6;<Dlb`\J[XWJ`_3WWlFHL:_@6DZDj
Lg\e`i^EmMT^O60kUd\TXnOWc_InE`i\_G>;SE;A=dYm2mDPa1e=Q6;F1_2VXUOV
0f>7<Z?h1SZ02]2SXd\TXFm@2:kq7>7oM6G?[V6QREh86?Ab_7jeFD>BhK_?NkFK
gW9YI>1nV=0gQ=3ZYKm[8n\EPUA\1D23TimTLf9O_T1ChWU[i^F2mc5K\PeVDQF?
=JTP1R=J<UY3OS<bC4K48Oa13D58FgLoafJO67a`IZN@hWU[02>oA6p2PG0YLTfo
1F02<SKB=Jd_k]Nh7TdJo\T8Y]\N?n1<P_KhhhUN>ZbmFaPK@:MVJA>X;?M?ah@_
>VLkD0_^:D<^>`BjRXjO:bd\QoUoeO;<lZ69IH1e5_WFB7XOemT2CK^gfgXJIGOj
?ICfGXS^:D<>d2X]:pK]ZlT[9L5Y5PRCk`N3?29F04Y38D`BGQI^50ojI;fPF[YB
jkDOB49=bcoBLOPIh8>lF55\HR4P7IBNB6Rd3[mJ\`Pm3i?S766>PLIe55<mcP43
DDeSnIHGH4DO5<OTaB?\VGmO`fl:>eIC^mRd3[e:2dHXqfo?\X0SabD2<fNTNmfE
PFNUg[K2<><efja5fDo=Gd=jL:V;@j;8;TiI6ZafB7dUZd59o35]eZJiWN_Lldb?
mKb7??ajU?;nKmXeI:N>1eDW6gZ^nJAZ0D_UF_8WEEDnZOgI^Z44C6eDnR]mRdb?
mRUfP>Cq^b<ii@SUcbD7hC<ld5<;1BLI0:?2b@Qlln7S?Ao4P7h`OkQJ5TJhGbiD
[QOnFGlA^ShYm_1<`L652b]IC`DUlS@O3lD67<lBo`>dUZXdPcOX^JJbg^ZRYTDC
]e79;JXIddLY5\ldiO39\\TSC`DUMW3X8[qaCk7S7R<mj^T9d6=K;d8NUJgMcST8
NAJ4jX1K`>@I8nm<>=>]Zhb2B5lQP2oS7EL[U4`J23Ho490Pm=D;76mkEVl8QfOl
M<QV6X^ij_cj<67@JYChh[hFGB>Q17o3<N<ekn2mGTDS3ml:e;2;76mV5mT66p7]
LFJeE0j]Kjj=AXR6F7G7K4WLJ^3AcnjBohEhdnJ=44DHI;gTbc:k67FikAj_ALc@
QNn<07A5<Hdf@6U=ofOb3T;2hRkNQBikoabY_gj2kViik9[``jSXWTFJ<VQ[Ij\h
QYlENiPJSXCl8AU=of_lK\`jpXFFR05?Z=FRQMT[aDW81j;P^@lHekiB]Yo8nF=T
8RN?`OflCG?oKgPDhX>o[m8`3bnQ]\:Y:SKl2m[4Z;PTY5G1_I0p8aifDe6`Q[m^
jT^fF^U[SJeZc6^7Oi=?]5^HB^^lZh?J<HIYgi8l2L6p>CiO8f4;UiJ93EH`N?V\
1JP`<`HIL4B^ZF0DR]gl<IS2=Ane7j3Z4FC<aP9_L3ZnMoRgiLd195036@QaC`\E
NeYm?Kh>OZ;EYXHSl?igf5dLek>MJ4GLQ_XB>QmooZ;qK_FH^ZYO`YEbWVmOhlg@
Gl`XQFI`e\g83VME2UJ>M3HDPEJj7[0NOT;=4n7:MMa=PV`EfSEJGT`XZ0F2UUmS
T2\2Ud8W\3e^1A<\W??:fLUkem3jg87HFc`E`Dd@]cCqRTOXkjW=ooRhIL8cJ[Il
hNJd<_INmD20AYAe2MHh172LQIbHh_WZaj4HFddkGVPDg63AES=?5b:Y_CW8`nDR
9aB>e\C[IP2q?5eCIR>SVQC6XW`C3CR_MhJc2g5lUY75E5oEHN[_TAX:KcJ69IgO
aRlemb9N3OOKXJOYB9dX]=@6ZGaD7DYP8e<>iRmU^D^=\0hdfgfU=[B;WoR\5XA0
VIc6jF9cVEhp4:chDU2f_g8>aS_kba^PW5WYVeZ2q\:fYR<aUf^Yng0SZemR;7Yj
mPCZn@K21KOil9EHS[9:;fBJP]Db0E2_]kP[3A@UE=JBg^@Sc`hTUTZJV:5X]e8i
K7oiN=N24WV2g3bH?V0OIg`k11[i0<7;IIbKP7lnq@?8GaRB]T12MHK`TH_mkMd9
IYMOMbPRI5PN6VEe40ej1Xca:RGH8EQP`[\BfgRkJOm1:]<T6nPkCNEJ5QYID8ZU
Ne8G=QE2q_ZAB>6^G4?ZJR01hEYgDjJ=giKc0\^9ACE;VVm<^3cHi8il`^:IikTX
Ik@[FjWGH_Y9EEcJ<;HE>L]=7Me@ACW_>J=7TFLPm<c4?5LRejVNaU=LfM^5^2M2
qLe7K4RW1Efe[@\=fGJk60_1CA`_R=;1\8jo^?Uhd_mSTMilLR__[21O9fNP9U5M
TLm\T:DFXOYEFE;RE=W4[gTRkI6>J6XK93UM_NIcHP?OE3bRafE=UCWhq7dg?\RL
23OU7Y9oWSg\LAh[d9b?kF]lnk^_AC:k5Lb]4EO\CFNNHF@?3Yk>>mBOS78?=L^V
VM0@^LR<=P1G87`4@^apolZ8=Zb?d8<OUB7Bb\LFH?dOo<4MA6ZK`8DKciNGR[AJ
Hj0^KZnF@mhFWD0HQeIQ]@Kh]Qc3a[<oC_5NJJn`Uji_eKWjRDLhS;`5G]\F]QJL
X`S0i7lOG2_EVWg2NMDpoVXD@<bCH>>_Oon3Y[;m3gqh>8AJU>G@hZnTBA[EIJVH
3VggK<FaaMn3R<2EZKSG?:DP3O1e7?[a4e8TAb\j^NUJ;;3CSG68WZLW>>DW1gLn
3;<O1<RfkTZHaaR6ROJ@[5OdU?jM>:X_N3AWiCH4>bq;R[c[S48iL:FC^4bknmJ?
m6ad@[lGEn>;N[SoncfRL1G[hReE?lhAVkE4OKSe<QCBLRaD`_mRX:jMYQ`GCnFM
AAIU:TX1@HpZW2V6]XSB4CJ_STmm=_j\LIN\\D`goDf>[7\LakPGYZ_4@`M6XhNh
a4U>ZHdcZPllg3QS_`P2gCF;@QUoA0DP_I4^JHT5G\6V`Y=`hi@^bH[1lF[OjMg\
cPb8LnnEKgqGBJojhdK6[<m_eXGcDEV6f=5TLL[hCQSB<81h3XKD6UZYh2F7Mff@
OdCAnLBe7YOCb=@Rckl5m<mY8]Fd>m`RS[^jcW9HREj>9md@^S`>3[IURa:j?CT_
GQj4iFe6<<qANS=XfoHjDL][a1jd6j]cHLHohi\NW7bNa:0Z1[fh;=43M`fi?9O^
3U4_M8XcfLIOO2oI@jKHnL]6<QNFB9<jZD2;R@DINKqe7QnQ<7NfO\AnGO72R3kP
_qOU0`W`DNLh7HNXO\VF_471Dk^4IWcN^=CYRgJfnlf2oFICi1QO?IFP2A@Ajnem
LaO`;IO<[<bHc<m4dT\KJV9ia@ad;0l8h6nDc^>W]KMag=7imc<YiJKMapOOMBMN
M2_6AGlH\1e5bP>0nF@Ijg6Af77SWGM71WWcG[R59AHmGCTZNk41Qbb4;GO3=Xo9
3KLiSK2YiZhcGFf<P8cGdgo=n?32kOFDIa5JHPdmVIe`9K_8Rp5hWOAdjYY81I1k
?WW?dH;jdCPjCQg6Y1LGY;T8G_P1:YlYhWa\W=P=CI8Hl?Cc`350E3[]@4TTkb14
Z?3cWXg8aT_oqK54W``pXf?]GC2$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module FACS2S(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;

//Function Block
`protected
=a3TXSQd5DT^<EVMFE9:RTDP>GA]omog13`RBLO1YYe[oG8B\Rlm<XGgBK4BP[Bl
I9hXm;M`phQKk3UdoWT>=U7hPb_\JeV6T9>KQ9knNF`B2UU=lZncAB1HqmdCo;ih
X:0hiSgdX:?:o;>Y_0@XBkghOmAcTjj0=\SV2AYP_7ge@\W^37Zq_T=IZmqA9[2^
Xp_QmCRNfHcW?;iSGHcL0JQaeZN\CRaAhUZU4VB6>Y9\M\gCQbXQAS0WI8J`p72?
T_`pQ:STAf]C7V5dA\[Yom<ODnWVnXbBcOAqBX^aVCLXYM:6H79FK`c;mJZfWHnn
IL[cHSmRpm]b\CWNL8\7UIl7gNTKRB<M<g4HH[GHpMIOHh7q7fS2ng8[V`n4E2l@
TSZIULTY[Z_]M^<j2h]YQiWjT5QmZZ@GVmRXLa<p1:QP1Y@koFhYILOiUQeY\iPZ
kLNMnVPUm][DqSBoPijcWQLml]jn6VejLk164db:_hdKm^ImlTDpXg6UZhqIlkHK
90`^WgLBBGQi<]QBD<Ll>`kO5VCn97na]nmi;Ufl>q@a]49MLeLPDM=Olfmbo@jN
iTd]mV[=N??89\p>nPMlICL_J5?a5ifCd5A4WjkdN_b71E1;@V=E[qgNJ2:np91X
8TeimPB7N=L^3ddb@JUUSS52>?N7p?TbkkHGRR1b>lIUbCOPbYGjJ];1\_8Cq;j9
83KdpE0ZkGeqOCm3]AJ_9DWKVKK3A8M<3ZXOF7]AD:n`hT3>;hkBjM2;O?3UV^=N
?3X1bKhIQ4oO3EYc0;kbLa4a:Pe2BRQYhE;IBj]5hilRmfY<?2fhBPdfILdcPKNA
mT`H6hhI@0nNP@\m8dQ>fRYRcCp?SMm8Y;o5\]=nIQFHJL:a4dZDkDfV4GilOU2R
Mqdm>oL83e:?[3\NXDI]VlLb0aT__0L;Gh36R5@^UFJiBSA51E8mHZYfOHk54M:O
`ogj0TMGaWjhZ11eVe9h=D1?L?m4<AJ=K``7V;?Sm<?AJ<8Q]22OW[nHLcX:4adh
VO`gdfcROLJMf@IbqHnX888oN5RDj;`\8=;i@baKm[Q4DK2XD1]bWXfKF6=a@>9:
3g38Y\4WhC:I=6>YA6Gm>;`3li?0ZO6[V@G=Gn:<C??h`K7f2U=b?`A;lH_LB];d
3fCdPT<0dcGID\=;8KIBn1m:jh\I?KJq\0?2`4jPNcPJle\`J8DcV]S2\78CAjBc
OT5iKc>XJ:U6W=6lM1VJ6=iM=@oGicPI680;\^5alTkajF3^GTNCij<>A0`HadHN
Z8W6\0hcGlFPW5YU2BD?kbNDTBo@YT=j`1m0I]NaId_^W2plfoV3S2mI\<X62KM3
o<5aoO9cNbkflGhaQgmf^T\Z^Fig3GWSjIM^N^35GklZc@Di1CUl<lX<g5CFF>NQ
8][O8ZMGooKOPBQ7iPXnkg3Jh6edW5VL[Zc_I3@Kok`ZNA]ZM8@cf^MhTOha5qHn
Dl9i29Pnd7aKE22j7_WX=KYQ\olhEcU9_?KZ^4\jB^oMLKe[S3OP\H[_RU^099A3
T=>KXG<VZI[9Y?`X^93E\AjTc5MFYB:X8O4lHL9l6jN0eh895G:<XbFBRMglfD1I
di7XPlR4:\kKpABcZHCUO\l7BhIRoM`BdSCKTH;5@;0laIX6IL][E`MYgSKi<LEY
6OL]M8Q\0of^YaVITaoam1fbnfj825c8b=K8<`SaI;SYP05^U48_ncP:`ePm4MoE
>lb:237\JoFTKTX7f=Yn79]Lb=YpUa4icncYJ62o>[@U8NKN\eOT590YVo]\21^@
Ze=UAmRSI4J\jIBm?EB^g>3?PJS8RljoKkARN`FUF2GeXV^BHkG>QO@@KPTXS[Nj
l<<1NKT\dF\54m]hkmOKoL3a3`eiF?gk5OdJ[KE6OWqD_IT@S]?JP\j4;\IX?6Fj
oB?1Dc2Faf=AhH4D015gO7AJlgIWcA=gV1WFBZIel>ZXJFb<`BK8YUgABRHbW;cK
3OY377`_a[q;TfK[bUi@DBS7BfoGF>oa677M21VG3GY=<KFg1>>h;I>_D7OlBAdl
T=TnjWTQB1Ub@:2?gd2<M26XcN8dWR[`_YLj6DJn23BSSKmfW5F7`5WB8QhlOi\T
WU:RX0PIgDB?Xb?YT;j4FjQLbE_:_Z0QTM81cpim7H0jPj_<V3SgEFWkm\TTj[XR
74MHW8^mWjOZoA0k_Sk[U>q9LHB8d9CQPY]?d`o;12j\J9KHFX\DKIiT\1OW;bg>
]Y`>`j9G44K8AN`^;IKh`OnU6bc\R:Ag9:YC;FS:WS2n]R?g;eC;@04eTS_0H?ZB
7hMm7;5M_:gc8fOmV?4IBI?@BoIB;R_`>F?1MiUO\bKDPo\MbqXi0Y`MW:5b^1Wa
j[h]h<W1RjZg8n^dbm9F[lFGD=B2NA8QQEX;j3Q?9m=NKXO\T7oGL^O7?kS`LXjZ
DlE:@0][FLcGhmEfRibkAWAZMlN[N0NDoY\NfifVkgJW=JX2A\DP1SW9CFe0nBkQ
]U=5obM1Lh;op^3J[kjl:n0b1^?@fl_dWV9I[S4JZ<ZlTAl29<cNbnO<SbXZ3Y^S
@IH2=5]59dZa5;B`Jn9]?^JJImjfX=;_BmdgJORmaoD@22g2e^JSGBoAff^hSkBi
`B:Q074ONC@lmcHYC;6ek3QmDo2]8X7\j68EJ@5p;bIhjTn=V:Q_S5l[WA`LFOWf
`KmJ5ac]SBOZAfkJY:lIWf]59QXDcRWB2X]6[oVa`UCiahKcEZ\DhMZoiC3ZTO81
T7YcmGog[`OlCXD[5RDlZA:Id3]@92=e^^>34jQJ8KU>QLW@\QgadCk?G4HVc>b0
Q1p2ELe]UBYe\c^3oKG`Y>a3bY5R2hnQ;XJFbgRoL[=VS0XG;GbcLTcAG6HU]akf
DQ25iFo15`1KED_KOj6[]9UWbX<<_dQGRM?[Ag83n<=XhK92=YM<Uac98f5ZbEJ8
Sd\<go<Sn?oD\MCNeFZ3[F\L8[OY=p8_jOG3H0=Vmk`VhTO;cEeDE<QV7JKkU3i^
XicEZ7TbpHBFUZ_]3UnLBIk@G9i[4c@=?5WLOPfR4Y_F3<EER`G=II8^QoCYNMI0
U7]o\G1MaTb99DA8QlZR<CIN:15EO_@YkH8<WU@=9_OF=YPg@WAZVLo7YUFeo3<h
0=OohP5G8lR8gZ<V_PmMQ]medli8dk8G7Z?q:jnkSVfa>`:aDKSA:;[;X2ZThW<f
_jX0fJ7eN]dRZJ8KS9YOgE3gSTQ`D`0A3IBakb5PCB:d^M5ZM<VPKLMQf2Ofj?:N
;in1[?7T3o@T1I0Y36NDEmLVMNnG<SdKHZf_\XLTk99LZbmhEO68oZmVMg<N\dq?
E69O9Bh:mF65n^9_L3@9jmQnH@8NWABPIBCDXV3aU5L9Rb<Go4n`WKd@AG]TkWYI
EWAD5Uk5\i1?YGAEdbKl_GD9Sg<f[]U@@B<cjUKNk`Kjh2f\JC`X1jGRX?cYB=a5
ZdR0=j>?S2PKGhBHlJXc37TFnp13QD3:TgNFbei29j=7ooR<Yd:9E9=0>h9GjK89
iS7LB?OignXU\:>NB_Ze@_7g?97ObKQVlR_Lfc2Wi<i=^2k0Vc22=<AUG@NO[ln:
T[MW8H;`>OBS93oM[`ZM9GND[iGcemD:SUOQi^O[3GM4@>BhScVDq4bMm`D`HG:^
J58PD:a4K\4[Z_n7=Bb5Gn]=`H^f:8`f:;2YgkmIN_mnYq9jWeJR:YT15IC21<eF
_Tc?0JfF>D^C0mjRV4:``FLFBjJnO5<OI:O5Y?\8XMA_MC?V@G@IKY9D\0lNZllb
ZjRlSlAmb@F>93c7SZPTY9`>MeXLiD8GfiM6V3o:2ZL3Y90>?IL>1X7H`a9=>a7E
@;;_R]fmqVU8VeHeMhO0E=jhoe1a3Moo=fK4M4f@6l?Eh=ZbZfAi\h=`CXE6MZ3l
Uf2RcXQ`TO>o0:lfZgWQ@HJ>Y>>_;<>AEihD>O3PYE;ET70nb2FFA?GC11Y0ZRYM
l_MgYM>`5Id3I[?EYF\M>E>a94Z2S`k`kW7qZFWKF>SH;[<YicHCDXhC4PCD\l65
W\h9i;0PjDQ?_8l72F`S>Da?cWKOH3X9S:\eD\3FL<ni@ij3GWE[dH0c=mac;GoP
Im;[0D5K<@T>Ee[hW`EUZoNe?JblO^_Pf_UV7\`Z4B\OgUR0f0REG7Rh3O:`7_p_
11NTR^3m@N\IX0kpHo6jFQ79b?FBYEl52ROAbYUWZ1<34W`e?2STBFG0_A@j5BnL
kQYnc6W4UP08mMRX0Vo2cJ2A;@ZU=<5KD;:RD4gNOjAVU1eZYD21[:bhI77W?`Im
B49Hed8Uc=Tmdd2BXWDb:@jj:LPHmg9]EgL_[hliigqNLFjGS]KfSb4KT6JX?S5l
\mF3NK\nU4T43M3P\l4PP0IliIZlET[lW99DlnK8O;>oh>hK>IOnD^nE:8\^\;JG
lmo@E;NjiF9DhRfbhYL7N9?e\TUbR^V<9=]ZDi@;78:<5Z\SYEBi^6dfRD0:ESBe
5dNfBpX^3BjN6gZBDSBj<UHhKLRHEL6Xl2nm=RCMaIX_6`M;j2X_jYU7Z?kNAUoC
`OWK=9Plh1=_=aZdRZ=\i2<2b@=lHOdK4RID19gl@a3A4ekhI?jd63T`P0:bZJHo
>TEjM?aFGHa5>A3@i\je<_i:HED:F<mYpVRBabMYMdi^>dL?[nJLdnElo^mKc7gX
]@S8ne45KhV;fYh7o3;OX6b97MCNK:Xa49F;\Z2iN]7OBZG`e1n5C:;\ipXC`FU]
?^L8ZR5FhVE]l6ROQ;`6V@mhJ3?kA4X:\[cJ>ikkXYEOiEj?dA2SBJLWGW`F9I@h
YQ0?UdF9l4\6CGIm]]J@jPIlB2<UjCi>i\_LQh`b;F_d=bZ8]^SN18LZ<\XIcMRM
PfFSMEYCHOH^\YQHh6^Xaa9JpFg@5:]hVdeXZjb2m^IX31C[hNAl]RP<`B<a9BfQ
0I>H3[c2;NRnlj2c]>MilK4g0oKa6N39IQ[c?_3dFBZo4[>jIaXSS>Y6bhMhJDn9
aI<`hbmHTU6FWRCfi4]oXoY<<FDik@66@cdJUXMBl?[g5a>IUD1D?k6p\Oo@B;R>
mC8QRcDUGTH53HW;kmI6EeH\3OM:<J1DTGcSFgg5682c<5B_iQ=5HONP39cfD8Zi
gOomIijES[RTa0e[ABNeaPgI6okH?fCJm7hN:a3i_b6\9Sa2dF6Gh2IK\Hm;<65G
3gi?0S\hIQPNk5R2\Wmd6Mp6=7VIGKQNVF_oWGZ;@Y;VQNH=YMo8=k^3DnZPEB_d
SEi_`HAEH2o[:E]hhXeNPRji:MA;7PF@X^A^=<Enk?jcC3k_Na7YO5VFXo>WKPcB
hllj>4lm9iZfK19DPQ@QGhS6W`PWeN<SPVjTf2YYEfM^;m074f=i?q\\HO=L3kai
LXWk]^Q84V1R7nl6IWJ7C?mmXF7e^C7DibRRd;cjn@d=fKI?iZIRWF71p;QaneB0
B@<ZH1eWCE`<he5cPGUFk^SG2Bb1NF[RKC\_[oS1?2>3^:;hO6gT;K1[2FBdO5;F
ZXmFQm44]lTX2QcPJ3@BKmYCMcQ>ObQ_9<b`2LN_C:=W:l^bAH^;e`B\C;:TYciB
QW0_D04G53d]?fJNC6G3W=dp[P[meMMhmOmM4Jc@;^ZfnB2_>3D>XSRelj0M\S7X
6bOVnn_SY;MK8PP27jb3k][EHMa^?:hLa>nEoOG09lWHfOH\f58Ph5W5YLKbkc?h
9gb]2221L^kVkV3Oo@eKPTG4[JWC<<]bKTWSk\@^m]jCm[^jL1Tf=ap<GjY@j<30
kS6Snm9J7:cmX]bVlPcY22E]CTO3\\KecJ]kIdODL\;=\oB@m0Cnh9bE@m9WL?kb
dhAX1O`nWa=cfLebK^9;mkn;5Jn[Yl\EQkTJ8^]94Z64de4;hPUSJ6n<C<7O_W<o
b?<H0;Z>I[<^UFS\:5]FgphFG8;7UDL?@_dWbJj\2m?dW@<\Q2AWDQWMDBP4k104
@a_TdalWCCb1cMnkC=KiNXZS865U`73gZDnYGkLT@3S:8W`:^Rcj_B5T?7RfMkGn
::SJfZjJefQ4D_om]Y`@oghQMO<]Rca7d>CO6QbeD`dS=aTPmha0pN3[l1Tkh=Da
D<eF5ETa6RN122MXG1kXhf>5l8k7^6MbI92RM9Ro8I;7<a;[=6CdWAF26oAbaNh0
VLCCH5b6JVl4]j`?kALKF4hYT_W61M=TldZXLk:E`gY6meOTHiD`;NYBCP>eah_Y
:nWK6]\Yln8DhVm9PT?qhIA`F`biC6O[8_Y[`I6`S`nbi5cafIU?q3ej7TXTZHAP
:^miFLSML4DLj2K;5QRn6FFRiE5Lkfj>80?49XlKQB@e:?RN[a68XkVQIXDIe=@b
830[<?\c2>`Oe3]\4hU0b:4^mUZC:6W3DKRQTECZU`MG:\fc7IJ[?3c3kgA6de=X
`T>KGXAdocZ5[KXTi@`qj4UmDi2KfL6[X]LAU=H>F`?Ug4=`[BlQ3QT5P;KE1LgF
hK3=7V`Qo5lEA@K5AGCS[<>PE=D^CUBHgV8b;7SOYPf<1LY`9Mo@bINCmNMYW40]
WfSfOUAWZlBf2b\J>E1njf^9G`W2kBo?dil7iaAlldG@FGK]`_pNEZP=?RMh82SS
9ne[aIN`[K<\FDeA]f1<>8>fWE[JG2:jdncBUf<X6^1;\CPbG`E[3<\5JeVba@kO
aC?aIj61N8XBDf]hKTSY<CK\o:9K`dLI4P2JN]:gAfS9hK`n5iPNOJa2_kR0V\k0
@3H?32ATPF@74o6:BpZI6YWfN0hn:<VS\\G;IPdGSTf@j5o>\?goYPkLbic5`om_
MQnXeUa3:lQ\mHWa9h39TU<O76JMKIh@I_BU:EoQ[IDj[SSQ=?[@I3LQ?Rj0bKm>
1dZA5m4`j5f2FjM>]KZl1PNgmZlmE<i=^RiDl^cl>]mXVKdjp\JU5C6?=:>h^Sgm
Mf:`4j3Zl\POq]=SYLa0okg:Bam6OJm=hi_hQ]b=ddSRf8_Qbg3mUMN]Don7_k>]
]IBYT<8OmAM95Pn<ZiWXgGZ`238^9;Q\g9JkWH3d38DGiI\3;N6=Q=e0nMehcm9L
G@9I2;\nG7Jcc]N4VOX7;0QAEKnBEel[?`F`FL71VM2pnIQPmXN9`;AMAFPF4C25
4T30PMV[lAZC@Zj1CcZe\k8ZD>AdIN?i?2Y;BFXb@XZFf7WZna0:E2N@MYb@l:gD
KOHYIfn@AbF;mc_71P6XZRo`0[fmYUYZhBhK0HPg5AXAn[f9MH\:\[_GD@OECF9m
[<2:Z^`]_Iq57OT[Xh0a[\ALmni]Y0kVJS0V1I4kicDfme>JF3WIon?20J4?PI1>
bKIdm64eFM:WkW[We78j[4em[Zf\_4JiSiO50T9HS4kTh?lVmmWOK0J7eC5YbMkc
HL?NARVmDo>52Rb8ILO1HkB7l_GBB6GgPgR9BIBeRpSOoc5h83O?7d\BiTAEDPdZ
4bKOLifFGIS6f9V:K<h`Sg8I0?GdRfATE8laoG4JA]f1WS>R@?:Mf=YL5:o`3FRX
>UaBQSp[E8>^7e]V;8CTmH>\N68`baW4\oi1dKBlSYNZY=NbPlcA`9G9QMlM^_MA
fK1SkhffJK?P<7`iM@KU\7HU4U<:3?^LQS]Km:IjC:@@n`DB_2C=lW\ZOO`UC`Oc
9KE\lW^WmM2jJU6?9H>edpIP]M=HDB]VdOnPbNY=SCmK<PN?:l`2j1OV7bl`mC\C
f;HaJg:02HRZZfPj35C\N9URIh0M813V1Ecm3[kim[UUT>RJI71\ZoZS15Nh\6=e
B_L@C<B\S]ckI]E83EaFDm5GSaVLoGToB3S^pd`G\VPT81Kbi^XGMcOMp6XE;]?2
OJ1^;hkPBgib>3jVj32oG2aGbQ8kXJeV:]e25V7d2;<bHkG:2U6X9;@Ek0dMU8T[
YiS;MI`NN1:h53XHBb<fPg1LkZI7`5Xli<8UT^:V_an;maWcW8hX9be7U]PbM4nc
^P3MTm2qY;HSDn:XhKA3bDFDCBIJNhg==CK;QgKbejNI0MLn[TOYKeInPP@KG[LG
dO8h5?kin2aE_MC3V^d_US;SYlCES[BceWk5h:[<mhF6RKC@Oo5@c]ML7kAW9;SE
kD8jIVf`OQ19]emUXOe55aq^CbVEoX>2`UcD?n6iDkIYIO<gahb_TkbCdE:ZCFF6
^dUDUioWO\0iA3hKY6YILF3FQZ\\n:9<o0>Poo6[?fIY]>UE^GMMYO:fTZQD:5OI
\OAE]mWKUW8XXLhV465`=kff\hPaF=`_W4KkbqI2Tn\VTH\<A3FM9qO4hCU?Y9J[
bU`cJ\SikTL;<dJn51@Q@\oROJm[Hd]a`1R[CR1\nKlmBdQ\cnN8Th`jIRCoP6OO
Dd?C@[CXg@eB3X3JmA_j3WD`JFGQ`<fn=UP9YDM`d@X2@1cKcMEhh]KWV2:nlW\E
]WXoqJBdZNLZVfE`X]fAei530DSELVlG`MTQJG7c9D__cbU\UXRK:9UAE<Y:@Qf0
UEER;8Cf=[ZI5eUnJLZbEa=iWdm2B^@jB;AoDAWm^HY8;:2@56A6T48P_f[2W3I0
74ifKcD=Y16in6?0ZG^plQ]9l7a84UW=F9_:QIYh@jCJoHQj6V[PYLf;PVQY;2DQ
^2\C9JInJ06YORZ?V]G7Y`Mi=4o]hcIiE=Um9UnQhaO>L?_g_8RUH0MkJgLgZ0[e
9>He@PiN1=186`Z^`ck6K26Zi9gCMjmFM`qDkY=99<fagBLmb9NhCOoHSO5D;boG
\S`oGYQelYYMO0ClNGQ=\76VTF?eab;=^ODMoV^66RRO]2db7[72O`YNK8LJPEJV
<<q;P3ACLK0?RE_R8YJgjcWq4=6amVKIfOdDClAJD5XlVN7:GiU;OE7eO<8K4F_4
UAHMV4SC6:4I2OhB_;S^^UY34BFO2J7_d9f[k@nI<cWG^gHc1IJ7;h7hEdL6fk:A
13mS>NJ@T\K>2eoI>cRegNY2Z3ee2?UTgH3ek@nIgJgfKKqU8ID0_?3OaCO\D8o^
PPb4JG24X0H39CQlVD0dQddRfD[Blgfe4dH@Q8UW4dUfZIaU2ZLUIDWnoQF[YNf3
I7[acVB^5fWRSCH0mg60Mo20oAThVh00fZl@UVM?1m?4VLW=^4Dh`N9\`Y?[YNfO
kdU5mp<>cQl[5g:W0;fKJ=<hee:hZ_7j8[>he5;HSC86cHlG9fB>9kk6QZU:OVPm
YSY2YO<40:dO]ob^jHD[N9jA6`XGnM<j[>bjeCi\Fm4UTaK<;_EdK@ofY5U?3e;9
:SoC<SmUXP4?Vk;`<bD[N9cW1IHBpLUXWU1PBFEYGT>\2VFRaU1KYl0LDj^_f0?A
Ol1a@I4gciEoaMkJ3mN^CKKZB^R>VLJ\U`o6_XQjlZ6Mg3W>L[\P3:0dmH]_jj0j
FjHXQM_N0o4g[bT]Hm[jTMGJ>QFBFImMJ;9VAA:P3Z6MgB7b?M_p;]PA5le;l8T[
b6iCNe>61m_bl;G0J3Umee8JHcC1nnU;8@o:YWS8n4P?JJ^7XZAY;cKc4VIb]k6V
J0_AaY]BcW]SI;Q=W=U8E\[CmR`oUGiQbElF\iKinYEK7eb`l5B8_O^R9Z\YTH8H
J0_AT0A5Bcq7Y?QZDIDYnPW=DVVUQo=KMboOJWiXQ]3GG20oZWO[AG@Qcf51U\dN
^8p?59^`:QgGAmk;AcOMVH`MGKVSnMGoOO=nko3;o]B7`i?QkNI<1h;fFj9]dH<m
T0;?\nLUgH>h>=BkE]8lY>M@D4VcnN1:HO<RTOV>?>k^SU8Km5;ATcgf^<RcbT04
nol0D1PIlUef=_>kE]846Q;5NqQl7J_:TiKkSgaAdMk[IZcb4IJLjeiLX;?F>clk
AGJaV7ieY=j<5X\k6LZXFDd17aQ[\@oWZ3XKMEF[0A^G=YNn]39J]NTKXN^T]WF>
H>=i_OWZT_\6]k\:ERW83fnY_0YdoWe1HkQh\:F[0Am1giHOq21ULaWQkHUjcJWc
@W3^m>[@U4SKgKNVXe94VRojkl^HUhkbULOH?d2F5oCUZJ2WL2O>Y4h[YUYLM5Od
J99g]?22IXL^_HkV>Xo@RMPTYS[J:l<<1NKT\dk\54m]hkmOKoL3aX`e\F?gk5Od
J[Kj4WWp^UVSBF1USaoLF1J`@Gbc\[h3hM6dPOmU@38B3f;;C0kPEYH]L0]=GdGN
T__a^Jei^AcS2Z4HoQc6WRM1B9EJ8KqIK0<6?N<TKCVi9n`b3H8Z_4Je[VdPjZT0
IB0GY7?ghd2Q47K@c`Dn`meC@EYG\kb;<1<Z8ecj[9J4l9VRSPE`Z[i1Zai;E1i0
naPX5<7aba[SL2VJj[W^CT1^Q5NL<0q4JO99d:LGNR1Cl[Q^EQT?6QGL_RA=IfKB
Jn^D0<ZC8_3WH:qGBKaE7eh>hUY=WhVD_Sa;b0^b@P;JgoBAnPckJ7d\bkn?P^^Q
T152Fh4g<8j9L4?KR>B3Cb\Wc\iigN7BC9kCW?TAFB^JnnNfmf0DY?L1dY]F`:_c
igG5BPXeX3kETOqRGd@ZU3hXc3EZhZBYBV?bDjhZQPLi4F1NJThb9c>KCK`3@IHj
H2jM@mod_F\2^PCVVQSgfL[=PdGmUNBXg3CCmPLE5]El<TpC@fVEX5<DJG8LLc\d
XOD`FbT:kbAC<EoQGVgek@2>3Sg3n<QTon?J664XJI;3RCGf5lB3CY3R:omRVkG7
Yd7PmT>nk0<Ja^;Djj=9LfOlhhJSC0fkHTJCL;L_AZ8I6mqj4J[6L[MjBCfFbjno
\D5o@m]1@ID7LGXWFT_?KI0AFNVQAo>VgTj^a3QH9@IROWY5hgbm3UW[8X<0[g9^
[3Z]fG^0_:Ejh^A;0_D;`3Cn3Z^PRgRWOK0k4hVYn4M:\`qd]bdR52_P<2`Y0hDn
E\=15<7VNUiU\D62\SgI0IMDaGE<IPE];S[ELGZmYIYQdegi3C?abOV^kQR<l^=l
XJBZK6jYT12b:jpmVH:5n\eSY9mhAlR1nKd_6F3dm;UYM93=;cXRhc98j1]Oi\XC
0U:NPVmg^92\KL9mKX2NK?;@][g<SKHATISkTJn4<@H6EjAdiR[YBL0LGe[S8Sb<
nG8nidpaHNeg@2C8BQSib_MXFQOk1IfLWfR4W;DcS58S<4jD`n=I=\Q;>in@76Sf
aIE>oSgaA1TlcWeP2Sjehc3kLSkg94P?Fd[CUFjJOZVLVn=ZC9Lgaho5j\Y3\5pn
Q419XE>WJHEmNQMN6_e3a7:l<`=lDZ2X;UjI3pD0TKSYO10\LCAdCZ=iW?hBlKRH
^DglAKS@l?`kPQ<6GIM1l6QMA59__IP29ROk7PDnnh]DPILI1XAAJ`2<o4fXnFLD
q]??=;_=;S`2big3[=T:43VXXHdKOMEfgWHX[K1ARe<??\0PCUL9fd[]Jl:F69J^
gOkI<@A<L\52:IUDVn?cQU1E2I<biMig?\L;gUa5K3IdS2R;Cf\VWgb7P?<KYn9>
p51<K5OUo4F>eE<lYSle5FF`k4=_`jT9oZRoUgl=g_3\`S4Ze<:Q@4?TiUflOSgL
HAoCCUFWh:P>m8\XmCkGSZFkjKgk9]YTk\l6_GkdaghRHi>jZO63\ABEh<Nj`D7W
qXOKRg3C0`DEo<`4c=U^GW0icMBL=MAVXZ3@37iePKPG>]_;]TJ[N_>ZfcQSIkIh
B]nlSU56GEME_3c[n\NHj9[dedS4R7^1qMlff<Q8Qe_YkoYfQk8@6cZ]k0D0h6g`
9Y7bR2Bn9WVAh8DAJDd43goWh4:5D8P>M_WVJn=b2gAYQGHUmQEKY:ZC5G]o43d`
m1i\13_f]6XC7Gc7Sh^jSVYd?l@eeC0=pT;\?gL>Y<AXe1[j9D80MMGo9TRS[H3V
4OFSjM:2h6[K<Ue8Afh=_4W6Nj]nNdD;e6;VFKlZJCoX]?o9ROO8M5QJ@9817A8C
dTZ`dZeRVUX\R\IRe0VJZ_g_h1IQC\4QqeJ9LO^dX@AaQeZZd@dXk4X`UYFdXdBZ
Gk>?PhWiTFG4]\e6c<E23@ln[XL18ib0E@[_<3]93Ega60:QlS@8Bbof=OkJJEae
pVAZ>Rjd2SoeI3]PAlJUXcklak>gSCfU@Y3N8E9=Y[f6H8eVRNgTJ;S8klX^E]jG
BVa>Z[d`OEB5[lhP9TYAdOoQDD70]aHM9YMQHCF9BVbXb@[\4[XNc`Rmqc;oUi^a
OkoSFA\IbWhLmJOjY0PbqCa=iEBnY1E_dbH;jXlic_LPPYdU<gWb?WSdAL^6GO?<
ROnFPlbRAdbI::iA7T>mXCWdCc<QbKX]X>mG78WaGbTMnkhQlMX`=GV;CPkGgL[c
Jg[j;6eYGOJQq6NM80Bm_cbc36`0YfDS5Ao5QF_VoP?PLT7VWf9m<oMEEX`jfPFl
8f@\g2Cb=>G4C6P^^H1O4lHVX7DB9lUJnd;=^[Cp3NY8XWphK6Me6L$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module GCKETF(Q, E, TE, CK);
   reg flag; // Notifier flag
   output Q;
   input E, TE, CK;
   supply1 vcc;

   wire d_CK, d_E;

//Function Block
`protected
8;nPgSQ:5DT^<5>XOW3bglT:Y9NqiL0F:UFfdAgP10X4Z9IK=TF=\H[qXS32_3A@
3=AKD;>[K]h:1ZGL?`1OE5oljnOl9=c3_i^AcB?:JXWA\W?f^2mFpC]8M0cqjL^Z
@`;7PCcV@b=RKA7RTNE^:21b\Fcmq^4R?>=0m7oE^K3?5QjPE5^j>l]_Zo4DE;o5
2T5mTLj:4S@J?;;DW4Z]AN7B5BhEXb]KqijN;8lZ0`5ALOj=07^Pn?4]1GOT=NCi
fG84MqABcZm]OR=j4=<n<biee0VZjQfoj_6QIFK?6ZoAZq6WBONgpWABhNh^pmUB
=nnpAM`VPP_a=O1K1=QC5eGQ<e3heSo=IME[5YnkC_P@1gCTG7S?X7W:A[6\e;[Y
[G^SASAi:HY\TE^2I9_H@6UnRa\]F0FMPBEAX;SS4^qU[d7m5047iIHSfQCV180N
AmQgA2abFHF:OcEhMS17kI6c4YmF8Y8;SH@AiIM:mhaDah3[6aqKY[o?=;TaPBa<
=mORGiCk[?nJ3AWR?CED<Y1QOVJk0:K5l?WRSC]?TQHN;Tm5^G1K??[81WSPlZ<5
?dRPG_]?>U2m^R@^>CE\1gY]>pX2LHjTC@`foDQZTPlFnA\KND`[JESn^U<cGaQg
Eb^W5G@0FOU2;e_`B;[T0O;l;SXM`n`i\TZIb`b:?>`BA[;kqYmKjbbpK>^LU6?d
N2HnA@ZZW2?La0nBH7>FRlBa8FSXh^l<bOk>TgccJjT7jblicIfROUYTQ;`86]g2
KO@KX>L_d<^K1WLq@1CX\Mq@8^=c>cjIm2jo19?@5XD]84NH;=Mn[NdB>OkBoplm
BLWG]hjE77DkYV12\5H6:N8jVQinCjMV8qTDfPFDZUB97ODDkiNYZiiZ8lbj^70<
GCDgXAB@47H:`ORWPBG9RACZ>:IPPjS;1D4FUg9QAaMU?m4b]j6AfD@>mc?f^2Ik
G]@26?=ffUOj50jGRn<Hm2DLX6HZJ2X@]5qYJ_YXLSjDZR:bll:B[mJoSD?`AE@\
5;Zb=9CaSlg1WMD2?UfH1hA1=:B76XDm7iMT[\<XmcaIG23Io^fj^bkQUE;e_i[<
cHJ>oW\j;32YR24a`kjP]:<?3I:[eKHb;@]pHfH2anaSV6R:D6cEFW5^]:PEdL[6
Pab9]k=LgY\Z;K<f9`H?pFnDf>Cqg`]X3V6NBmB2cded:HY>OQHeIIl7<CaM54;b
;7pLdA:=35h[VoD6b3V;2bfIYPKU9Zc_a_Z4R`E4HTELkhcX>n3n6BBjUAIk@W0n
@jm7Vg`Nl;>ZjqKo9=bg6$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module GCKETN(Q, E, TE, CK);
   reg flag; // Notifier flag
   output Q;
   input E, TE, CK;
   supply1 vcc;

   wire d_CK, d_E;

//Function Block
`protected
JHb2hSQV5DT^<n5bBSahA@Gd6e\KmJb^mOHnf40Opc\701`9j9fY1D?`?W<8<D;J
2MJm6\o:V6g@PH[f[;MRB0Rl\pi8H577ZB^2_cF8f>4\d:AkGQ7lEEC9>5oGp6N5
a4Oqn9O8@QRc3NCTI=cS;geACU<XjhMY211>p35Ao`:\LW[EPRkM7JIoJYOlCYDN
K<O1]\:L2[ZOF903C<RJ63k3FRDMLe7M@0ml8>R:pCJBWhnROXoZ1IGRMX[KJ5D_
]=9:=:N?5^@6SpiG>i?G7G?O31KC?UjaEX@4hk583IIcLTgDiMfeLp`mo0CmpV9m
kQEUqAA64LPqP7PkERC[;PW7ABi@\mE=8Ej;;Fb7Y2JV3gYYW6dXpHE_SEQndKde
;NH9jR`\EPk2<S9dhacd:c@l]2m;UF<`fl7RN:gHgodm6Cicaj?JkH\k2BZKbTOE
FhX3`E<[4ZgI@?:;X:0dNX7WHLhp?0jcQJfU_8oo\QWA<CTkSJgc9]h`[Ue4MW;O
_n=R>o`7MFDWN3[@@H;c4UN9KY`7?3O4:J_ZVIbd_V8I:MD3MCa6YbP4YTegG<mB
5CqYKkl@MhK0WX6\]WR1jOhcbI2?N`i]lil4;;>[\TLo?QhREI]@o7n[aL@b[WD4
g\9Y93l^hmQIm9ESDlmP<`4][qQ7PR7WpD78k9d@cCdln=Nc[4?Hf90mV>S]XLT=
A_b4MbADUjBP[]8g<0NF7[bC:l2O[_V3pXAOGOWijb:B6GLmmBd_@135=:kE`X\n
LWW;D9k:b3nTc\D;C^4JR\AY9AebP67OUZZG9Dk`EA:;N[HUI`6\;;3WpLX^eLKp
<@MKjY<1KWjQ`_2hi1;LjS[LkN0KJcZUiU>@]bpJ5k=4<mJ_O^7AAd@[WWAFn>=j
0EIH8IJTaVq;PmkOKYbQV\^:ok9<kA;2YU89SiO?jZW;;_V7S83fogTFiAGjU5aQ
Em\]I_\BjFgIkTi:QoHYQODOVfDJ]geecHfh>PM;=M_20]HLZQ18?<Q]oN6^^`H`
X@UPmii:ZdPpn\`Jn7aS88N]TS>3=XXT]C0Q9>3EkTVZImE;PTde16ag455WSc6Y
`koechc19dNZQ@4g?hQ;goNC2Vf<:hRFZn[j>Y@@6k;9Vf@?_Ib7BY3TD>IH7f1V
bC?D<Sbk1mX:pPAm6UaqbDoEm>PIT^0D6=NW^^Fc;<9V812h7jF3@MC^UPq_CX:\
J\XB`L1FOSOA^FmLLUo9AW6<AYIggh59GRYTd7>\@<ni6ob`eghNSIC>7cEAC:fI
IoFd7qI7X3?@@N0N[0NWU33U;IidKSNC4IP]p^`G@Fam$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module GCKETP(Q, E, TE, CK);
   reg flag; // Notifier flag
   output Q;
   input E, TE, CK;
   supply1 vcc;

   wire d_CK, d_E;

//Function Block
`protected
hgk9LSQ:5DT^<D5a_WEP=]:]Igf<K<ZY>VE\<6ahR=NMJK8bo;]?16pVmUHZ7m7J
`i0CbS]c=q[ZhMP^81J]R`g[GbEOn37QULNiM]d^]VBX3eGB5<gW`BVRSKcB?dKV
fJKN`@6je=]An<C<qoh\VC1q@JeCP_8@iSKP352V1@;i\ZOgIWThYmTRqD]g_K@4
WA<P<AQl71m4>\Pe@cmY@Th_;`jHUL8il<b87_UlfdhU?i9>I>;8OgH\a4H\pCgG
f;Z5PC^ZUYel9Xi[1`22J3\3\=\;\jeZ@q>QFAFM2e?`?edE0RmcQaFcgd`]7HL4
\DmY447K:q>L[T37q=nOI_0Gq43b@RZ^Teg2R?6Jej3>9Vi^:h[LS6E@;?>:0Z0l
pbDWYgdqPjAbc=jFF1R@Ijh;2g`1D37o4NB]GWg;7mO<Tme5Xc[\HS]gkccH=GC]
@>\X8:BSPgVOa6dV_12ZINb<AFW6?]gJ:]H2P`gLVTdMLIp>3iFH\`<2LdiQ@V3A
>CXBXClB76VC>lomjdVK^YD1^JlWUlOlWFg]I6IJf>FKCW:>[Nc::6;FDi@N;N54
P@C3]@gCQY\5^lk9Ka?Fcqhknccm0;8;[^[^a03`E0`lbT^c]`5`;]8Dnlb]9f;i
9Ah@\foN[9ki]I6H8_;5QdhT8NVT[]T4Sjfc<?a=fM9>p46e_ojqAB;NkN76mO=C
bhdchXFlnQfohNTMV?hKNKh^<Am84AREi\leYWPbUQeRi3^:F8Z4G1Y0P[EI5IfT
X`;]F:J5_8PpI@@kCeq@g19A1I^kc?g=UAgTIYmPk]8E<4?PhB5LW\6pbAjE0Pm6
Y>E;DgdAUdJDd4\;chUB2D[4n=0@mXp=61:RRFUZF;`jX_0P6kb:Zi?SWM`=FC<8
9>qna_ZKMED08CWmcaagLYYcH3b;g;jh;bM=W>:48RCo?0m?gB1EnaCIgiKY:AkR
5941VU_^g816_:]OR;2nX^dP9FO6g387eB^XAH`MDI`5:IF=oHGE55^<LR7:5Khk
H0dqoKfj1XgBcgd1AGWEKE_0\B`<if[KO`iZ5mNE0bhU_k3SEeZkTa\aX6GnoAcj
L_lLj8K5ITH=84C?kfe<FYN9P\847Y0gMEffUbU5k<8IhmfIiG0I2>4H?KQGDZi9
]ENaq]fPOXWq_eU61EV1<BeHn6;;ad4:D@4@Jh2m]@cZFl20e]p@?01B1bI[1@lf
1Q^Q>lR3KHhAIjZaAmbk91GHK0NDVnQPnYPCM3[olACGR0WFb2VK_n6CSaiKcpbl
ooAQ5PF>=FY2D_AafU?[k9b3e[RS8^6>hT4iKW^QR\7dGKgmBTWU2keAH3;Z`MHb
>1b=4>qNlMTe^K$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module GCKETT(Q, E, TE, CK);
   reg flag; // Notifier flag
   output Q;
   input E, TE, CK;
   supply1 vcc;

   wire d_CK, d_E;

//Function Block
`protected
5Li\ESQd5DT^<U7lA]V9VJkGK6fdOjlRT@hkdVKEmQG3UaBgU9:68e?ngmO`JKWG
XhGpmdUffoUn7^Ybf3mOo[a7m2BLC;_Q<Q6?fRg;Q>PqVTc`dZjToY_0]5K74>N>
iceTPbh2U5n7Z96e\LCU@D_6U9WE<QmJlX7h]DQgP\9Eb\Z4>`@VpaDlTKMqe_6C
Dfaf2<X4KJVOj<gS@?FO32]`Yl3]pGUQ2lAQ8?H6dcmbCARPX?0EVL?GbdGMT^CZ
f;HJj<WRDY9GMULTm?`Fe9mXb7T7m4HeqdLXM>5m1V@P@caTF1G]IL_5C58IP9@?
MSomnqUT`7O<k0Pln07kCndf^UVLKca2jBJlWK6<g_[R6pSMO_C9p<dj6B_cqWl^
YD=ph;l^98kNOb`WX4?D::1APf\mB8I6J19fqVj_Pc_GiOFPCb2=KIDXd8=CjXUC
>b\J;FX3e[f0?I<:C^D8Z7ik?V=gCIVTldSH\Vb_=kU=Ldbi;_HH]<3RnShc:Vjc
;fLJ;\iPKhnqX5cTD;PV@K41S>Jh4ccGN_]TNmJYX3loi00e2Cg7PK8M>B]1DBJ8
JcD^[niJVPXIX4CU3h5[jNN66@UjCC?bN;>V?SYOX<l_VWKCo_qLB9[VQ8_cSXG7
V;eGFW_BmjWVlH4X1`OBjSXJEUJ5>ng6R>J@2<Ja8c7TRa`i>kQLWhmWm`=KCo<E
5[?F7FTBmpTHRDNEqmUZ=dlbKGK=dYE6D4>F1?5@?gJP<\ZZaZ3iI9J_SDRf?H2K
bnkVB_1?i8ZKGcn<M0;P4D^SD7bUV\gWbF^iPIOap>6QN?RqXbZN?ld]\5@oC7]:
0GYWMX1QKNF2RO;>o5NZS0pXO98e_=:RUjWK3W@@<`3Z<27gLXSlNoTUIUpP;adW
D5<Q]7GfUXMMA1`o2Aj0Gp6Fnm577l]OOP:_V?ObMKIVg<QLD01lT:k<?H`o2SSe
J0m\gR]g]GNIn@dAo2;_bB\`LDg363ZaC_42FadgiLk4jG^_cIM6go25<JLI[3k]
h7RTMC0HZ74JigQRB8C:5mp9WOoPUI>2Ia9@VBjjb6;`]b9gXegMO3S0nZek_okj
G\iIHY0<jJP92VA\`]Tb32<dlR]B;]_=E2MkRa[b0<QR_Mi5K[0SeEhj_85OQ:FX
:3SMDN>deL?d8lfn?jL3h=Fq??7589pN0QjVe7ODDPM?9BO<\@Mq1@00R8F8EjBE
b<?_2jC\AWPb;m15_^JPWB8D48qR^QJM@UU<=`B?cjJK0`An@Rcki2\\`kl6XQEU
=h2D63lAUSZ0XBidA8?09V3cKXZi^g^FY2;Q>q;<TMcEP$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module HA1(S, C, A, B);
   output S, C;
   input A, B;

//Function Block
`protected
gbi]LSQd5DT^<h=`7m7V^nqX_oUaO1fPj7m3VTOH>cil[YlJGGI`P8e;2`AeQNjj
^kJ0URa[ZAlKC^95g0_aEVYRXg\qmNk:^m>84K@WdT^477N^M;iA]G?E>^`1QK9;
Kj:_hamoY5[JQfiNL;D`N8i6q15QGampFZK]4]WCT0PgHTnk:cWJnAeb:2Qd0^qm
VH:M=I=aA3]c]eNATKXPSMNT<03eSqjCRfg2<pCA75L^p<m?RgYNK4gSS_:]O?n9
WXhDQmD4Z]:cMk`QMCnH4mSaDf0\NRkTkZ4HcP_co?bJR<:E3?3P0V>jb>GNg9?g
\[5:FA\KjTLcQ4Q1pjV>FX[BE5A07[2^4<cBOZJkE`1KF]O5_Ugf][n_En\l?>=Q
5D@IEfnB2PFVYF=:VicgF6?X;0]g>FLC:fRY\QoJlQK\?P8;:hVeLPQK0dlUq\T2
R6Z493ic60i<mU\eG>IoacBb;`CZJGZG8nB62SWS]@jXM8cb85f8AKWDQTLg\7M4
;I>6k=Z0SRd\B<4enZYS3fHISpj>H;EDe;G9L8Q7RZb1O8K][D]]NL7GRDbi`ZZF
bcpXbRG8]cP3ULPm<nO=FHTmA^>OiF1ILJdQ]`dKYmi@;i`?lPkSHm@eNhP8;hU5
JJNX=c<nXScYNc6FEM7\_eRB92ZC?RmZaJ[2APqXUK>ibLD[DiAg0=cKPXIT6RPn
jdo?f1CEJ\7@E>VjT4Yo887MSIAaRBao^2G<K6XXPmYOPJg_9j5QX6Q0QMdi=7SC
^>Kf\1hdh5pgMeX`>7GT2MFU3l_SOB0;?WXNJg;``eVm95Wmjn1F637=[Y9Ql=nL
a><T9=X3l:BgT1HDFI4DVH0J?Hb;>BCpX\iVZmqf6L6jWJ6@M6fFB>n4JTglY8[_
cgN6C`RdTaKeFo=2V=kVcSZ0SHVeGJNM`eXL[Kjf=96;^I0_YHmVYC`n?q9Pkkj8
;kelRJH>Bq@jFBLNbN3RZX1UTDI1o<iTFLPL@A64>dh9;;X6in_U2=O:h5F2g5nf
:MaG[jPEJY@Zo0ZRj7d[7;0jC:LnqF^YG?IC$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module HA1P(S, C, A, B);
   output S, C;
   input A, B;

//Function Block
`protected
^hYL^SQd5DT^<Qll0EKfLKY]m?gTAh0^N>`pBAb6fUJQSQ^ecPBH3oIW[WOU::57
NGToIN^jUoZYFJO3]Dn61Tj6PVOpQch7XAkNb0>]g[M?g^BCbH^Tq]@iaD2q`TWb
LW;3S44ac=n9Zm6nnA23BMdAhXqXXNcZNi^[S]<O;[k?4H?MG:X?iPj\lpGDO?j9
epA_3GQI30OPWi>26IJ4a8HDoIe06]1P9L3RATl;E4B905@=I>Y4q1j@XV8pAA`4
^1=IE\BX;JcdR;?lMn27ET2f`VfG7]E]oZAD=^8WNFjbDaOM>9>HCWORSi0hmRZA
8DQW??Z9j3e_cKg2C^YBico8H0k6]U9R01?Nb34p4cI2:PjC0;QHbGa]c`QLI]BD
R;V;:Z[WHKFIL97Jf`G3W<>H_6Z:MAd??:;7nYTYBXWoDi04OScAYOomB^VO<U1D
eC`IAjYPS@P@R9fM;_7q<QfmUXm=E\4=eRo9cI`0KRKDR?ci2B01G`Bo7T;DnK?:
mZ@;OmZ=fLPdVcBRj=[U?=F1OGfh4:FVQ]578ojailT^?PCUp<J4Q>?P9RZ:j[P6
a3@BR:2:;LVG4=Rd44]X[LXPM7ZG`S<Uo9:R5icmX\f0SN:J6P>16KMlUg9KJSfl
9bCQOjS`T:i;QQ]5hJeX:XY7pYn\C48`G?gHhMHcne9TH?VZ39\^3c4R:W`[HV8J
UKkO[6UHoc4WXhVX]RT_kF?33b<ke8V6SNgJiU1AIFi8aSF`f1>4\6oaHAmdO8oI
q;nhZidLGU?8?OIkC?=6]?GPD9<7T[1MS:YN\DjdfL[ncc]b`jNYI>NDc0X\n;9L
Q7\:i86N?amCk`]en<2DE8bN7pg4VU46pWa6AE3nI_6M0]YXjacTq^d?g>b?YaDo
>BPQ20ZV9=6kTA2P]239QL^J6nVci<5GU]V9E^Nae8hcZFRfK?RW?^;QV_8[Pg8E
LKXL=W^qo5K8\dl`7hh0?WMiLUZd@WZZ=G^KKi0IZo1nW6R^9aDFJBDcQTM4:dR_
8EE\JnfHo4i5IMGT<KC6iVc=[mpfB52Im=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module HA1S(S, C, A, B);
   output S, C;
   input A, B;

//Function Block
`protected
Zl8F=SQV5DT^<Q`1TRd^>:RlWb2eCb]ScCTEDP@4X\i??ln6qIO9K67T_nTF4S:8
XLb]SoCZnR:bNMK=?VE06p5990GO^[B74EG=YlPL6keW>;E13YQR2f35FLIWi_Qh
l@a@p]m?al2qJ\k_da8\>d4;[DYlCZ5hJi5EgIf:lXq3Y`_UB@4JM;JOLRKA7_f^
lPi_Kh\U1qac`EYfjqlAMgYmqOca1\NeY>Kc\Yd?7l7cU065d_69nh68ECh`6`5@
C_0F\k:Ll<7:n];;maObk8Z28=e48:?ff:ilj[3S_4@OH9JGn];4[DGVjD_`66M9
pTD8n16@]@`H7<Al@YLXV]b<VY^^be43;2D69<^VJJUb36kl9gkfkLBTQ<D=:Zaa
=lMAQJoZXM9>]O7W94ReLT7?Q3MXH`19NbF1iOG\TGC=qfkM5PlTLK7HEo7a]FLi
dokGgK5L;>[_jNBF6[<E5SXAOSLmZFKoV@4cg@GJI3Ye3OcV7nGW\ahj5CCHJDHe
\Lic:9UklpbE<CQoO6\:\4YhHMReNfRLPfncO=Gc?en\^Q<j5V^6:J`2g[=m?<?^
1MCPhfle4GbX6QcAM_d]?VmB0Hj[Q>>JY5Fm6k\L?d:>lp11CfHKDQUZeV`\IP56
lYa70mU>G^D[>q38e^l89[bD;QMi?;EKl=F1aNgM7=]SemhdMgfe\4Qg_GgbUe\n
8o_SUXJ6U3d59o35]eZJiWNje`AeUdja`Y6SV79A3V4MemTdJpKa4>EaYOk<93fm
=[=Ii\0O:TP][^jn:_9flAm4adoaT3Kg8KWG;^DaWM<ag5aog=KZei_@T;3F`Th_
L?0JMCqWlfda2qHSl@O0c5F?7M0O5S^A6:4F<oB36IHHhA[:N7kcV;IT>NX_hd_U
71\VeOm^6Q2eg7H:1]D9=9SVH2D=;=TDqeZVjAj_bYaZIGD@m[64`P\b8?C1I]VV
RCDYne8>QhX7d5\P=Zce`>f=h?aUfnfD[qWUQCUMU<9>?^LP2Ca:9eRo;BWU2JBN
5CP8i6M=1L6=8PWM0mh;S>dE<R\_Ka:B`9W<eLj`Y8mLLMbfCEo^qK9o?^U3$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module HA1T(S, C, A, B);
   output S, C;
   input A, B;

//Function Block
`protected
MaGC3SQV5DT^<<7bPN[aa>T6WL[oBj`Y`nXX0QZKDU[jF5?FIk8GfjoQGBPYVop2
i>aHCa]cb`0hTgo60]8lGQCocIEF^_NV8S4\O9`KegQg7\RW?GaLJob1YW50<qn>
[SD^WaG=jl^ZkeYmBl6dBjTU9Kb7d0aQqI]>ggTqP<ck@[oT;<W=i[`8RmmF>jY2
8BY`60pLUCcSDHEd@e_Jj6RNZc6iEcK0_]D0dq]kMhjkapKgE3F0pC@5_[W0kmol
1BkXgIZ=cSZRNAR@EojK_WK`A?OhNLO=EIP`:5iO3\PM]OT0@UQh]KJMGnBAi=e0
;WTfeQ9V5XbXQ23g@gH3RB3gS^`[b^JgpA2g7UAGj3lg;EJ_eb;bHG`NOn7?gha7
61`b03]n9HAXCO>aEA4=:aHgOjAQDCLeZfZ8Ga]]>VkAWgQhKTXglobU86EhTQ<D
mWf8=S>Y>fB1q=?EY_ZEhEoL1eLVChi\L[KbBSNIX>B9b\kQ<TUBB2URFL^I`J@M
okA5ndC78275Jd1a<:A4a\<_cY>;8=ncF9d9l<eECpoAWP4Z?g7U6;[iIb72<f0<
EWSkjjgR[1;@Je:L<[kD;5@OjjqXXI7CDm3XJ40D0f5o36jgJK5W4XMjRW35:mM5
^OXiha?Bl5gNhE<0\<`YJT9S0Yk8]jjA9<4[UMfG1=[oXU7F[HadcBDQ0lUR`\@S
W18:egp`ZHZU>MZkHFiD]:A2hlZ1>:6oaQa=mUAj[`?387kD=mTocm`L;kgaNOei
PG0Qo;mUaIY16nk]]4@fZomae_Qn\HSI`k]M[ORF72cT3m@`B^pR=1GlJ`eU]lDC
\>ll_m\Yg<oAFa]W\2iZ;cmXc2@^XGleR7ET8MGgG6@QAZlEI<:TDWFBhTN6bl5V
71Zh7caMkPF3DWoq46?7L4ePY@\9W48VY`pAZ<AFbq`=W2Kih;JU2X`Z;MZj@;?_
XFJWN^V>;L5i=UKm0f>C3e]An3k0YN]:c22Y@kHk8>`;k]3T7c^O?73INUl7q0iQ
edQonH26in3gP7XFjKNQoR:\\3F_@a[g]@ZMlCcl51@AfBOQO70[VNX?oc4jf0Od
ccEb0nVe]9>8UdIpO]>H69[$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module HA2(S, C, A, B);
   output S, C;
   input A, B;

//Function Block
`protected
EFLi[SQd5DT^<Xdh5k8m\DOkSaIBmO50<_XHBIENOm?l>NYJNU<ND?MRD]LZUAg`
4RUkiD0E_KKlpQ2KCHK<>193^85><X7EHW`5462SL2V]P[N60=<>3HlFiY=KmLR^
;bNTQS8;n]01ga^a8p^X?fC`XX82Q2FaBEc9Y;1BSDk3[M0fhphK<0?>pi<bN::q
RR>SdJdG6HeZmeKDP@E6]E:@oSqTZJVRRaRMY:?EdTAc0pXhA0SlpUDXKiC?dACC
HX:9D`LFYc;S09O]cV:nqGbdWV2:a8IbL3>_RSG8Y:^<0hgQcfc>phE@]TiGq^Cd
7ZBpS6FOSe<f2I>OSVohmIT[WebJ`^kIFMIkRBjIDAm8`hngo2hk17_Cj9V`JVnJ
<hX1kPGgb5AWNkI53iJd^1K^m9[BWIWGAW]`f5\5G53No=;pTUo:6XkmnVlPlle0
g?gg=2EW=h2J_@UIhmiaRmJ9RQ@7:PV3G?VW:HiYnE648QZdMo3kq_\=14P^YK33
2jnPMb1S_8G8;]4M;cO``[oB^OEF3Yfk`o6cgCSS<6K?j4fPX0aRnQVM3iYnAX?S
K]iVZ?n]Ad:Uj<FhP`1HnRVCQR?ZkCdOqaCRJP<;]`]n_ZePTD3W\oo>LH;Q3=97
dKFPGWBINSOZXI9lFnNgCZOg133J32>7I1YT^8[YYB0oJQeS4Qh`C>Yb==i_jp>^
5Rl\Pbn]SHN36bb2`6FJBS`5_BRJgLGgThho7\BNbV[WmaLJNniEjL6a6`0O:Y>c
4RFoWI^NWnWe]UmeLn<;GUm_8nFJgClF8qSiD;<:gToVI]U=VjX4Kk02l9T57Obi
oS1?YiAA^<Ab?ISI71ek3DABi0l:\GD0aoS;<iU]>nY\c\k27T0\@6C102kQo\Lc
o1A3;pMZC4l23GE>F;OP?HS3]fQI`08B<51UejW@FFXcR3?;JUL_GdlOd:ee]Me9
9XbFToM8JQ3bEZPF;jIe1AH7DhpgNKkL?qaL0D7[L:`=mV;1eLBKenZgS7?_E1_8
g>jTW=GUFe1g:VgNiY<o7DNH]69VEWKO^PP6a5MSB6GE>PS^2<BCc2D^pUP`FdTi
`==MTKifj40?C@:ACW47dG4aanC=S:a6_?[38K1\_j5PB9dQ@M:gdj2ODXPqEmCg
GE[J\\XBflG[WU]9C;JLZ;XFB7kcjbdOa>faCIWBADGTLlkh36B:IWeBj<DjEREI
0jTee]bZYeNcL=qC9j]nn:$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module HA2P(S, C, A, B);
   output S, C;
   input A, B;

//Function Block
`protected
O;:10SQV5DT^<45aB?ONh7daB5jg5=qGldGAc]6n:2JWChgMF@UN72b:nQ4d_MKb
oKf3\?m^T:DgK;\HaECpWnd<Ja@8486MP@V9BFB:R1T@<^B9I`p;4Q64OqF:D9?6
paS1B[J4`TcoeU522K_ee@a584HpCWh[9Lq5n=k6TZ_X4BJK^QbX_n5R[Tb4Z<a_
b9]ncf2dIOqce]j7MAl_7eThl]jh2cVQ\5=[GZR`aIp=SW:\7>;78gjmN\]E=iR3
f6L2JGWO94qh><I?Q4qGX1c\lq;bIhjin:VBQ3S5l[eA`L4OWD`K405a3;SBOZAf
:U=:LYPhUhjO<\Y7b<UYo1YfPPODk5XL`g4Q=@PCWETlBfC>o>h`AQKmWZ<b^6MJ
n;5f7pZ5aHj6O=@PG5MiN63oEZI\K@52;CDa@IdjGBNQTmZZQ@NekL=YWW:Sc:hB
6DOWaRW5CK=WJLQK>Tn<QC;BQX]g?iA>PZc6@2FKM@TlA;9h9qhWni25\4ij[6E8
c[nS_n?`3fLGM1QILDF043>9Q\<PCPc[3GM\jj]YVcWHh]:iIgB9\Tfd;kY8@_jR
ZZIFR^TjbEY]d:qU516@WWW]4L=_=B8AG78?GXg1KCICWJKeLW3A>ojgk3AWLYg[
dLIJ_DEc32W@F3HUN^h0Z9V@_cQ;6@i`XHdKZ4TDPO89nJ]SDhqb5n:2QehIiCbM
HYnJFhfOUZUKM0JZI`0bM8NUKkj0Q3m5BoLM1;6ZX32<Xi7A:OS=FZ^qPekcRAS\
Y`3g_F6Q^P_@9fF0C`<3I6mF;Z6l2VG`H?5Q^o?1NQE^M8STH^3U4>6\P5Aj8:nn
O\j?^]BoMYgfanCQLG@OKgmA086q3J?oE[V5BSC8TKZ]\YimN8Bhcb30;fSg_E];
7oXO:n7]Kc[AOFnSdK@LGnO8gKM>3n1ghH7IcOEnB6f]__2EpB^b8O1qUN68AiOc
JQEoVV:bE88lT;<hOlmK3aI4:eFKj34k?:a_8nicbZW6N4>X;FkZ]aP7L`JVnV??
g?hh_[FJOX;A`DkAdBpHjb]5VQXFN7nN?5acfO:EPG4Hc:WTd:;\5AaDmYhcS8U]
8?=g<hhQ7B:;oIUOS;:Hk4cebj7C^XOlMKE^?qUW\@K:L$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module HA2T(S, C, A, B);
   output S, C;
   input A, B;

//Function Block
`protected
>\WhYSQ:5DT^<EeY;NdWP=fWgPh7alNVAAJHIdP5aNoqUU>EgMZFMZB;Xo<RUO?T
<]XMV1An^7;Ljc0peVXjU2CA;6<6Ij87k=916_<DF5p`6CejRp2]UK7?qI[8i9bB
cQ_V_WBDo57;3:Ih@=:pVob?AG@^W7ao9BEOfR<S=YFYI[MRkJD]2H7Bc[Wc_ZDI
2ATqlAMgYmp3GI_JeN1@fJlT8[>6LER0H`<9nB4;4@p:P3R@2\5[hniIbRD>\2gA
mTaCE:j629pBZn3AYopfJ7FcXplXVR`Q0NBooa5Min][SSk2CLPbh`HW_3Og7`CS
g3J>J=RT=?X;W]0UOY@?:k0:?6eCBbdLFm=jYVIMW^]YCoVlko]EWO3N>RiWC@Nh
W7hATpLS:9h63C<S]A`O;=0KAN2FHWbj]T6TJ83>m?^F_DH\`Z^;6K;LMSdaR6]:
bWCdR0qXi0Y`<9H5\W@mkXOARTW3jBaFAiH^0JOlAAP<WDid0@cE9VgO;B6bPK@G
LmmOU_2PV5dW9GB>Bk>lQEdXR457100XjmKl1b8B=L;jYI48GLpiKbVBiIIieZ8W
02SJJaNn8[<>oPFBH0:5gK<I>>^<^DEW8C<RiK6oRY^V0oE<h`2:nA_;F2ehm?0b
0flZj]4YbTA;8>]qkUB7dEL0eNMAXTA@<OZmo7c^TMfPeoZ<CTXofE4TR8ZjbVTb
flLM9nB^eYM7Tk]NFC?Yn>33=37G20@AS2dSF=ilTG7Jlj_O0U6\DfSpVRY\KQ\A
[@8k<O:_;]1:8GfLjfYC9ce5_5CaUVH8k0_a_8l32;FL8]T[GkQbVTPSkgEG]jK1
m;in`Hd2IPBCTGeLcD3]=J^:4kCb10Up8<BgfPd6;4B:kM;n_\TPTcg=FZGWJdTD
]2h3B?[>i:kmNHS0YLMF?4j;6YB@68oKOKXin5c`RZ_GQb0CVce3[je7qJV=2Ymp
W9ECPXU4cOVL8cR8\PG`o;cML>;PkmdIkZaV>VWSgB__`d[oZe^gTJH99]aeifjK
EXJgS:FjB0gMi<P>MR6[XL08S<pWbAH_H\HUhM`80miU8dnU65D5fbo1k=]X5Q^4
HSmk\m2S;:\=MfIgODOaHkAfoY2Wk[UL^]TFTLo<gU;i`qmIc\_2C$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module HA3(S, C, A, B);
   output S, C;
   input A, B;

//Function Block
`protected
WA5aESQH5DT^<;dMFMW@k2Mgj1jWf=[RTc@4c9@RlXl^damgWe<f4k;=qDIZbe8N
@ON;cDX9gdZ1FR2pYo:DW2\gUaam6PL<kgS^P3AT1?XbE6CAeEDiIX;MWfl[:aEk
?Jh3O]G4JEF_Uo5oVeCd^=b8pWf7D:?p;Gme:?q1i:g\^>dh@BlaCigj2ha_iObc
JUS:?q4c1MH<N3EU@g]7@\e4=Z_1Wok5mY^4fq9b^SMVB@;N_LWfPaT462JF4=Yg
TRMc:E>fARKVd2W_>0pc<J4jmpAd]IoS<80gYjPg15:da^lgJ@G=pYKOW`7q4YiM
TDfqa5;:P1pVEQPUBULZVHfVE`FFJXaVbH8IakOOLT3p1C>chC5H>AY20TcmWfFK
7noePR57iI8lKbZ>M<9F1bRRe4T9LloaOiKIiWQ?binT1ELPmDRm3NJ^`LO=e5NK
=lD001<:d589YCJpZ42`E_j7QF[>@cDX[7jb>l9>=nY4KE>RjT:68PiW@77[DjRW
M@jI1l14[eP7NA`8_dZnKJ1\dhGd<4hQf3FdHc3RAgM^:=n3RJhIb7@gQIbpcPlc
9>JP1;n0`In[GPLV3gh1@ERV@AVEL4m?Hj<oFDQOIoX\6kgXn5;IU[3>EWo?>3dj
c==jR=o<US`8XUR5Db?n]h51pmPHkM15aPDHE<I6adRB^VfEokCTGM7?YO[5fQG@
hoif?PRSb8A8_5<;@ADP;J\9Smm]K^@MP7cMjK2RmEDo9Sf8<W\lYGe?44_Xp`0b
4kJ?]7oZ>4_7\=cWJ?P7XLfEgnTTJT]iUg^li4BMll\DO]DRB>16fF;315^nJ`=X
eE>AGOe<Ho\]>^L:<9HJhIPmg@BT;??^qB^0;hI15h_3OL[m4BObFOEmR6NhXZ10
QR7F6dn]JUJOHPeXHOINgU1hI`?T[>LJMB0R8oU`Wak:eagYZjBfNqUM1\?>p_ZZ
RmYE@I_hlgA3hQ?bf>Ik2doH_YAD]6CLdh\cR\Y?HCRATN]@ch78[WJ]B2P>g_aP
LQONTMCDKLYnYF1p:kFeM_A4fFMD=KEdZiQdPOm^dBGmkUMDnAX5G^fFiol9C8X=
aR4\LFFlcXX68]`S:0X>PC\nl[mkj_T77JqFFT30RMROg>YfeXJ]9XBjd\QR[mBe
8\`6VeV8IOm_dI8VaNkM[p>IWW4_Q$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module HA3P(S, C, A, B);
   output S, C;
   input A, B;

//Function Block
`protected
B7;8=SQV5DT^<LQhUYd:i];:he6jGZdIX6:LNahP:aEYbT>e^Q48M:f\RC2S7<En
^aUI\Aq:UbRd4H<J:H\J8nh<P<Y]_4CWA3akOZ>G^cIQ:VJbid><fKYOlT=aN5?L
hKNo99WFomBqh;@0hel3A<M5SbCh_LH9K@1`:GLjlh>bD9gh68p5ASngHqC]hFF^
p][beMI0U2eQM7c;6NknBX_jXjSJn5mpCDg:_VbBcHU\Sj6^`V5nJS@R@;K`C[hp
mlDWZBqce>T0MoHa]g:HE6FT:<>IOhBVmpga9ch[CYi8m7bLZ1Llj;E2JSMUcqX<
QoX1p>U5\SEfqj`4KZPqHj3;V\4IIOC1[J;c7l2D1LXagf6<NEhVUFGeo930OM^6
SOL3eCPIkinm[:>Wi<EPB?X\@Vg<?N_m]7]M3g[3N189MBNV9W:PRC[AcfQg2ibq
dIl:_O5I>dg[@cV;_4CP0nYYWAfnJNnmNPl_HT:S[@3JK2<AadB1TchkjGXnm>[5
53MjPVLJZ3m?57KJ0RGC`@bm<XEWMb\1YQJ]O?mnTV<pE4;kHc>>gHQ@I=Z1Wb7@
0be<dnaMO2_b;OPiGQ=7QN\3SPeb0jZ>WSTjYjd:bJ3H;I8?NWI:IJmhG:J<i6V]
D0C:nWn3p^TLW]_a>Q=ei?P;BBo\X>fS?TQBE`T0kQR60H>N9N8c=WiC^KE<K3Y_
RE3<B11ZXXC:A`0B0fi_[6AY]KXclM^_ZL4WQQ`dPna6UUn\p?3HSE_KNdoenE<A
[n]h_dan@]eBf5AS304blK98mjSXBU4K23C^_9H;nhc`\h=hoQ>@^5Gc4pcHdckR
P40fUWac1R1n]A`MWRXUH@mIX:@^3a[Y4]TU:P77IQMKkc3DblA>Km9H>g5?_A0g
14\Ya]TWP]>:em14U:lFQZ=JE2^GL^14Fp:ZAW<@6`:`YjDh0mNfF:^MmdC7Sa[4
_F<UQ=H5@dKl68ePfL=;N1[UQnjkm^=IiTa_jONheJo0dWUDC]jmS?bT]4q0VZAC
Sp@W79Y0`9E98b68YijScOO?Bg=FlS:Gfo[DXKA0[m\AGia=kP=QIbS9K5dUb6e<
5J@OVDaofk=Q34A?@J>WqNbX:hB9IL]69OJilcW;ATARKanTLN?e<3SGiJWDR6D7
<TD1W[N5]Q2FN26ohU4M5NU`F:<boOM>hJQDYQDqI]ETdN:$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module HA3T(S, C, A, B);
   output S, C;
   input A, B;

//Function Block
`protected
No6U3SQV5DT^<X7XL^OdY\e9pbVUHkEA3[CTD@8bQmK\Rb\ZR7QMn4KA60VdjL?_
n66_oe2543JO@UKKI\_PWQ_?RihPpEAcNm<oYAT4o8>DmMMbEM1Z]Q;ESkleq;RZ
:91qDhl?C1p4acYLN]f4iAidlno[kU2?h@g0dEEX1pYLko[1>U0BcO1hZH5:WllT
kAV78Q\YTqa`S>=RN<G<P<fmFa`oPMY53nS77qo;Gn4?p57]>J]HNbBjEL]QJ?c>
YINRLdCp6<cg7Xq3M?N9]hq5LjJLWpIN:IIM?8c:gk\N<=:kbcaVB>flEEb@J57M
M6hbLS0DXN<Hp4I:AjQ<F5BFL?dRVSKZ?;cRYJo[^0Om=okWji=C@3nj1X1_X4O1
GR_:MA8a9C1Vh\PLh;?e0AY7PYjP[jJlST_\3@Z7[3;F^Ln<mW;8GOY0q[8J;;\0
o4nf<=b?3;o1bA;DM[bYa:aVV3aQ84?C?Cf`cX@o=16IVC[VBgT>V4KF@_flg[:O
kLGHWJm9TMaQ>OSnkB`g4:>LQ=O1c18m=h=;q;l<9>P2E:038d2l^QV7Ho]n3RjG
_:VbaLdEj1O4\1idPBKO\JZP>IN=U58;]52ZoG23XWoIh>@?7`T2;^Ym2nmS:R\^
\p0:[GQMc7hmhhGd7?llf`Qe_nU`j:3gaV9]\eYnZ:NN`f78\i`8hN>:@BKlWHDn
cjJL7GVRNcfSLG?4P^WhLhShLI__?`mJSH]W\_Xl2qARhhFQYN6HI5O?niO@ZNDV
3LBf2_VH1f9`T8i^R@2ffHe;TJi\8Zi0WYNmZEADl9Eg=mCgdeg2emBi83=?We^F
XWMAigaKaie[8DL=B;5Y>pX`DHRjd5i<omX]]<dLYcg]`8@J]Vo>l0@4\N:<h>K2
e_gkfZBWbUnV0T_DJKV]325?_mj\iPSMF]OJUKJ5l6<Xd?X1H>q4F^L0G_dSPBlf
4K4S=hM7`BoVH@qRTQF?>qkEOmEAWC^;hD`XW>JFXVD[kHAO5E@Q6SA<jn6T9ANj
dL3W8go[Q76MWVI]B[3812kENQjJ`9TW9KPBoGd1pDJ>@2CND8]ln5`PQ1mE688O
aE:H48:l`X0Jabf2mOhKCjC[Aa\ldO<N<joK]IX32DAV0jC^JaC3Xl\2<[Xql0LW
_@2$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV1(O, I);
   output O;
   input I;

//Function Block
`protected
X8@IWSQH5DT^<^T]I?aamkbiiDPg<Vj[3F71SPqLPh\60QY:XK;;HFX2cgq`K:5Q
b2lkEh>blIYT6Sf^5`=JE\>DijOU`[\1<oBEWb9e<NOQU\iD6`9pdYbciSpR_6eZ
O^PGAJPF7:XSPXP>N7bqYI5ckabq`bA\HmqU4@KG0giiiiKAj1TFXmAJeHKf24ck
X9kXVHZL]W8aZEUJQde8BYkTBe0?2OLd1ioUb2HZaQ0Q:WiYJ=T?mq]9dMKLg$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV12(O, I);
   output O;
   input I;

//Function Block
`protected
OOa3JSQd5DT^<:FH5YVm7fPhKTfM1R3WlFUa]PkI<]B7>YV;kh4qV1`eGfbfH;:d
InUM6`a8\j3W7e0VYdWHmP_CIHh>WnQ3\CJ?Z<D=qD`JZlgFRf9Q4<>L:G4^6VEK
9DARP:1LhpifggD=q\[>6Qb]76Wk]\ahm2NIKhZ71q<\][S?ApE4fcJ:p2B=\jfd
Z:2jgZP5G]XakCg;\O?M:3HdM]31<j190<XWckjT7=jARS38D_C9V?6\j2`9Z`A`
:`O_55^aW=lqU0N;Nkg$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV12CK(O, I);
   output O;
   input I;

//Function Block
`protected
e26>ZSQ:5DT^<0Z1M_lbJ93eVjcS^<UTA14_[O^`V95Cmc43R5lgEHV0RbMB77:D
q`AlVIogE6fWKQJqlbFGE^LjAG4fZjT<;?DTOJ`PlHY7o>5;Dcb`EhPfXa5g>8@=
Kj4Eja6BN\9:YFf0Ta?lq0nM>i`qBm5Sd`>j:>F13X^KA@RGi4e=qVDHC5:8pT8h
=CHpXNnQNN8UB0nXH7gkQlh:Y]>3ZgZ0KSSJ7J29J53^S;db4IGMhf]8[U4AU2;B
VOI5XLn6d:1a>OFMYHgT`Sp;?UFHPS$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV1CK(O, I);
   output O;
   input I;

//Function Block
`protected
h2Ue3SQd5DT^<;X:F0MVdLYNSfJ3ISaT:[C`IPVKgi6o@4WWOV`35`Ea0KE\SS@6
7d;LPjF8B;\kif8pWXTbeI;P@l33ni8NSN1qMeK=8HfIWKm;d]mRq48O??6qTJ\>
k;G1F\lZ`JHfI?_NT_T2qlAM>:h<qWIMB`bJH?U=FmY<E;LIJT8Tm@ePq>73fGXq
@gQi37T6]=JhGhWFln4[;JALfNYTX`a\Kcb4YC=g>F>=nj?NJn1a=g`;12_`ibo5
@O^9Uo=?HdVoK_PCd?q_dMZ;5h$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV1S(O, I);
   output O;
   input I;

//Function Block
`protected
dl^@ASQV5DT^<X51NLkS[JP_>UlQRga9pNAUTOY0iO\1J74CFD04X733^6EWkF`[
5d2b?6;g6P>kLmVp<`lT7HZ2_Pfh5d6ALe4C]3J[nW\YCG`RI0n6cSPk1BqV]:2E
nq:2HD^BTSfZ_3iONlJE`Z8PZ9pH34>UFEqY4913`q>AacAhYF]nn3m=e7SmdSRl
:ac0faSVVmZf;4N6Q\k7307ATTP4ZFV=jRRf5Rg3FW>GP[IUh<aC5Sg[X:o^qkZ;
L[DgPXdf?o<p2Fd806T$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV2(O, I);
   output O;
   input I;

//Function Block
`protected
jWS:dSQ:5DT^<;n]7P:Xclb1j]0Ynod^Caa>dC\ETS=m]Iqb_@[joaNoKUDElBB_
L6Ia<>nb5fJ[TM9j\VHXa@n4IXIp?di;CP@?9[RId7E^\JbcX8g9:LL>P>1\A3?\
m1Q<`W@`I?Mkc2TV6EWf?6l>Y`96pRYHlh`qQMh?HeKbH@]OH_^lMSI0M\hKp\7f
N`DepeXnn6k]2MfcB94V_^F;k8j71P[ENaP;HdjZT8mB6]R`iZ0m=2YR8Ajil[9Z
0S;0qX702_`pLje<4M<SA\ZTDg6T??CG@=Mg@bGRaY2NaCO]SIl7e9eg;EoXh?_j
Li[BFfT\^6DTLgbdn4jQWEU56JIhS2pVfgG5Uo$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV2CK(O, I);
   output O;
   input I;

//Function Block
`protected
SO1^9SQV5DT^<S4HnXk[9R?U\D4V[_cDW1RQnIM1CH[aL7PA81feCZJ9nk9pI;3\
X1lK3jj>o>``\86@PaaG49c2k20l^m=V4M40jBK7HWp:FOoE36DaFo]R=Up;R@E0
cqS^;h2Mh1OVdY>6nJ42ggTU=CpV:<WfDRp83RWZmp0[61o<aDoZF=1GGGU^P\f8
LRhXT=^InBDljXjaM550TUYDeJ^4LolnR:U999cbO^02LQoO2IMB;@BH7iHmqe@=
V_`@$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV3(O, I);
   output O;
   input I;

//Function Block
`protected
\=R1ZSQV5DT^<lnaePJPfl>GHV5hUP0M6=E`PH=S01N_Tk4Em4X>88C:m<]4]7L9
VJhRJeRnegqe<`j652JU:ALC;9a6E15[JG`p]TVG4aW4KJG^;8Vi?WmUEJL1kP[>
IGBX1NPDS>1mo;_`g2SKm_Vc_S1SHST\0JC>q5ZQ7h`pZZDUj<T^P;LP:e8\cPWg
ABhBqNZ3^BEZqcln=CHpdEWUVG;6a1]^<;jj1dNia4i0J0E5>FN[@OPZS4BVe1H8
PddB<c[WS_SAcCJd<IbIdng^cE^_3JRW\SaUBQqfCb5a^7$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV3CK(O, I);
   output O;
   input I;

//Function Block
`protected
>;n3_SQ:5DT^<k]RdV3>glT:`4apY?BVkZTlE:aF]li]_I:L0]c1a]k;n`dHk=^n
O`fj8Y@[l4CgmBcG8o\q\Eo^NogP6f^K<Jq0B`0Z=poGOao:<mE7nI6?GRV2h1I0
Fbq4kFkBAXpf?6;=0_m6eboKARIaWj>]FcaCm\k0^dXMY9MeW5U;Z=OUoB9OG1Uj
D_D[Z>ecJH]PiWl9BF:pXXk<EXpan>e``PTN>M:WO=oE0ni3?0G\Hck\DTFmcXc@
?bWUUmZP2EKQdRI0m`?4BgoUUCFa6PEEAVBmX:T;[D_F@pfJ8=\dn$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV4(O, I);
   output O;
   input I;

//Function Block
`protected
f;V7USQ:5DT^<64]8gF4A`@RRTbF<n8LmOHnfG0cp5NX2\>QNlT?f[08OcPA[HFh
UL:;EkkCU]iF6i@ZBLZGG5Y@\En@05oRLmE=<i?Beom6VL\kq61W]J1oR`H[7@I4
:?\a=6Z?hmDWHUj9P:6kSBE7paZXM``pNc42DWiYn=;\]eFgBUEbHfWCpNBLfkFV
p@`7W8GqE]<Fj6B\UGRL;nTlIj8d3k6Q8CPf:iom<^30;dIf:cian?NaiR1KcVOR
DcDhCS4oE7\3^GmfVhE\C`d][4qHg>\K`@$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV4CK(O, I);
   output O;
   input I;

//Function Block
`protected
dC\6ISQd5DT^<\ClaHXc18e9ST2lA<PEiNf[P6]U@@if<K8`o;b?76qGYKO6UNA4
hHYN;>2TQfgUG0IVHk03eGIjYkmg\2A<8XolC2LAJ6nW4l89`Vp7AMB_hdok_85D
^E8A=]daYAl9ZB1P9M4L9lI?od^X>1qbMkb_MpMS>=E<;kZnKmgBn]IA7c6@:<pM
3^lWBaqWFcJ8Gp?amo_SN6<o9@9E;6[h2q1ji457Njb;TSW;d[EU0JRWZ`i1ciYM
2]73a1cERa]kBAZm0UnCQeAQdY@XS\\Be>1ZQ4?BbdHiV`TGXi0Wp>27WT0b$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV6(O, I);
   output O;
   input I;

//Function Block
`protected
m0GJWSQ:5DT^<;7XFU^NUTUY8S?[c>fI@dV9[0OaV:GU1ES0PK:b0TVTINO8JKWG
NP>pENVUMWQ4;V6JCAJ==`T=RVFZIj\^3WTpe1oa2?9gMWB;U85hZIWEiJ^aOU[K
A:geWSL_@6TN0o<UfNR6S3NZg0qNN:9bDq^[Jn;_h87kkce=CDl[@UGM>BpM@FJ@
_eq9[;1fGqYUnQVQc1@cDSd47I41H6E0`[CY6[282IfRDJ28eXPXVih=]1g`C=Od
UCE@k`H3`kYS<_^icU59;R1]Qk2QpTUFAk_V$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV6CK(O, I);
   output O;
   input I;

//Function Block
`protected
e`];bSQV5DT^<h=`7mNminpOLo[M`VeOkcl7d;5GIKa_c0EekLmoUZ2oL7<\Hh7k
QZ?o\ODU[o0Z<hhb<N9]eYm[AM;q481OX`X_>;]61M9kaR_kkP<[;S:bNS::E]<;
HW00C4m]h@O`MKmim>gqZbVhamp[WFC6G<n`FNkkb2kEaHH7b7_q4\j_f`Qp5DMB
n>q6Mf9KSH[18^8joaUn>E]__[=cKKi8FSXh^igKO?dTgccKbTXBblVc3I^O4YBQ
;`86]mRKO@KXhiPc:_=;1paQ^K^mj$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV8(O, I);
   output O;
   input I;

//Function Block
`protected
JRYKXSQH5DT^<d1Y;3KgH2mTSogDAh0^d>7qRlNTAgT>EnLoHi2^HaA0pWW[kZRS
ZdJOP05R2g9=ElU]lX4?=M_<?f\@Yi1X81>RchZcHRmjH<<2bhea?fO^<\VRP8>p
?eDXcnpG1YF7e=@7V3X`=7jN:AMS]S?qK:GXlaFqcN@>nDq9dL4Y2E;ZVH:L_o8P
<LWlPDVD055774B3@;\Dl>QT1naYJ3`SLmZFg@S@4aMOJea9<72_CO]1;3k@fU21
7p`k;FPm2$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INV8CK(O, I);
   output O;
   input I;

//Function Block
`protected
j8G5lSQ:5DT^<1LiP]<g6C1ZWh9Fg8d_CQ:e:\?SX\i??h0KqBZRf>ZnU1blLM64
GS207cG57<WSA^D>^4hYelMRIFV7[]a5X^>>4T>:D3EchIlX2@13Uq8cPNf?Z:j4
Z@`BX`G=JFMK@210m9CUX76_iokkT:mlg5hbC[koPhXRZPWnD;^l6GHF_XC4^^q>
]4]^Hqa97C8QDUH5n^`YoG8EYUS2bbqhk4hQ]\pMl>^HBqi2C;5=fY[Unk>aHOW?
kj<=9XZlI]UHeNg1eQ5D2o9018Vj=aLHCo_>j;<kHFGDlRiERQ?4CCiYkdhFUGjd
p_TlJCNh$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INVT1(O, I, E);
   output O;
   input I, E;

//Function Block
`protected
>]aYlSQH5DT^<1GHfkZZ^bVa4kDBZ=h;Y7MQ7QEeXoZ?k5LG7_dHhjo4GB[FKoq_
UHVnGDKm>\;>8`p[AG?ecF92EG4fXnaiLRjD:?fl=c40m=9B?DNdhaX_kR?4Wgec
^q9LjMC1pVfJVGQ[aQVjn9TI1VSo]g?0C>G1\31q2f3gFi5pBG=O``pWAXk7XH`o
C2b60Q_Pg4`TQ8[]@pH3]T^AVeeK4b[W9jQlM\A\IX[28=`Q?iK@RJG:Ma=KJR5V
`f4clk9eF:=VCQNZPhHD_YYihUO@kChE4ZnSp8k1e@5B;d^M^_aNDRheP@59h_Mo
=7l[HH3lNZDflkVe1l7ZDG7Bb[jgKK@8[6Z9kF2G[S`[`LV3U=l8l]7lmG?5]XFa
\?B:TJ`?C[OPc?YFfVSgLME7`[gL3_aWk3HljTJWhE63H2>[WI4L[?bNVEe9[b?o
?Tl^mnE:VI7OhZd`7KofA\J2c62OeP4h:GU56DKkE9Y6qHOa0D_6$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INVT2(O, I, E);
   output O;
   input I, E;

//Function Block
`protected
7CFZkSQd5DT^<8oDaVTbUZEU@V4Z768E7TS<l4aZKb1:BP\i[IPeDPYDT3gWU``]
Y[GdiD0E_^7>pmV7H45a81hTifBQ@AEJ1[Sj9i]PLYi<aEgljX?X\_N[9koIYZPL
Xk@gZHHPEAPnM9;i?qQV2DJTB0NZkBk^qnCiffGpLABc9iA?F?K`i1Cj8ffRF2Tl
26D94`p^OG\4\hpl`6kO1p1BADGe^Y5fakh0pV;mo4_UUm8UW\>dSfW]2GgK7NIB
APK4Z:aYboA`k;IUVeIOgcD?d[QnNQY;01EOoVCfhC6jBbD1=oIRFfWpe`4QVA?4
:la:h:RbE5EBSfmoPk8o`5bX=S18nK\`mNo8oTF^ZA0^YTC:4KN077jnEh`9f6iS
5>S3VV8E2@Qim5mGW2S4XBNde0?Q?LG:jRf9H]XTi^QalbRfD:S4IL]T8<aelAGK
gm5jlQRGnc:ZB?m@bX8\\5AZeeHYTHD1[MRZU6LKf:XK0_L@\:SPUc7UKUW0QA0p
>Lm6Z2Y$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module INVT4(O, I, E);
   output O;
   input I, E;

//Function Block
`protected
VM]dJSQd5DT^<4ilo13TU7daB50VK=p_SbhW@HamhT6^VhC<;jXN2\`J2PQ^T8k?
3IEblIVDUme=Vc4`<8NpbSPI;JJ\<aPH]MaOH?98l4lkJQ`hdg1qL_]9KQq3@j[>
@5@\c5m1=IKk<G;J?RJ:@GN7bqJkcB;NWpImOAVLKgUZkJiFdF1=fHijWdghCWAG
`P5@3Pp\>EDJTq;3K^mN80mm;QJeV4:O9?OOhf4a36SZe_>C`\L1CcIbmabW1LEi
jKS9hf]2FV5HG40B2g1XlU2lJ5Nf;hMDPiCX?;n?q:6i^oA6;Hm4CRAXO=O^Wj=o
<YTmdgRZefY9VOiJ?L:aXX]7HU`>?SHifTk1Zk1ZX:n9]TaPo@5g7iPSlcJiUf5^
IE:8DI=ViUC75Dl1_i^O2So;4oERJO>PNon8dWhm9Bk>JKc:[=[VR3]=oHNbmamX
P\gfWn\\ab52WH:Kid4<Mj[CS:GN]R>Dbi_[]<[Y@@IPI\jj\8DRDV;bq_IV]aEn
$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module JKFN(Q, QB, J, K, CK);
   reg flag; // Notifier flag
   output Q, QB;
   input J, K, CK;
   supply1 vcc;

   wire d_CK, d_J, d_K;

//Function Block
`protected
HAQKESQd5DT^<S0hD@\ni10EKYhdT[TZKdJKIdP5Tfop6CM>4^VGdbX5:LK5Dn6M
l13HL]\NY:KQHoJiaDLAN<Ti<ZP\WKcKeAYBH[Qk`_PD]f7qL3XV<ChEHS::oJkF
D`bfS2N8ODA8Z44]El?Uh8J8QaapIDjCb?pCmO:4WcVCIhecZkK>b`BFHJm1H]LL
Si41jQGc^@G=U?_7`Z63daHdD81i0:IfJ?NkTZVjj210kkTd3dTdHO8kC;pbE<Ce
SXid6R4SF_U1oUoMa3nd4q]:lEbWnlCcBQ5>\o5c2bZ_VRo]=qZTel;NhqGO1;c8
p6iWJdbo]_BJ82bNbZEagn``pTDfPKJFiNIOjcc2l2N95XYMi0j`oE3OFLa5g=P<
m3UEZFdDTCUWY57D4=VG1Y58K3WFd`d;Y4eiR_8UdCG5;2kn?iPS3I\5YZYoE=Q_
>;RH2pn?PB=MTGH5KIOla=gRdin7L]ZEOCZjbUmohSQ6fl:hW:=kU<\QLBbe1gI@
m5Z;3T8f>\M?\;ShDB0mT`cn0mUS[BCT42B^6IO=2c>X?7<ZcglnqTZf99]qT[BP
MQb1Q2bFlNo6U1gULg56LKjIVgJ6ZmGT=Ep7>n6H;OA2n^e8P><nKiJ1ZZbb6CV_
M8NMb1p_IY_T6P9<:LUkW90QCf6P`YV:V=i@kFSP>MOo6q9h@d8IXlO<FNcY<ZVM
EH:c`4AHlM3V?60=2qUWi]=8<:EABQQ?ZKP`eO<l9nb]CNAQdZg]E?_Qk0G6K[Q=
FbIn73IgXZ?1mj;J9]^FM[\\PFlFDmd26a^eDbeMN:;WiA0DWcmPJ]hT3h87RIff
hL16Ig0mCj9eja]NPOpIdb8T;[[kZ@eV1i0=45>99an<g_JRAEKGa1W]hlCBX8Ak
PV1QaloD8TKP]<lnD6XLfbD>el9S:RnTTnDFR`GSJ1_Ha2`f=`?R_ZcG[@kQ`HMS
8Y9^jTGV7Ib=A1l_Uk`piH[el2;G=cOe`;AEDk=cOUInXl[P:g<CJ48oDGaH:ioN
q\0DXSLE=Q<d]U]`Kg=\3I^iNG:_;\jK32LDRG]CfRQ71o>ET^5D<`gCDgVXYUOo
j6[aGaP93Co2=jKDf5Yk9W@]3R5MYO\dLO16CW:E9dVoPQ2ReLEJM468=5RgCZ5`
>pmoHVLXX54`YUB4UJE35QiBoWPYARamlkFLKJF3m;KTFSDQ`oLY;;9iC]jF\Wfh
b1TG7R4e_lkfC<^gL:3>DmmH5]QDC;l2oo:;@elDY\7>7YAc^j4E_2EZk]gaD<PN
C2m0L;qd3SWDlql31Rg`_7\0e3a7`J6>TFW^27Wk8ZRn4nDcUfPi?ZTT@<>N8j;8
df6h;X]S?pOGH3;@PSnDoBE2W5WmmBmE>j@>c272RP9dOWKIp_XdGXRH7eI1QHd3
_I59lSLh5ib;VhMEdYc\U8cpnN08kkF\j3I8;lHBC_7`]^NeCmWHN6n2I5B]3YIi
4@WjD_lY;?<1fL3[Z6^I\kML<3oR\_ZV_Qq:00eLBcW]fY_0PGGWZ^SnkeN^]]mc
;H^Ke02=[JPPSYG3@;TF97jbL8GK[O][Kofe<M:;F1T2Yq:XcZokG$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module JKFRBN(Q, QB, J, K, CK, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input J, K, CK, RB;
   supply1 vcc;

   wire d_CK, d_J, d_K;
   wire d_RB;

//Function Block
`protected
o1I^ISQH5DT^<_`a0]SW_LJ?Af@BcfaXS0=8b3_lo?i]S]GZWe<f4AFHp1`SiTZo
QCaj]58_G:PGT=?4A?J:CRPFDGo4jimk[ZZ1Y[S0GSbB9dLL:BaW20T]TfGGonXp
eim6FAOe\kD8b1OMJkAfbF7GCb@bjo8X:E2D>Zk3ZBOO6QY?V\P=FGi`I_=BR2F]
9\dH>Oqik=ncGqm4FQ`XR<CZha?gf^688\K3YCo[Ni68^glaJR6c8O4Bk^i5`3a^
e;[MLM>\GGmHl^[02ch\^?mH7J;TAF[H8lK7<]pNmZARC>6=ITe49FC[SMlCN3:m
9qSYHdUk9ZJMHSTn0nVT\Q;k:H2><qm_<Tl`SpnMZ6nkqi[;gn;NP1ZEb4ZmXL0;
La;NnN=4A<7FZ6k\fR0OM4AfZQ>F==PMf0OOC@kiZo4<fVQ^kA>JF]hUnQOWCb88
@g7TKD@`_[3_k:8C;>15XESQCq>XLUX<ogWhNjLH4lUJ:4[TKRNZ:`MN`6?I529Q
2U3@V<mWQLqQ<CDh0HTSo]\0TQ:93\0o31]E3?l1L19KAAMTFlYih:U=>\R8;7U4
TSS>@JFiYd=JFj2c`D19:?RmW89amY\5^\kGAV9jdbiYJ]bahM4PiKd=jpLX`lab
ld;1kXK5K<N=>_fP@XV[[ofE\BKM`B]b9416WiYm6GM1eRbiXBCYQGkREfa@4O7F
85ZS<^ib8\gh40BCiD9o0MYS]jg>OGPDBbqJ1hokaj;DkPWSV0XSiBN`nE_[DMlN
I[^B\MXEl\aLCH1M4YM;=FYH80b\l40B9UI`7YaQKEFDBIJ@Vn17n=f>:]SC]?EP
hKX386?=cT?3RpCPRSZ0pcf<]S>V8EE2KdooDhg[\b`p\UYAPIHeEoVC<PkS4cLe
:fC^`jGmTM77Ac^bFBpo3k=K^UHmiWK4;ELH?BYZjI1ibCj30]nk\fp^_^Y>iF74
1RGW=3=?R7T@=U^=f_TgPgKXl8QN1q1a]k<1Yf?431dkaGA>NZQURJX?ikb:0kY]
api;U5<4_Te<nBk[SkH[]4Io0WhbgR@Lq>RI5?YCIO6BZQ8S;V@Ai1o?J^]2BO2Z
OTdgQTCWBH`BPbbiCGU1@gJQCi1R1f>>:WUL^FU54CE]Wb_DR@ee;WM6A[_RTCEg
>C:hZY5f1Y]km:S4BL6UiD;e9^9MM3H:H\@fL2`QUnBj\p8E[V\SZ0Z`ai54V8gQ
5gXhl32@ZZX]h1\mcjMl1ji^2mMGAZoK1[>eKgRmLnIPLWe97>KAbUebUa<?7I8;
MLS7Vg6;JLX9Q4fWBamVMIST0hEaN<6;dNMBfIEkLdJ2OSD>X16AZkql=goSPj8a
1LJL9Z07a928ae1[\IV[2b3``^H0G]I8J\GEZ?NPn1oH<M>WTom=ShVma4c1c4ne
>ML<\Qlg^YQ9K7`IH^ZVAc9NXo7=X[a5\<d\;\F_VUROUWe:PS@Bj3G:I4mcf8b]
Sh@pA<Y@WiceNB3]OldHX]KPU;K=lCP]h?n3eOUSJY?@ICQ3:Ad9_4XHYgGU`8X;
Dm4gQR>Ze;NWVV0984YNbO6T37Xc@?9>]ZNKdW9DC?T`Ua>ilgooJabLUU5WDZKU
6Z1FDBO?0oZS2^E1pMU4YcnqPo?]aimJG7TQ@DeJ1o6P6OD5og`Ce8L07GaPAT`>
i@Sq<OBYal_O4hoLOS1iaJP;<WX>S?B?7;bDJXE[Ad95H1Xq6b0lD=W@1bQZWg@<
Uf]XK:`V:WF\\PoJP33?G7;aYoZ`c>PWiR63ELUN3;0`Y8R9C?;q0MJ2JU39=kO>
VXK\8VemfBaIfhI4nhmGXLTQJ\SQd\4Y]]6^?Zam^2eOZk<>8iMobY1dZ5`kofL8
UR8Y@R9j9cTTVom_2jmnlF\U0CfoIMMbeZ4]igVZbO029[piBImZPqYYZB2kRCJ=
[;HITPPo0FQIQVk[maC<T^PLaABnp7E?iij]Zdi0=;?_@WSh]OdKX=GA1\mdbSE@
egDp3`C4V>_lF@\?oVgiTooH[]Lh@:4A@X_cEYP<^Bp3O]CLZenO^<ZP<Z5N2A5i
I51i=ggSYpH\1GZX8kN8j3i?3R1KoG9f^8Uo1^7h`k]MfFYRVUDZlM^1fK^B;HkW
\d^0;SDGb\L0J;V;gAhnqYN7J_hTVEK6:nLd:4g?^__;S0jg_kY1`Q1V^EeoM2_W
KL6LYf<ll;e;[[P2ePPQGVPOmlXf3>Mp[K59b6YTg7H=SdjD3?c\=`N2k@BT=e]9
7`IA[=AVa77Zi4AK6aO7;P]SB>`JRA\2HE@dEDKSDNpDH_BOLS$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module JKFRBP(Q, QB, J, K, CK, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input J, K, CK, RB;
   supply1 vcc;

   wire d_CK, d_J, d_K;
   wire d_RB;

//Function Block
`protected
eoIAMSQd5DT^<XTagY:TLc=054W0@\d4i]Lag\NJA9B1mKE[Gb5lc:WUk?g<X<E6
^aNIJAp5l`cJ86heiNZ1DL^2>N3o42;2\A0UR4g;Q[3V?kfS]D_8=J7QRUaEON<=
b7q1gAoBUo1lQ`PX8ZomIiRNFeUEdTTM9E:^5V_Pjiboc6Uh1\l03D>n>OOViGlb
X\ZZ7qe]3D^XpNGJ1LoX7GKjk65YG6WYT7\hXj`?5HGikYf:l>Z=_ZFb5?b^]A]k
naR=f1LC8@1aBP3f@eVU9aj\;iLQ>hIYN7BO`qES5iCRBh]o4RO3jj6nEVhXOfA6
qBe]AOJ9k=Wh`Em11MZ[5XIS]79gqiS=`fCEVYSDDR1DFHeAinCSOSG]W2Z20_8:
>:kpb2>PK@2qNUZ\?kp]LbjUR]XWf`HN8:J6UmhOQ<\l^ee_Y_Un8m;[_APH:0FA
lE2=^<eOXPb\L:1l8g5T7o7=4h\4_15Z]?gBLdYZSM`84=1oJlETG7UoWBFWS94p
gnBFkN\LZidY8aY@@Q2MXMjdm^n38SSJK`LakN4CSW5\;`?^`9em?bGl?iF4DUKB
\mkiJ3BC>5bU9\Gb7=_bnaBS47>\;9F6;KSXo9bT:LC`m2p>B`cg@YCoM@o_:oEW
]MEf3?hAOMT9Z\_bACaLMPT=DhoDR<`Y[nPe3]N<7>695JVSgB@`ARd_j4DYbQco
h<K>e`PC3;75n]mOgiEMT>Hq=C25Q_8^UBTJZAL9g:m^D4FN;@@EHHb>hEK@5VcN
d<D9<@ni6QCQJjV0em:lQgEia^V4fZ7DU3oeWA[QNeRY2<E\dHiMJ>^dHXm^fWKh
c>po=Rjc>p\K=a`AoCYML=A>@5K?K\SRNH<ZQgF^h3VSn7fKpW5>1hg5JWgimVkF
HnCRHW\A1AW<@T=2qj4oPHZfN0?DgRPGbYgJFkPo^8K5R_[^=9ElpM;DXDio^M=Q
k:^ZZ\>C;Mbf@3]`P[aoXk=hTIWqS5PIk\?Y0PEE8^Q15EXkGAJiVXBLVonVMLXp
<QXe4jCi6FVDG]lAIkRnIFGMHESB9iK]jXJmLI>0K1I4Z58kX>RAL;66nGk5@3Z8
k_k3RkC8j4AEV@d<]<a;9k1hC?\IBef^OigQfM:OdCklIJbRiGN4;H^3]c83jnJm
Rd0WVF02l3F1pJ@N6C5cF_IOZ:[U7obg:B:`KR[GAJb0K]jJbF?[TXhk`Qc]k1Af
EGWIfAFNF;9Gc23ZU8;jg=UkOdiS5if]jfi8R\V2]`c_Vh>M5MBFBR<5[?TN0GL[
4Ne8\D^I6o4T:R3]k\igBqX@Of\e5KcF1SmVRd`76R;HK?ML:fhoa8L?TW[n9K\b
Ra_jQWk`7kRD:RI\ZC@YnBBBZQJ5fW0@LReh]LWW[iCiGP]Y;Ti=Q653<\cE3Y3I
g`oFE@;D25FeUKUP_dAj^U_8G@\OnnBFn6qK<Z<Fi]>E:G<k[QncaoecUMVR3F6^
nA:?L>mL<Kn<\n5Za<2iiHdHVnAGgQ_OBObVf67QFWp8g6>ZPA2:PJ^4Sb7;f[l6
\G7?:M05O?Uf1\0=VjPT?8mT0^TY9>A0=6=]F<O3k=`8A8j^?b5_HoYGQ9NI3TW`
Snh98::j_gC[dNJQCD]Sd`lR`;e\PBOCjFK8[Q8e>X3LUJ6EYYj]]6WpBhVI4OpK
lk?TK?Q95oO9Th?5Ee<oPKUoIK`XCGca?N\;EdhJN<po7G?h0l0J8NEboincChWU
^Mn`7h3jD_1m1hWN`Z]^bApQL0`OH:k;3b:OEeM]X6=9U7JZ9RoI=9lmEk8^cd^;
Z7T`TJY6<45o_[IFmKP]PESTcQ;\XZ2m;cV=0^n0[S_MD\T>TF4jX2j^gQ<I_?7S
kXdGjdh3U^LXLlNLlpj4>4gdqbR?:]L_jEne9>hF1e]E9a9_6>@Q8n`lhR:1A\Ip
H_EBVJaO<d9]H5nTV?IO=<e`T;dfqD^c9BgnV4o^X?_m[TB;R>>>Qi@mMI_Ol_H5
deVqD02If58>=gLgV?S4g1nNhmb=4b0VS?A6kaXe1JpOD801\5M4>bEga=Imao1R
<\hPK2W9>IN>BKo]i:KgeGo9?l05dS_REXFM4IZQiTXD1RgXoB`fSq\hL7JPoP:G
L>ldEWIK3[R?C@eD:4U@5FCd87^0k[dAkg=k:U8;P]=\4l]o0MfA752Bd;H_5HKa
p`BOJnf\;Ubb<a638Gdk@FLLI8?VP71cmK\XJ>>C31O3\K1AY<Q4FI<50XMBRcCD
LH:2\h0:JV?p4]mi>9c$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module JKZN(Q, QB, J, K, TD, CK, SEL);
   reg flag; // Notifier flag
   output Q, QB;
   input J, K, CK, TD, SEL;
   supply1 vcc;

   wire d_CK, d_J, d_K, d_SEL, d_TD;

//Function Block
`protected
NElDnSQd5DT^<g3:L^OdY]SgqlfCWG[aMo@7`5c:E8Ni2i1JGoC=D>WmWaYoG`7g
:nSYAYmko9oW<2lLQGL;q>^1ie?G0@^0a7RVhCM@DQSqGJn26kp<NVSZHXUE<gjd
kgWi2]^6e:ce]6g:4[]IFeK]9C`^G_RQD`gRCG[;@2_EeMqXm<`[IRNVUZ0mA:0b
U`bF7;]3F]KLXE\Pk5c7IQ33<anbUMGjRfi8<RHS:GjMMgo<fR=:3OOmU8hpRWRD
LTEkJRD;c49A20g_V3g7\Cq\iCR5AY5EICjSl>X4MQV?DlHToVND`5kmcEIeQ2fR
f\8`L:_:_;[`@4@S=O01e1Lj:^]IJpAjVGWDo7Z\h=P0B1Ig@`@\nm5[HqUOaHa7
f8>^;UB96bgomiH\Dj]@;M[>4C]iY:qBQE1X@dVL67nTjdmITEmJ^m2>Ng@Zogb<
V<]qk`GE^1f^FR<jU7If?1l:NoLO9XX\O0L\OPp:bYB1X3b5Jo95>Hh=L327A5@1
Na5Ycpek2M4DQ5WfXc66oYN1Pd[9X0`iB_HdCbPG0fq]Xm5LXLbf1c:@K?C5EC8X
VQ2S^5ZNG?fL4SIT[i_dI4Io6KOei>01gZ>SCNFLfBqY]FDdi@_oSIbC;G:dFFK1
P^]^<=EDGfU5Fcq4L29EempigBWh^pk37KOlA<>[Z>6fQV;c8iA7l]cS=L]>GWbh
XB4HeBRWhBGWO;;SI]27Wq2jRhCGj?niWj[>RUZFPB:n9l=`k?e?P[@]FlQY3`7k
J`91J59NNU37:h89KS>I[9nNF`7]Q\Lg[hgR]?d>f6]VSb8ZaT@5b?mkc;Q_nKnk
ZKqC>Nc>Zjbdedajm1on]19Zj`2V8;lJ2`oaR33AFl\dPdQGPf]JZ[YV8f8:1BN=
@D@;VkZ5e_7eZQj9ZBJ2hl=6g8?Il3Qi@Dfg>A4_YF0AfK:@lq6N71KMqHM8a_jh
h0ha<UeWM8[hn_S1l<[iK94_4ELfNYmqPZ14CC<8i3Wah`h6ER^lV^KI<aDTXX0i
B8Xq:Zk2PTVImQ?n0DIIM9RLeK`eHo4X1imYFS?<Bbp[AaFTeoZoo^`UeAiCj;4E
Wb\E6cAWj]H\LVqc9o^Ac<N?hZ=1V_d3ZfeeN:NQG=U2YmlogaCjh:f<\5=Qj:PH
GeSP>GDIS:do_>10NNop8VcFC[^J5\KQ?hK;;kj7=lFF<Gj]Ee<FL3G:<j5KqGhe
cTP:hS6TlE\`f<o0VVU\L]RlC=Hb`J>9m;f8pd<I[1KJ54Wg?B4kS>FPlFHl;6VM
U@?B`]VoKP]6p<H3\lM^_>1c4ibEKV7hm;gSMGSmg?BHVIQkTqXlS;HDA:AL@_5Z
_C9cm1IBlgO@c9[@7;0ZlN`@YJ@@ILNSU5Jlo@PPMZ4ckWWMX^L8WZ?0oP?Z7:0N
;;KZLVlNYAU3=SgDd^[Z86?h;G02K_bZ_?`_KT^J0XCNb_I;B06NVT0UE3g7f7Zh
0:jDYpVB\8n06X8T:fGVZD?j\^19nQcYcT[NZ]Ne@JeLlbU2m25``JD8F8b[gg]@
:\\T69T\AaO?XUJnEfbl31U6L>kY;gE:cZjUST<cUT^W`<=M<Wl3B=@FHQ\k`>a3
4hAOSa6\\57b]kTUIF8T_?=T\p@>8jQTTCnG?Z=K6QFMaBN[n=VP?4BVZoOA<UQ5
FcB94WTZ^j4XG>5aNiE7lmP@omPZO3ab>5G;nEI<5`a`2E<ANDZ1Z2i4f3IlZ>lJ
m>AUGC?@hoE^@nM4\YX7gkVMnAM9oTR0KaIa=M_@@dRRLq5ekK50DZ4]nNWbK]kf
SF<C?>ecLBLgPO_R1a6Ln`f:0YYVgo41la;X@a_M@DdcJa3FYTY:PE@5F10BjD^^
aQBhmPkjoJoUMCIRH=fM<JFeebR_<SLc=47:^mg_m^^:`0BVnPIeUk64Xk4Rc>Fe
mqOinc]^J2m``;ASqU`MohEkTWX0nUe@9Tf6hc?Q5;27ORXJF7]bU31VGjXc_NNI
=HoY0Cl=QjY2@B3Pja\31:@>nK6eE^0ng06:K`c_3DocRTZCM0i0@99YPiaYV_[g
6Zn8EGNdaXljT[=oeT7V4Xl<QccpSH]7m;cb4Y`S\mbmoo;ejhT<k\RPjB<O>Xf5
3@=[ai5TZgAS@\Z<P[:NNV2JM4P`JmOCoe\[dh6B1?9fm=::kUdiaK<aK6c_>\0i
B?a`4o>OGf3I\=<alMV]4>iNZ@j0J66>Vi<OIDqO:Z8>=9Cc1RYkXP0iC1B?=obe
d=deTdL\=>O2oIOVQF\ciP^?aNIAbe^BolX5PCgOF3O<7JK>4T;57i;;F0j^iK5S
Q:`JioR;_a5LLZ18MbYR\[gFMB1d9:0Z[al_HbPJBhmYR7H2kb8Nb5_ql=FmjY^Z
FJDhR3N<578kFZ<7ZaX^Ki8\Z8YEe6GRH=a[g8_A8X@;^W0D4`QhKgQ\l6EGA[iE
[NJJWLZGodocKTe]MW^ESL4QHe6Y]?>Sgn2OUJY^2L[2];dNEa\^9nMWY57WL7I1
X6N2>O4<qcI2ih7qSZE4n5iN>P[[]>63Sb[RI:Mmn[6c5X4E8^?j:Tp_R=]jWiY3
jS]OK1JJGc5Gc71c5U6\TlMf[c8Qhpg>k\Q1fGnCKDAlk:;PKa=Q77>1oSG5d55J
dYB1pX=kl=h<8;P^9m^9kQTH4OLYFQOQL`RH5K9:S5o5@gd_bbiF@k=odFNEQJTS
3S_IUen^^3mHEDEqGP4D4D?M<CTfcJT5D8EJ7df^Lc8W6@eiF42WUk@amXJe2Gij
If4N[DSK?jhc7Zncg<2TZDS:Caq0VaPSE_P=7QY7c=RABJ=l_[?`5hj>OBT;IqlP
dgIgn$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module JKZRBN(Q, QB, J, K, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input J, K, CK, TD, SEL, RB;
   supply1 vcc;

   wire d_CK, d_J, d_K, d_SEL, d_TD;
   wire d_RB;

//Function Block
`protected
7?E@kSQH5DT^<@CXN8;DSk0dhH>4NVje3F?1VPpULBB_M3o;64<`=\OFnYCikC>O
AH8LZ`H\a`akL@H[fNCdh`\0@687DOfL=E0RHaIT<:XfaqL_OHGm2f>`kYPd<kNQ
3]3T;fGcE@=V`]^@beP1?\9IbN`6WKA;RCVcWYWM>7;mp8`5<J:pKb`lDJY6dL[?
`D:J87:\^9@9hWO8gU;>GZO^nYFQRnCDRXi@DA<>G7Kcklaqlb7Dh`]>V8b4O11l
>;PV=?aKkiCX<a59:]_ZS<=O?4XL9G;2828;hGd[R1Col8Q6[<a9_SDP@3`imIqa
80l?MU?XLVJ:=8jZb\mido`jJqY>CANXPoCf17_2fah4O^`30A=9Tp2XBm6gP::=
E=mi8<EPfF`GIkMViLGo5^<D_op9]97KXGNc0Q[M7gLOnQBRFNLb4b41O0oj];?p
FFd3\b5L8^11A=nJS:WnI7@lM<1MiO3\g^@XU7=lI]ipKYPB2FjAoD^AZQ;DbiNZ
ZWXShmbI\ijAX`pOg@@XgB:V5I:B2i?PG4I7;4<:CT@aBqGH9bX0d_i`7\kblXXR
kVacG0RfZjo7P>6AAIq:dOT;QNLfASLhZ;D5]8=j9>5lI0[_;^6cLeqa\aL6DKqm
FSoVNpQZVKGOiBcM431:]eBO1QLYem7alG7`<e<KDGI][NMGA?^aU[E<RnQCWUI[
5OAm4UO=669o^]j21a6QVh;:7dViWJ@CjXSDk@4fYPOM>h>=``q>;Q[ci9GCg^V2
d:B[=nR1M2dHi_3aHcfZAl6<1a[P;GW;lf`JAl[`Zc6ECMe6ade^QHo4\=`XDbDL
50;PbBM`DdRSM3\2X^fV?1B6>>^JAi;SjqE<_J17FL26Q4>K_DaXle[^EaaRAHMY
C;kQ]b<MYQ5HCQaSk9FQa05?[U\B[<3mjRD`dJ5mHVakc@o9ZYdI>FSc4j:P:;`;
_eE\ge:OE3q00[@<jI@Afl^M5PnTecS^2fE92eJTZDd[?WlMRahn?e7AJZ4XXQBO
QTK=PEqlP7;InS@HI4?gAGV`]FHCm=Bo[mC3RQgM=TS7dTcIY9keJL85>l^0DkGM
`K5aLl>HLTlBkjNA6T^TA8JN_=:7_Zd1AkBAB9P_ZC;C`Zc1:q_J>^;^qfcm;XS9
ha4TOYBmABYSL56]K5e]Rk<>g@XWVj1qC?;;feB8F3Ubo45Ql==fFIDE0UPmH^Jg
FBbq7[EY3=kV>a:oXekLhV@QDV?2SO5ohQOOeCVRfBq[lWPYeaY?WbVSQe;`cHJR
?o>q^d=`ll>ETHhT`cJTf?KgL\EhThN[IZObn6<p1XADP2E^^geA1@>51T_\Fh@a
H^7Kj3`b52ii1EGEql7i;CMh^YSlPoO^A_=@Pa3b;GY[U]`A4<\e`Olpi@SeO:SW
FBC=_RcE`YGJ9<l6hkT[Jbo49a]oB6Ppgan_RIYBQLEg51P;VbeR;dHTKiZ[[TEQ
cHFopNEIF8gcBo:gYjWGJ_=>WG;R8ehAC9]a1n1]A1Nk=AEUo=[IM^d:5KXQCe1N
:7>oGZG8?Od]EB10DoV9@<ZoH`nJ4R<YdfDE921UNNXjOQ6<=Ui90ok6ngfGKHEg
PSMV^NE7C;O\j><b4fSk=S>7FCF@VLdhq=ZYKWSoAaFmR_278ncDaT\4DF[<C\lZ
Q26]`ZOmVK]TCaj[XoIU^1d1RK5e?TkgiWSKk0`Vkf>KK45e1iT[mY0j=60_8N^\
eD_OiIGK8d:`Z3Mlj=f?2^NTOiNFWJU1===i9JdE`QY@=I7`<=5V[FcMi;@`qe@a
XHRT=eSU\gX]N8_aD?]:^YRNDmgT<dW_8mm<jOF5@nWJ:Sg]^mMKh@8VF_@@aH]?
@IJS>@VEiZ\WHh_Wge6T9WYGniU8Dif0jY`VMcHFXS5dXPb]K[6G\ECg?RM\:eR3
0gmWMKDVLI`o2a7O3RJZ1[A;q@^YM;?567_AE7QD^aoDTP:qV5_dUOhdnN8]nGcm
cOdf6Qc;GPeX@XY^SF>mN:GG8BiH^6f6c\n^hcAT]CY<RO]5]1U;ZL?4HT=FSW@J
>PD`hO`aeaC14<L]_YWOonk:39?fNGUO?iO8354aM>hCIdf;V=j@4X=i[[=SUEZ0
gGTca1[1Y9Zq__kcHaSQMdn@_k1f3UBjX>A:XTiLRV5nX4doo_4a^R@6g0@fKPlM
TJOci>_NlLDXjA?McbN\NFdodK2@\Y`IgnQR4i=jNFcnlH1Z?dFDN5ILbXD\C3iB
iY76KfC8fjEV4b3Oe^Mehl]RV_fkB]qA\73AgAHAlgT;elU=biXdodm4]Q;OCX0g
gWmm:3O81IL?W1?=@6BQWPgl3?ZUfILYKnj2gQETPA31mm`<PEVCfR<7D8G;5[>0
nVMAi47UPmSPY>_\BF_hQOQBSScBK<XZmR3J5^Jd4S3]0iGJ=qU;C1FnN_3GJ@_>
k`XggFHUIL^JiQm1K[ZHFF@Ib=l@Ec5c4L`_l?J];kPRF0:<0<Uj?BSokc`XST\o
0N9A;n7aHKRE2]ae<bn@UZl7EaJGa8]h5PE3alZIiUe==9hC_MWmNZm17QkNnnAn
<do:f1f5>hp3=KjUh4:>WnILCjHmO@C1\<QC8AQci0k:TZ2FjaqJ[_LnO<S5mQO_
[JO;CU88`G5d7i^k@2UPFk?M>9e0GOoeXZoBEZEP_>`c<`jYR_<JV0cc2VScbY\M
16YfaRW_c;Ajg78JNao^=FkC56f2^[4QaC1@bS^hG>aQ4o<W01I>2N0;5Ya]k6:;
JlQA0>;L_59qaX^eZhpBVLlDVcEREc>@1MaOKoSbgB3e8PU@hZFZ]FUH:i;h=pdV
PXOnF;]nbiT39NQa9XC]AM8Wo?@cSRCS`gShmE;<dqF6[0n3X824mYL<bEQY\Fhi
I:A44hdJfJeAL:gm]>H;]2c1?59cl@PBMM=U3HDj0alBYf3Dbl7gKW9Q\KhW>o>a
2T9Y@bkamdN:;M7U:;l=l7=[_hohloM\]YMapGO1;cSqbho=`PdIkINHiGNPZEag
dj0qZEBogmkMen10[PiQ1VofD=idZ@WGWZ@hGGdnV]pZAU?PO?Q9aBgX\dhYaIII
WcTb;okOaRmF:UIUQqoF]iY]b54NE>m7OY?K@Aj9LQMfD0YMB97L::FIpgSX1K>\
U;NCNK8MJi;?ZS=_KT?RU\cdcd3mQ@_OnfBFSdOV?K@[RJ>6XW@^VXQl2kn>T@]4
RTdqN>kgIOTnBHZ3SBL?B9;_9ZNk:>\<ESF7d4PnP1ml7T6[O=B^g@[R0YF<@cX1
PfiG94MoS:Eqb0jojL;h^N_=<U`B3HVPC6:[bK]k[mPU6Ajdi^EaidL^hn2og3YL
PR=c6;Eaj]gaa8JW?9g4mlpPR<KHQH04`>\NC0`KdMa[4RJC=T\G1OcINgiElfD:
0ZiNM\fFVBoCmKobjOX`iLDo\bnXQccYhp>[<S4bJ$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module JKZRBP(Q, QB, J, K, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   output Q, QB;
   input J, K, CK, TD, SEL, RB;
   supply1 vcc;

   wire d_CK, d_J, d_K, d_SEL, d_TD;
   wire d_RB;

//Function Block
`protected
76>?ASQ:5DT^<R[MhJGiW=C:L:HQP0W2aPUFXmO;Q3B>>YV;mk4qKf2H4E^VT>VL
V<1YENRZccG:mkBp0m:2T<If101:MkZXW[l1j8ClI`Gikg1fk[?LTBp8@AWngqOW
[bL`]XHe^md3QR6ao>[UM8Vd?i[[TcLRThjg@fGal4[\5=A@^IofmSP7Yp90<]o]
`dkN_i@F\=Vj?9mU3F:bmTAB;0Q?:T^AY>_e>AYcYk:XbY8\eh?Y33<A8KkPYBX0
kOWGDE\^pnS5MJhcjLN:ajA:>j1a7g=6OT1p67^Xd=Qd`aLKHSiD;?IjQlnIW^ap
ajg22Bhk?E@HWf9MG>lY4UnWhajGd9;WiMT\q:@]ePC;F_dJEaj1Znc=Gka^l2SI
0OQ^<G4noqlod3?45Gn`^Xd84LVdCZ^mZY>T?8XMmJ_CpB7K63CYKmd5<BhPRS\0
A>]b2:aYPGUZ^@XqDH[BB]UaZJ:kZlF76gY7B6gZYm]P8CqW<fJhi?d60CYCEM`l
6e3J8UgP[Z_F3FIjaGBqWE\neeI09QSUeC_W?Z=m0GYcIPRFRL1YV9Pq>ebJ=_Np
OJ>ID6q5J=falGg98I]3T0Cdf7iAbC;b6<CWd\jnHL5?WZ_;6FY3C6^8D>JK<bnh
6VP`TlhX5OA2Kmf5X@=15c`Q=QJhRK\?]\\S:fha6fo\;89Ek04q1`[UfR6E@S1j
jNcEUk`3U;bQR5W2^ELcY5fQ8l`me?d5J7:2YdlM`SObhe5CcUgF9GMm[]SolZcX
aO0fF5hSo\<B?@nXGHYGH8IBf_YdaE\lIDpI@4@ST4[XKhQE2afXP?02HKB066on
nE7oX:\D;M0VkX=MZ_@`L9SE<>OpW5>alGEWhoSn95akbK=Sk31M3l_<X\<8fnbL
H2Qi090B_^9F3ib?>BkoC7mMZZhQF5S6oGMgNi2LZ@cmDL>nZ3:H:cD<3;E69BZ4
^jGCpg9]KBV54WS7>AGAM0PPgWo3fCmX<iZS:@=FCZgmgolc6>;CS?Ih><=A6jbP
OSe3oYG7Ce_YN:kG_PGB5T6FFS>^INhFjAVkILl\I=V=eK3pUbb3d^qKPDoNJ0R;
BM;d1<VWeNhi\9Yh=kI[0EKR8:a6aqLTAo]GLG9_1;jW>4h70TONJ2LH[>OHC^kU
Eqm_W?GG1LlcMOmIck9<ZAYE0=H877mGL[dJQ<=Tq`c:nS\nYfaeP7AcW8S>daG>
>TTpJ^4\84BfIBBdGml^nnjgoU@E6ThF2Dlm^<?qhdPmFeR\HKM4[<k^`]MTiE=H
YL96\6UU7[Ua`[Uhp9TLfRQ_JdgMES_:AB`0gXo9U0lFQmMj24P6:<<p>Gcj\OVY
Ei<@\C7lXcfH7F3kE154TcVMj6bODE0pchf0I24;3o1BGBUX56kZ`om2>C;3K[BC
mPhGqffY2a`SPC53`>\l;R`if=Bbig_<8h8gP>m2@FkaH31;eiMJFDeU?4cRVm_F
j?XbRc976B^[nL[hlD=F3e1[DYPFG7KPDFSRE?mg8^oQe:]nnEZYTa;3k^k1S]S>
=Q\:nf^H>eM2Pdog[Ia\FO@j>eRXQOQXpaGGRST:1oMgZVi_DLf8hD>E`EbfhG17
<U;g1YbGjeTe7UAc[k7nRSU^d3aPLTK\Mj03N^QK;;;lB9Llc0EJAFJc2l[m^D=K
3Y:9<\\5Q4=`9>jTNcSZ;_UbL:_I8R1F^aGHkGaF6Yh9o?^T6c9M>IibO8GBqXea
@279jnY412G0i>?o>GBFm^<qGEY5j`<e0<GCZYjEi6;^:i6oM]7OB<FN9d8JbUec
S;L9[6>jgJ=[M]OB__32_d5]hMn[7j`EA3SOLaN7`@RJ1D@ST?XfGCL3<CELkg`o
403M?:D^b47h4`[5Ad]b\CDTGZFWZlA^<_RIX[fhHWb?4N5AZi]qh@hh\cH9QOXW
o\B;c?1OMU1g\eV[:PTGIg0:2:e_2MZm5oGdQXiPOSBVPokP80Qoi^dC4?n4e[do
SMY^gg02SBYleWIXIoH8Lmce[ej=^3OE42XDZRnHTV>4Xfjf8;k@h4?3I?><iO@T
i3nIlB3m:cNQF8?qZ\DIQWJBFnFFX=W4UR[b>?<c`HAK<HgEC?8WFoYo7dZ\I1KZ
:0IcHG6VP5f@SB_KTARnT74K?S8N>[Hb5dVZ[1MJH<\h9X:\TRE\nCNhR]NIC0Fb
HHYWJ2F1hCiNI1J3k2US@<^II]3ReoaiZoqO[bVV1>>=5GCg>;EjGQ=K1C=<;ih9
fg^>QGK7oThm\YBE27Z4aE>02UlbBLFd^Y4nWHKCn7=IS=`LJ@_ZZDV[P4T<[iU_
ObZTSAlKf74[8oL^E`QEnWlbVBWTZh@mCYnRca[o2;`UkHIj3e?7Hp[So2EP5>>o
:1C@OE@G\4U97SmDNTdgbfTS]iZR7J]T8=c0\?]?BV\>\P[mOB;m^VqlZF\bIZXG
YO`7nOPbc2I0I=0U_0;PZCd0;Wj`YV4;A?7fW_3G\DlRLD5<]L]D1F;lndhn@JSo
d:`N\?Uc7Al8QiOS5\J_HQX:R9ORQHcLM0oZSWLR<826iXH>8M\94mi[biUdmYF=
@[kGDmn6mPD9To\q\D7bm[YM6l1jPOj\\jF;ZMVM6HEBnRMJ]oca00KFUJkMQ[ME
T^ERPSXLa[o7Qa\9\>Nff6X5Cl<IKndGiSU7?m?[?m86CUe:meF0DS6OcAeMdGZi
SB<n;?7EYbYDC8ji4h?Lofe]0HnLc?8>5@@YfFhNpZd@4k2pEYjJ2\JX^FlZfRTU
Ri]cM3e:LL4@k55XUcf>]O7Ph=q10WeJTnY9P@HeDJolTg:C>fQHQlc10?fl<SWD
SS;?Y:52e4ig<YgVbNf\JMiLSIJ7Z<f]<qGmVW:LEeknd4YWgIG;8I?OSm:NC9;T
:T`Jka@hlc]<Pqj]TeNDLAk=;PTg5Z^bN>9G3g2Vboj5RE@dn:Z_ASjW8]25[<M8
1JJ\Fo10oKR:O8@>;\Vm6^gLggDFGPJABhXU`]mY;[Y@@:WI7gaQEDYjL2?>Hah8
^`i[<ELepO\_<^@pMZn8X]YmCWbBGL6[Kl68YeD69nIKkQJI?gOQ\2q\K=aUAoCE
FLRA>@5K?K\9;H181bcP^hdVSBZgKpEaZ;b]HB_TQ_NH8eK@=cA01n_K9TcXcZS1
1JL7pVToCQ48Z`>?=7964YG:`?k\e5F>Yj>HaHmZg;iANMPW`V5ZX:4LO8HU2X3D
IAL7L]@U9ZM9=\bqSLhOBkF=cdBm]f<mRYE_YIiO^7c`_;\MUiYMOmhb[XD`<kNK
<KZF]01B:5[?hTi5=g2M4^1\7Qqk[AICQmTOKOikU`NcoUgGE<mdJ>eKXUg6VJC1
mO5Wka2YU`m=cn8a13LXAV]LIRo[^nk4eK_kmqk]^1bai_AX@M0L]LB@=54^c50b
UpD7>N2I=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MAO222(O, A1, B1, C1);
   output O;
   input A1, B1, C1;

//Function Block
`protected
VHOWZSQ:5DT^<DUDG]OTSkFQJ50VI>oLN`jQaOlnVFIYX=lYQU]_a4iZRbMB7<WD
qZXRW08`HQnICUH=6bCbe04VGEI_BR4?nadNiPBX@6F4W?1Uj`_`_U6mhYb<CX<l
hoK2pZ7<R?jm9gm:8CMMj\m0Wf:2eIMMf0Mh`ZnZSSURi^ZR05PUPe=SO=l`OcfR
qE`PH:7poWeo[oV;P3>UD5W<keWIWc5Q44g?BDM1RlpenKnR^]X\FO_CNPWlJjF>
J\dS3JnNU0pCUGGK[R;HPQX84\[M]m30P802?Gm:Jlp@b1RJRTYi0UWb<cU:f[cg
@@klOE7VjLJoLai3a6TqY]V\jEIiEW=Ff]URA_?=f;6E79pT0iSQ@K?a6Pg9lOnb
Al`:=0<NQ3DH?>M9fmR<WjLRWip>LO:DnTqZ;gAScqLifKHP6GQMM^kJN1em[APW
n]KHl1OIU`d;KBjQJMTZo8Rn8cioI[lVa5H0PbGC9XP0UTV7:4ehoSJYWZHfS[BP
0a5jc0c?om?]Af8QgYL0?F=3lX^m;jTfR5oepc@]kI;ZZa5@JjV[UD`BmEE1SoY;
iI56Q4iV_`^fnf>U\j:YaJI\TUNAMD12T3>dGc=RjmEA`5FQ>dAT\3OZSBAa7fh^
B1O]WFi=N>BkBF<iTabcFBAU7AGqIcM:DFGFKj]LG`h4=14bcX?<4:diJl2]N[jT
\FkY8G2m6jZB@bl=]UNV@5UV810LIO[@PNflBWf=X464OYfGh?qBhk5T]7XgcETo
66>Y7LUdBQB0JoEhWDa]J4@eXkT7m;[=A6>cTS=>1g<fV[e8nj[B9:QCGXF<bZ2g
EG7Z;1gk]K;e6egCiTLJJlNN3kkNg@oOJhGKXR?3kpB6ci<;:AL877S:Ha?[>mbF
2QA>Cn6XbVR`a\^@LPSoCbNolV[J>U021L9=[_`Q@:BCn29S8@DSC?cPNJkH1R^3
_@PJ;8=GAC8`HMC;icTR26_IZRgMk_W`q=<DWB<0TcR?fj6f5OFCJLDmB>:8:k;T
0_Fgj8@o640S7oMNX_oMBoE^PECl79WU\=MeaG>blEY]flL;JaRT_V2q8G5@OTPd
o<gI2ak]i4ibM\A:PKL2I;iYb7X]KJp>gE0<7d[8[S<L:L>i:G\kUa9gQ:1OR[K<
C7Z?@_FJKY=`VJGV?nVd4^m@CZfEcHk;dSBe;i3>84[Tj^]]oXRU>mjOnHhgA>Vm
lRBI@;4A[e^VM7JDLLW9[eXZ6q;Gl:DL5<;2dm5>@bbl0G=5Pc8aCCG92699l2FV
jJQbX4RThi`8Q]L@R32I_N7B[6Z6:_@2nRA:9KbESiU22o14V\l[OCI;X388mkWV
`Sn:j250aV@^dCeS]MBjpNoKCc87fd7eoM7eGkKQ`j\MLBO9e8F2l1XSH0[lH56f
a2A=7>3>F@BXPBllIMeiYKDc>eWBT>jP>5JMU@82;H_:N]2q83KY:Rpaa2H>EA$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MAO222P(O, A1, B1, C1);
   output O;
   input A1, B1, C1;

//Function Block
`protected
V2n^HSQd5DT^<2KhIFRePNV`FlJa3X@^YM]i>V8^6KY<nm=gSe^PlPEWRWPi0c@5
dcENM4FgB;\kPhWpfPYmE5]KNaW1T=U:nJB;l`[S06pacTBS0ko^:IjZIQB6_GcJ
3XCIXo;76W=eJbI6BoUeblqo?McFLqdcgG<@ePXgD:RULQ\<E_E>Oa9>Cd?IGHV4
qXOl_o@LZ;=VGLoXC[SkS4d4]PYb`El@qOZSoQiRhc?BmW5:[:U`m]2YUZK;:=B`
pVNOGj?`ejIo03T8OXO=2LdgT]YKJY0lRe>WY8SETq03K7929EmkO78nj^e5IMdo
2mAJq>2CY[L[qoZPdkO35ci^LT6XMWD2YGdMMHL`jAQ@0mEcqOJ>ID=pN9>ZHX=?
GV^<NFDCWPj2?MNXD4bNeR=eWbAZXHKJOIZ4DV1lWl?PQfiLPibbVb=_3fjCA1=O
8gMTLeI[gDPR^2h<kKi9K=kMdGD@PHO09U?Z:Z8PYa]PO0O?C`qkO^SiV3:FbVaf
Yf37OFBWRCFD4KZ6F^Dd7EG6ROJY1eihaA?@`S6Y;U4`VcGboQ]n5?i@hUW`LVM:
b\I7VTEmTZQDOmNiITDIK7DXRIAb?;<Q5E:AT:SjLLh9NpHV9M_0P>SRg@V:fQWJ
aC[M;\i1chQTNP66[E`XliibF>MY6BjE9VmLSJ7alhC`3@Rn>U0ZCgbQk6J04klF
gSe1;>C0pR85EoTJR05HnbeRY2a8B]H;g5A\Q[BkZibGZHn_[CH<AlUm4V^]Da2M
l6UYfE]k?R@D=V1oo=hYaPhiB083;bl<?BcL=kO=]4bW`14iLB5;j^1=h@mTQg=q
hc8OZ^B;JNj4I<C`Rf73D[\Y`UUe?SO8MT_Jn:CgI?U<;L[GojPQ;W6n1kf`IQ@Q
G6qW\85PD3;U:<n;b;0`11ghnNYRS8?Ne44n:5@IgdBoF[M@aK>VgTZKgQmQhV95
lF>WhR4]c^Qli?>MQ7=34?<:^@5VE9VMET5K:13c]4VEdTKc?fU`;IF2?p01FX[P
<CET<ioZCe;ooZ3=n6m9@68nP[kaiQ=a\C7M4Q3nU819n\miMC[dI=jd7k0c3f`_
dFNmcAeA7k6;9SIJqHCg=H@ABSeX6bXI[QFinC4Xm`0DTU3;Je`LoVDTDE0?CBii
14;Z>YHeT\V@AiShG\KeL^n8B[h91F9XYVi1WUIUALdF<lBohL>^4DD\ZPVQfH=S
OCO>@19EC2oqdY;^:Xi[k^99Z5;Jc5Y=@aQA5BYRC`07GSmjhEciB;ZiOF542FaW
h97Ci9H95h04GLIOX6KLc7jTfAI49HdCKY2L=F@3^nF14UfFgEZWVkLbJ^@DjGC:
6><f;cp3J?oE[HKB3XIM4_nVDECJAV>456W;H:<CCHV_BlmAE2T9D5W860>UL0E<
>kS9gV^5=nV^Ec9Si_HZ?o7WJU?m`hC3Ypm6G5egMbIPcNSX[:ARA4Dgab:0@<PR
q`VVKOaq6[P?C4U$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MAO222S(O, A1, B1, C1);
   output O;
   input A1, B1, C1;

//Function Block
`protected
d:ZR1SQV5DT^<O`iNa2IWXJJ>UlQRi=9peZMl[YW@F36]`5U=6UCf@2nQpbKjE@b
aLXk6JHQapd8G5YnpJCYTmhBB>=FZ8LgU2_:;ea<Gcg0R<a3aC0p_1NLNg89l:8f
llQfloUc9\MhPiGU>:MpQa^XXISAT78eG4Fjl3gimYHh6iFEkdZ@gEB_]nEcb5M7
iHQoN@K2FM0jLgWkfS_[?>;E093qRlM4Ska@^\WQ<T]_l:4<<o70flNjgQ@q3ER3
[WHkD5o1k<eZC]QbaN]4D3I>:1nf>QAWPe<5pT=L\S3D;IXGTgnL9\Y7?l7bc[Oq
=K;PI>@G[^WQ_?F=G1FABE4T9W0RH9aZCC8ZJFjkJW[DeTTqWN]O5L[qE5j7A`p7
m=O9bT?=3\`h:e:\X8S36:9FFlKUkFfJ:S?5jQ[Gc]aln0IdkIkG2fA4;\LlVgj<
g5`OQ6HQfLc?kh<8aCbo1KFY0\@18Oe87C=IjR\S6gKY0:>Rfd08ioP:5p4_MBe[
QC<7aM0g\=Pjf1g2K>?hHKi3][`i[6L^onN?Z_i>jZ:ka9P[k`P1dJh]2k_L2kQJ
K5ARG`U8G;P9?KeG;0375doNeOTng5Z^0o?doYWG6ii]FAYNP`T=qW7JJj6cQm5B
WJXEeX:?ZVC4?k3>9LZ?OhC=`lTf:?9D854L[EA>le_:B5<[AYW<hF7Rh<jEj\Ei
e`FVia;akak1A3nqhYoGjmPUZn]:3PYG6M^d?2TXZAS0I:m8Jab=e;_TcNDk714A
KSfIY<DH<cH>6W1JFlHSSFSJ_1B7=2HXC;M<[MFD;BX8i1E7@0ke:;oSmO^F;6=4
inh70R`:0WqX;:EGIdRG43JB<KD6TVVNjdLlY8EW[07@_W@7c[jfCAlU`=5?]>:3
BUWBd]ba^QEX87<=4cJ1XVl8RJ^<FS\5XNn0Tm\bb6;L_5NP1bWd;Dn1Wj`fJS;Y
mpK^SYc3V5S9J\blNg_3ciVV:bnd8KMenhWl2k=aFJ;c3LaV\hPN;\jP6ZLUO8c>
_iKgMMWdiBU`UF>YoijQM7o0pb:1`6D:C6KR`22;S>l=7?36aY:X<db>TMM`JHeE
^2aUJhh74Tn@074;Y[UoCaUi2A[b9eHYdmHC_WEiR]McG9BKGSg]f^iT=M29WCeE
[DSXMb[Pj8oD5VjNAa9pk2Zi0:R`oo;EaoZoOHcHFhEA52hMREWkXciq[olJ5XUP
GFEjnR5OT`jlGQ?`8X<<[BZ\<?jRH]O:UC<Fa1?H<dY3J^mNAcSd\::\5JWMXDoS
2AbLU^X_@b9`f7X@H[P=8m2=:\a=W]6VW3HM\]7TBg=;ENQd9lp?VKeSh2Pe];W2
81mebdl^f]=KCo\MK0hE^5cIRK\H=KRFT9BBd`3CK8U;eGeebHBQAP0]aRHUX=Dh
YK2B;RXg[_m\>p`:Yaj9pFCSicoh$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MAO222T(O, A1, B1, C1);
   output O;
   input A1, B1, C1;

//Function Block
`protected
g=Lm1SQ:5DT^<L`K8`7;1lJ<:=MMVo4ROZ19QC\ETSPmJIq]OUknM0hOeHLfEhJ0
KSOPP@E=WO?^n10ACq44Mj[9>M7==6c`VGfjQoOSF8;9FKn3Zhq^94YjRqVKlnlH
@3=VdQ=OAQ46Pn2V?co2=k;5CO2Hpmk^ogQ156^`ZT_cMZiih4IgiL?oTelbp1Nd
0jflBKi?3EA6OI:C[IOb=?`]XX5Gq\3De0[1Q8DmZHRYZOQ1>n_AkoL\ciR<pbbj
Q@a\oOdkIi>V5R^1]741S4RjlnJP7oLDSG<<YpNn[h<<7m@AFXa4Ph\:_T2nU>GO
qLcXF_6np7kUhZ6pcMM^J]hKRo]BU0EjloB<bAMIXGCSDll5PNX<dW;hGoF5MG4U
Blacl2;IiU6[OTE?PG?K=X]e2Nj>aY@8h8c1>L2_=_i:P1Z9`]dVcWkh4NRY\B[c
^eK?hoOS\Iq@=g1:_\RP5CSg[l_651F93HGO7qkUJF[FN<WCHFILEkR3md2lRLE6
`Hhi9OGHaKMd]QoU0cH49maQ6IFL791Q]D\PFc9JL:HIColdbONIP8k\RJGH<o<m
Sli87WiU[lDd>?RT8PL1<j[TF?UD8:3ipEKQKiamCUK1VUm`EZllWmfkh6bT9>5[
fR<efjaaf0oKGRm@[:nX=S<Z^@53]<CPSANKmfQS\i4@HSg]Db[Z\JeX@CnpleZ;
gfPjAjjQ:POFjO5R@S<cO^b\KgTo^35L6>36MFZ1Ldd5LalFiHRn\e8GAIJlYFAR
UF=^b3hhHj^Q36G8e^L:YPFWd:ci`L>el>D6glLlc4F\:<jUWWF?G2p48BlLPb:;
?>eD@Y_KUHG?2887@@@8I:COfO6ca?J<^1gdlUJheHN8UVnd3=H9`f_EXUj6D<B6
kJJdVVMVcgVaQ;fg<hTR:<>JjhoCa?JWQ9YXFeDc9E3LEMVgbqdbPgnSEa;XoP[d
fceC2;5m9h95BScg;b=KC>]K;SCc6BVE7W=72JDc>lklhULYL^_D0HR956[ma7W2
HFRJKY>N:G1`p2d=TXE?@hNa`?kiO>ggd:^68SD[_D^7I^e@?>TjEnTMhMc0[J>`
q4>?b4Y9HBQd:bMJg>V<h5F\D0YbWQWT?]B_kgbDF[2Xo\`Dga[8\KVE>Um9Wl@I
Qd0Nh6?6gV>E7WMR9]jikUnBLIC>lZ]O59?oJ7bRZ`GiKOaLf7hPE\0K_jWqkL3R
W>gA^JWPIW=djTe;42@1B3?eo5KE8O4;dg18JYS>bC\DBo5IFF@A2;A4kWc=G?K6
OYD8SoAdJiN6iSKhB@KZ>KAie:G4kSaF3g`l=7NZe=ILAAF5RenLSmqmN2Td1AX@
7h0h\DgBmS0:@FKod^fn[J`al6E@FY?9lo0cnU6O@1?X9:`L7YUjK=Y?14K@i8d2
NXGTCUj_61=`=amglp49E@E6qcPXhKfo$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MAOI1(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
DT;\mSQH5DT^<@SDDjU_=LMQP5=IQ:ePO3R2`0?D;j[akiW6SmfaCZJ9>o9p?0m:
3809JQ[Z`Ml2HLBXeUHTiSo2B5mF]fke>cH1Hi3PgJeXiYpV;1KoT9mEL66QUCA`
K<KS_4QHA30Y>qR?M\4OqMdkj2;a;LbY?inV[h7]ZI;U\H<fUR\dnTlqQ0P>JLnE
5WIAWn1]8`bo[_o]DgKOZ9E<P=qQh?<oD7>24ZF^I@NhoaR2;I^e:`5N1PSq]RVB
hAO<Z>VlA9YZp[>GaRm=pQlH^[=qE9QSgO@BP3[1GQeXjkXkJ>R5L<;>aSYFR1Xc
XPLeDTYA\ZEbZBLK6ZFcMMk1K7a;EN<<KYaaNSLc0dW9kfHT=6iF1M_f8lTL^1WW
3K5NUaW]EkC=F[X`i9qWgG^c1obI\<Eg0Q=Rb^\@iU]@AVgQ:_4;Kk6Pf8cb;:na
hicS1QqN2<9I1Nj>jWE:io>@V5o5_Toaf?[EVk:<[C4`0N5^F6>o=8h>5dLZWQ3A
=0Z;6b[N43Sk`5k:52WIagS5@_RbS8>CGId7?77O[GIe\d_\7;S>X<D5HAn;>p^9
ofBOcD:Fj]Q_98_7eC5oIK5N`Ka@k5\ASljL\V_5Z1<N8hD9S;F:4O:LWbeC>m^[
Hl8Cli\V]3IE;PnBQ@0Zf112BR]j]VnA]:=joN3U<PbU4?gBe3]BpCj:?oYdglHE
H0oLLgeMG:k>CbaJ6UoFBFThR2We<Km`@]10T]8\fP2a1T=6:Og9gCe9@A5]WkDQ
MYSHSD8Ce@5p<IHdC?Yb:@798]`bVIUnbgU?aBm6kON^AF:J_iY=gQhPAJ^<09P8
ACUen`^fRM[5<;I@?97QB2U6nJkhN1n9akSTZ]9e>P<[_F7[]W68G;Nn=cl^?[kY
M7qZkDZnD9o@hJjd;L?00_nBHMe?3^I4TLH_i6A06ljIo4IX3K^Ra^Il@^5mYkFm
B@PZB`3E`l7nBiiLQ`\I?C4V`BQF8e^jMTiOiXAVA0CbgA\YXMZgMaKi?p]G?[<h
2<k;=5I>^ZkXJ10iS<lQPSJL>p?T1TETaN:@oQM6RdDT@5aY_BjM?LRCZ8E`9da^
Cig5FSW;9CY5jHeZ`gQ5MYS?;]?;3BF[LHSUX2;emP3=ChYkWPmMRa91IRn`K?T_
;iUUi5T6fAhnh1D2pBWQ=G\K80K@E4>6V6oF5`X`C5J<1LV6IYZ2AH]kib=FFJdU
bB;WjH;BR:>5`M^7BBbMenH[A7aP0jY^[gNbh<ip<Z\ocn7m06:?fBd[\V8@:gKL
UK[D0V5F5N8J92jc7fKU85?C@oenR[BU3nd68SHd<NH4a\jS:;DgLMnCiQIY>QIE
4KfW__GblN9eTUM>Td0C03_QY6XM2Wq92?``53[E1DlcZDTUF`?48C;L3;JEb8XV
oh_<6Y8JXITA>_JXYcJagk>Al8KN2289I95A6<9Z09Tb9E;?AH^1nkSNm?TS\]F1
oY_Y=Co8M7iB4?;i?_^aWq_=QoM\YB`H5JPegRO\7[a;[=__d9_P6P`NkWE=DK<e
F5LDa=RC;5j@ieSd?GmiE4_P[1W3`DdIS7kXJa9RS2_TEY>BiS46I8fNf9A_4GGV
caFXHMAlhM91qU4`e6bI>[8;@E9J9ILkKdiB@21CPMo=8^M::j<Z^aWHmQZ1lKI\
KRLDkB1MfIZW3Ug>R1Bfa9RjUROb:R6F;0QqBZVikIbH<F;MI:MKEIOo0k4JP729
dhfo_WCkqVUSEkjc>^F172]U0oEKd`IHFJ\B>T1amQ3`ohoajdT?6LjcdK_8j?0E
V\3OV2;AFVfj?fgVKgFXNR@IP`7DSefGl=200o@^K934l=Mn?eM_mWbZR4WcBGBp
S2B@Il9M:he@OfL;ZnS3RfgRUM4AAUjn:h0Paak43O3BJP:XbE<>4^UdKV1R9KNe
SQUjPU`W8hUE_RQ1diR7SO6?\ZmdK<17Lh0K25Q5Gg<oQ4Wcl@00b<p7`_kVN1F2
CQ?iTM?5h[Yn711eAO^?k0L:Oe]M9faYbFjaYDR7`g595?b?chHF`]I7m];mG71d
Cm8KJc:I4me;hOBbTQZ>8?QoOfOOTn]_^j^X<d>]bjagSpl80lWi24[74ddZ9gSe
oJ1?kPmOm`5OX\E0T;?^8<GOE_gC?lc`LaN80IebH7W_cjlXCSm]FF?7f5P<KJgX
b?LPpZEBSnH=Do2IHFQ1]mdfSO[>nQ7Y5L7WKJcmEMK:b<Ohlnaj9n=IaEU9gS<T
8;VP[8@mnMRqObmFL8qLYGQDL3$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MAOI1H(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
5nWBhSQH5DT^<=chcUb[lSWXcho_0eJHmhNo@T7iLFT5KUO7G4_nN<9P1<Dad<ad
LJhAJegnBgpTNSf:1\[A836Omj8B0d49U1^6GlA?n_N2j<VdFn_`QG_]Xp^]3Ukg
YjakYbYIXXWX>U9XmDWZMbe1d^N5jRq5;P_8LpjAjd9Z17oOn2<Qb<iQPi1?:LeP
?O\E_2A8qZT`7h5ZIKJ:YGl<=YY46YGA4Y^NQUL3ERZpWWE<VeC4cAEhlV63;biL
O=JJ4\GniS[mpg5O`^^Tq62fN^dp_<o14SBJGjjc2m7cW[gZ7X=iTWZ]U7Zn3ZL`
TO^HR`UG[LSC=Yofll89d?Wl`dNX_LZS;4[abTN7aJIP?D27?TjX5KoY>[4mKZ6K
XkdagY`=2T^:QFL1:DqDFGECo2U_ljE<:JV0ZWT?cXcC2]PnQ>p^A=BV:N>\TQAS
?\QZ=jj63AL7;RolFM?QRj@VY4F7=ZX8jEj?2n3N7hO0K;nRS6Y^=]mMhjX[SDh8
]YV@NCmD8]45W5lBoFH;RPo>FX]M:AO3RDeAln<bbpUGK`K5K\KkF<ZRk@1T5Z@D
Ig^Im0>\R`jT:P2l]UNIUiMMaSW9Non@H\k\ROAnd>UO;fA\3Ln8l<3OBB3DTdRk
H57CB`kScf:TmnnPe`1]HL3:CoE4G;IGqBAU0=em_VJT8GBB^1CG]Q\^8jMQH;S2
505:]Db?WaN:obg<@4=D^Ec1<InJBS:FjB0R0i<P>MKCnZOO11:BLnTp;<[m=><f
OY=VGfDXWfmNF2U=>Q<1=6@@dnMN6;]U0SWGj?RW0Hb_=4E0VQ5O:O9h;8[YKfGB
Y0O=k^\aJ5_8R\@_LGg?QYWCZn[VUB2N]QM\B:PnBjiC86qVB4DeO1Xk1>`g3mG<
WYM\F<I:=aP5[`@BETN]Abe>49P=[I1NFcG3XoW7J<_DaMgV:A=9MfAOYM0Uajnb
kZ1TfgK8J@13E6ERETh[Ko:@L<X1[D<_A43`?qXQbN2;ej^dKfLgX;G9nHciC^M0
G^[c7LVoL]ZF@KThD9SHjakf`\U^j1FLfTMjCBXB6iBo]AH]?gfb:5JDTgGYV_Bc
_W545j_oW]A>D\Hf9ejo_kQ2gO:np=^l1Z[WFVX=i<]Tb9Ua:ho:[^E=BY4U<b3O
2Vc;mnh[R80MO_HiH]Um6O=3>75\1SAb9m1]qM_55oR]eiRobgEN^HfW2GK8KQQn
S]LA_OBbWENm`jk>XaI;_6W8<BN2>8QOEd:AfMLe2KM\4g5Z=GRZdf2c`bDpFcNL
nM\o@jcb8J9bW;4e\c4==03=:km9fU_6B\3\jIG@M`\?\7fH@5=`]6C0kCinF\7L
h0ojcj_l6H[<lE4`h4d59\hGn`aoKU_bR2LDS2b6NDe9k=JeNBpLeEQXOVAF_nQ1
D2`AIWcNmZEIDl9D@?4[oYXjiR<O?niBXZEIjRTM@]B1^X]\bcaLh0:9]21R_HGI
G@JK[WYj^edmSF3:?YR:oSfIeWSb6CWiE1b;F86ZopZA2Zje[T]<`94SoDLE[FBO
aS]dDFFnnA3@8BEKJI@TiEL;jRBDD?J]\GcZ8KS`eNZ]RTUId<o<o3@HH>h;^9B8
C3dIQFok4ec@M1jjhXnkhnm7E6\8RL^?pnjX]YhTV`6XfFWaKHnB^e2KCJ@DanO<
YOCERhe8nW2E3W^c6W3\;0ZP?@3AB992knm<ZlmIfA6UIdP;D0LaDW`pG5=A?_J[
0@fV]6kYJ61510RYYUCA60PLY8N343bC8>FBZVPEInC^F;hkqG2bh?4n;NeZUkN@
8:EM\ZT0hniWHQ1SNfVUhM1J[CGH3=BgUc7g4Km2d<_1bZKK=G1P4o?YGge7Xg?f
m`=P]5?N<Zi=\kXY0\VUlcWnJ4U3572IF3m0gX9qnnVG3;GD=QjFm?gKS`fIU<R2
V9A4\012Q94cl<PFl:F699^WBTPe;7E;SnmlKCG3nHTMNK98IQMAC:gO^i;RR>C`
39?e9SC9f9[mngM^?5D9ZD:iJII2m6qCXL0IfE;JX20E_SmW[oHRCOXgF6T5Fi[9
IDEMjOocl4lEg=9I:0beBMKD_PiibHdCCGO=CE:^XMF;NLBfIJV7M5CCF8UkHVIa
IKIKSLE=ELGT9h_JkY9gjqH^e5`99Wia[UNWf]nmJMU>JNWBH7?cn2G:hCGEWQWJ
27PL<ieW\O<`BV:bN_VniaHZPX0B0X^aA_c4KFF`0]CYqdCKmc2qBLHekO[$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MAOI1HP(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
F8V3PSQV5DT^<19KG93?glT:C4Np[5ofOYMSH]4A;IoOTXA3cKqgWMES8:H>VR[]
XDdYc[pR2cYYnpF46[;a^hbXBaD=jN]>SH8[f9;UgOG4j3b0qjK0QF5LXol]a3c8
H]\XELQ5=SFal^>3PHGpS3SZV]m1eAijBV7:^WQgdT06oYaiR]1PpH9<TF\Zpc:0
=fGpm5J^OJCOi`7MLc5`bO:]nb2gMbDcQ8hCKKDZS@Yb[@X=`3f`DI<GaY99U7i2
lNoNmfkL@;2OU@ofcAUAiW^>OS5bm\5U8^mTjKPhX6`[NQ86P<U@ST`GX1pQJ>PY
cDIdESc`Z:MZ:RI3@E?i@fSTAWVZUATZiPYQnSgaCBagRook^ZjKUJil`CaQ8GlK
Ub8AlXEJQXjh9HD^WdAS[70Eb8C7UBHcVVYXmA=\IKOH>T^F4qCkiEgmOb>SWg^1
0gg_2f5j1KSo=2>VigZ^UIWgK6ORK66DTjUI=?OKTp1ZZdG^XRShiaAO>YddHLc[
9@8oOST:5<=3FTl@dB5jfI4bc\VSKnlieE;hhFAEbB1=>4bNQO@EgUQ>m85f8hZN
:TLhoL:3o2J3M5A`H3F9`bA[gVj21RRhpJ;WjiDLC4A]@EOK<9oWY>;KX284UXiN
>5C`WX6iC>3@FJl^EFVgIZ\O>Gd52QZ7<J<1E9QaHCD6Vhk?T5R5dMJqTRVSBhmD
[X?BL7F2^jC:9>D=dL1QJ_SKUb\fY^;=Pj2g?]`S3LJBXBKkFIn8UdYST<EDmied
VifUL\e\E8alG9nbCS8c_3UR>b=M2BeRl]emh2UikE1aWDqgMeX`E=FTiMIU3?_F
OL];?WXQcgP^`egm97iijT9F63774YdRl=BLUljT]=X3l:BgTETDFI4D0@W@:Cm<
kC3FRL7:@d4WeSLI9_WREoA?Y9CYK50L`RMFOq]m2B?QNPC>\gR:Oo>>FHVm6^g>
gnOF\@Sg^o;_17C<8;=2h?1nhkK6A0:N[l\7af]dFjF[?ab9Q2Y4??o_;YBJ7[Sa
Mo[`n=mgBo7c>PmNagjj@PaI3F6lpG]Z_fBK39``MQUDKJWEA_9nZBZ;JG0<KQ1?
kR?PVF9VJ;T7kJ;eW=AVM?7bo6YjfG;B3aHZP\L5Zf=4=o4cm>Qpil`_OJ3FjBbi
]ND?J`5Ij5IY^F_L;RO1RCOaFL[1R5Ba`fK8`1?iY9^DVh9eF=c[iknj6US1PBQV
LJYdA[5@:oe1IM]=_>F[<C32Fi_In473T>B1U<2=AYqJjoU:cJ;;d]STHKH1T45L
?kNX:c^X>[6[F`qoLiB_dZA_2d<<kk>o`_d1XW6H4c5ECo9N6QYe^diKfEAeXV68
496U_AbN4WS=eD_oZ:oKGeJ]2;VFU5cIl_h7c_AKSngNJ4RZ6aFm39W<KCYo;HMX
39j<Vp:j=ONH\ZS?BV:<l0eWNG;<f6TV0FacO`W6EQP@Cl9=<jN>5<ET7^fMHb`o
D]Se[c:O?d?dbS_?^ni]6:Y:Xk^KZI4_7X:g]LB6UOLU:Bg0lbbM_e1M7lPMp8^N
=QN37Q8HF_3EGkKYLlJ:TI\T?Dm6d1kg3EJAG`;BiLDhARGJhaMOI:5:>e_ik8I\
<lC;E]8B2^WJKZZSQ=6pE;ij@>LJ<SPSUd58mW5bCh4Engd]LXZJOiiDoK1KF1aN
Y17e:S84oj`DlR7oCZm6ES4kjYMNTSf6``ngg2<nm4E:S^]Db]>\kiU5VU]J6ao7
V7e8m^9P5mqYRTG1=>c1Fc:6kl50LbnWg4Z4Xg0GmmFeChKKWA4L;fAH=R_NDLRc
<jU2K0ZVUAZYLP3ZlGjhF9?jFP`^h=W9dP>SI[GUi?VWCgUJSBFZ5YaRdYWM1Z6T
6q1m`RVB`Xl89>BI`JIB:hkXbUXgja0MCQ:9]mZfj0`SVSVR2jNT]Fjj;YEiY@Uj
[Z1ZZ;ml=R88UdXdjiNBdYK9EiJV?8RL7UK9k[H4_Jf9TXfeCfBWNC09pk3j]S?o
j@H2iC1H=QfaO_JFZ]2<1\o^3FCic26^[\`3@:4=3Tj;<UATXcD\^iR5dkbkOI>d
0kHijY?62n2XE8oqmDjd2>q\Ni1<TW[UkobBgFF=U4LPYPopMcFYn;>$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MAOI1HT(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
\:UANSQV5DT^<N7X8S>9:>YgRJiWFT0=mOHnfkQOpd;SV\748DZoFmLoDM69Skh]
Q>iYh_]kcp7\oW5`7k99::4bL_YVFaIJ<3g\i2VHCmWo]oICQ9hQ:36Icblk^Xj3
Vj4fFje:a6X[MpWFR\Lmp:Zdf[B\UhCghA2HfUe9BcB8Ch65_Lg[n1@p7IJ\5Fll
OD[dh8P;AciMGm9_NgJ?_03^@dqeoaog]MecV<No]PW;1][;[JNYDiTWX:GcnU13
fZLMT=bo@oNN]`5IBJNCK[gEWMELDa=nD:LpK5eUA7fXiQN8Aag``h\i>T<@OkFb
ffU?p?4X_JE;pm1eihnq9QbYg`gM?4im>aN?W5ZF>]a46n2G2[;\5;=jRiKW_DUH
95GiL<>MKBDDc]c_C4fn9V7]5on@F;<R=bL@cEHLWYcWhRG<JU0jf;jCCDMg4;:U
T\\OQ7WlOkp6=eWU\IAkfXHdig`]EHAoh:1HifL=H1<T2gj<kEE_di336FPBV1ES
1BRQM>8h07]6;=J_RHm5QP7?hn6]7LUjO8E@3N=<IT_;2hE@Tl4\1;>g<CJLWV^h
iq68n43QW0_N5J\P59HUM]Ql\2;[REID5DfQ[fLN2eBNOHTD>QI2dGAj;gJ46YF`
VA\6q4G?^dAkd]82XA^;@gO1]mo?1VcPLa6Y_:__T6GNe3RJ5R;[bbl@k4eXEKUD
7;KTJ4;1<;bi`Zl2Sh:D9Y>\mFB>Eo`Vb;I5eW_c=iK`^4]Aa=7kTk`;Qc0qOU0`
WadiL^7WNXJPiFWM71DkgAIWTN^=CYD\^f_Cf2oF]Qi[hO?GFSU:@NjnemLaO`3I
<mSTb`>D;a]_0RdN:nqaCk7S\hPmoHNk7>kcRHM3=[ihfDYM4gmkdD@cl?[HRa[d
g?<SJUa6^5oF\13KFK@adH5=Gh_dj1An09Q18]h25o5W5U:O2O5CdiR@j[PW9@EB
aJ[IHdDU0pj?PK@k\lV]DKJNA8a69`9O4q:[[_18Y0O^c9cK?8T=gX8cjge0ZWDY
=C=0K;108cNJF61P;@jHiO<Tca6<4XVTcI:1mSQX:[]`V=CdELJ=Wo;D`am72Rl_
ib206@@WGoPCnPo`i:Ne][C9qES85PJBZ<:K7mKEjoWT]@cGV\GenY:W\9bhKf@i
UQ3EDmo[gl>_A`d=bcJdk;]EeEZ?NIM\:8N]XR?MFe6fi:0L\Y?8O@Lnf4b5nj5>
oEeRV6X=6MFbB?8pLee48]SRTg20XjEQVl=R2Hd;mNH:e3O9[ER18KJ60DQ18l@n
BiSV?\9ORA0^AO=lLX6O?_7mAOBP_IFa;ogCU9q71^2R004^k;W`N`c0a6]FA4ND
_^QnSGFIobck<\AQD23[j`S?n@K1n6lckUeg`iG7gaWbONm1kQW7]3;Cg6MeG8lA
7i:GoZKioIMWZe^^n79XS7Nk4eD=lq]mk1^_IMQT4_UAaJTXKeDDEHh5W;93bS3=
VFL8MGL5kMIM^9]W3MnYo\\8SZBCJL];kH^:Y9DT^l[53ieCKeO8l<GdfQW12Z9=
Q`iI0CIGIEFmGlX]TcM^p7oG761[APb0mb@S6Zg3=lZ6kKhLjfQY8oN9g40kjF^O
SmX^i692Xad5a6Q;8aHQU7fZQ]A7_9b`V9Q[JLf`himgR[Bno?IlNgN84TmR;X^G
FfJ3RBF0H<6q:1HdPSL]f3de^cn8AEaTbUGdSo8B0P\5odV;F;C5of^OPWf^<9NO
UX;E3YHRTT6R:VU73?kSl38DD\k1YSa;>Oqcik9o1QXHT0?K;[@^E6L[I9<nBS0]
[el]lWfi`BQL_8JMP?>6AU@C=8?BnWe6De`c`O9AY^DKTSAlGNU4Ca6IB]m]E526
F3K_lHX3ZgW?WFee2SH\Kg3h<pZF>LHPgW=YmloH1SMFinVTE@5C@aSn>Fkl[Xo3
d0]@9GAG6jI0XOLgeP7j<3`mH5Zk?SG@FWmY5FCPoTSa8]?SAUH8][m_YX0lOf@n
NE62:hX6HFD`0_5PpkR?FXIY85^TEYXblXCJO_X7;aGNZnbONB4iMW`qhicon5Bg
UT4E3PDk:74:6FSHX>kn=_HbRX<RgD^i3Am`Qo;bLKo?mhY4M?5QL<mah05o2DUO
[TUUbPQHXeF>Jl36WnB=V6K@YXJ>A6\2dC`JdC>?V6U6]GpHOYV8<EQJ>9E6h>fC
`66kA<6=PVRNVd9WZYI;=IRlXn[\[<d7GYeg>`7iOCbVOWFHP=LBcJZP>=470aBj
@Af4Qp[4T<C2p>0SU5LT$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MAOI1S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
]GFMoSQ:5DT^<n]R5SU:<T_d2Qdh?VZmE:LiM6[@m:J08K8`o;XBM6qZBShSBI:=
Pmf9`W73l6i1DHYeQc:lZce<;S]50`q<C@Z_;Y1cdLDigRi_CS>BFDoJKUGdCTY@
WX9mmLFl9gEHNZM>FEN97;K]AZMcIB6OdqWNMOFbqMm?88Qcnahj?@Q977QS=m74
ATNCQeT@WX0pGYZZ^0\cGXg_mYXd:cW[b@HTfcZjLW:65Bqjmg4@:^96aDU3<1iY
<D\7e`f^]5UWEcBq@h7bkhPqOVhbZBqR4ANO^d4KI?`_LGIg@YXgI_6AR7Sm^n_H
LDZZ]S5O4cgmV0oK:6J[;nQY7>;;F[XRMj;\n_LbgjneCd`<k56VX[khg_UVc96A
Lm8l0o9COHQl>PHgEPeU9pWXf=jL:Vn?OfnaV9_c5HDh1kGPoC^mA]B^HJ3_X71a
RD9RXJDnFiWE5`mHmZIXC7W_Yo4mI_OFNKjeS;DXnViLgDejDJJG=]h^g[]G0HR`
@`VliTGCm5^]qGCU?HnfMSCm^XMo\ae0;nHGY4dO<783]^@\SF>;0ed_bFB7^5TH
1gn2SHlUITbb2Gf^Uf^\5n;JcaPYRAaZ>D8G;F;C\4KOOl@[e1mZQW7EjffnRg6Z
H:<qanH2c3RnZ^Q@JUV4a3PW>09Vq?5P>em@[0Xn112Cc9SL<[LL;of5CJTibHK]
nVH<PPJBW@j8VI^9U7`o\Ijh>mQJn?@gmX]TBWRPWfHUfj8L=DEq=SW:n17\9<=C
RjD@J>@I7dJ6HUgGak:`Y=dG==6dBQ\O<ZL8IdiY`:mJgV4=GRBE=Om67AM;76PA
m2OFkae^Yk;]2<jYHoEE6=dEOUIl]l0Kkl>AhBI2YmqOca1\Jd6>C=2lTRDl=1jM
Oea;V;VhU?8X=ag8cVVLBMn3G:R;l:OM6J]SGoN>8^iOQ;f]A0RLVXL=e<@N5AjI
kC?]9Qfc>0iD=3PeJK@ihdd>]kL1GQk_mp2SZ<5nX9bj=7N:\3`<>5=DjKKCkACJ
j^[3okONW7a5XgJTZV3cg`>Gl@mf1;0aX`2\6=>S??QUiOSQ5mNOWlFMV>fLR`\0
1G:3HnaE>k<Am[4H>b>OK=ETp^m4M7ZSHFVbd`^ZhQLM01@i]@N4Y=X_7B?mUWnf
Z`9^c>k_Fj2f>X:ZAS2d:nhOF^7:]d\=kLE9R7_9gkR:7Oeq0j8k]>I[X[\mDTO@
7Q?EKejCU3DhjQdDe>A:10<[>jm4WlN`gPaR?39WI=NNa_I`0bam?h3kc=:G60LB
ZNS=>Lb^=M2Jdgb@_>nM4@25LcaAYRj_k3eEVApOocjkPolj_:\oHNmNKgX1T_j4
YT5ET7i0ZnS^P?]bdQFNX0Oe29Rc\?<Y9QY?FVOOPYl]ZcO?<_E5]HMPLCGbHjHk
LaTKk6@FZ4R7X1hc6c1T_L=jFc\O2ph4=1fMLOXhjL=4Vm4:DaL=6Sfg@]5b^IIY
;2UhRKR7gOm9G@jEZQ6<DY7Tb96c<RhG8Q<DA^7lcee:\gO;=[:h9FX:VHDc;WJY
N]:[C_JlLhNk1KZ[QmG`pHoOCZe]C2i_k9:M77@nd\OBKJY08c4f7VU=fY4TePoo
G_9?@5Y=p1\Gl9Goa9S=Z\i2@SU]][nHCfT@k>\oYmLe_51GhLcab@KLEU@fXDLl
UN\BEe]m=1AkfaVDdL]_2HLePdD\UYmp8eaCdaO3WNFoOHUIl:_bBXiH9Dhe3T?^
knJRN6Z^in`3A06Jkbd;f6jZ8iWQRW`H88\LQOSYN:j:A\XMd_N;@?U_7DgCIhNB
jnfVH`[oBM];RYWN^NJ8oWqcCa:Z];J5R5TP<I0LTf[\=[Q8[Mo344oogF<H?Emg
NKKl6VQRdX;nTBmnK5X5iWTcWfJGKODUC5bm\L5HU7E`;@Xm[BTUi^igg@:l4aTW
D;R<Y?RNnkm<>qBVDhCG;5cZ18OC1>gh\elM?ldJ_PJjcQb4nO?PZfZN`<CAd0`<
n>E13Fa5k\?INlB3al8EY00B>HaKb0N6HPEbKV`JeEHI0W>4b_e:FK;J1Pc\TUTj
>?bnqcPKl5bMJXFAAF9UE1hjZfgQ1;05kFR=hX[?m]>Mg<gB^4[cP5W5O3VZlB@q
34]JQ2^^[SlPjh_f0:EVOmeM[S;[mN0JmHYPIQfZ:D4<P3RW]\AU7X1hCEf4l:ie
3i@5EE5\SAUSVV_QRNNDGHq@\n5cGp[T5?gVf$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MOAI1(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
`UYkCSQH5DT^<Q7XhYJ1^0oD><<@mQnHZ_<m3nYQY9@_JK7ej;:bGi=60lO\JKWG
WGGp:ZRoJ3]c9LNXg\Nb`fOO<cpnJFZ<FglXDOXQMoFCKAF1lYR4T0:23aoDfF@K
iGn?_4p^^DVB1qNRd5QU@15\2d>;\FoAQSn3A[IVfdj;De:QqZEcP9@@VA3?_JH3
YB]gI6Bl`_j49?]K4T<poM5MRHoL8Wf]Z4cnbJ=I]aV?iPh653a^qH2O5Fmjl?[l
lhl5[6efhQX6JQkGiY3ARL\4::PofB^9^Bc4YLb0_C8Tq6=YA]7Yq;506o1pCYh[
FM<idU6kHgS1HAW@Me2KhC=C9emYm8o50^iG9E`9NaR@P?JHm9=nH;7PhgEDCB1^
BSORQUD6N0U5;b]P^?[J_[IR12>Fd8P5`jONgJ3X9\WoI>1oUUqCmV?]?b`^7`XB
M2V\D65DR<`56nm:3]`2BCBl_FMJ<omT`;M@Q4`M56;^bje=]:7C<6;692IO7ZY2
1?lfDhPJ5@aeam[koG4^B2Ifl7R>g]b>@6Q;nMmU_q2B5I[SCSc\i3WGAf<<19SB
JhGEMkDdjCIn_HlUiY<3PYif7Qo6FN]ci@jZ_W<Yfe2jeT1d^;:\;:LF6ddm:37]
4i=K[Ifh4c4n`Qd[Ed4JX5gJLbM;=2DBqMD`\JVRPgNd5UL7GD6fT3jV>5laIIb`
QhaG_MMUTaP8@Rk[5=lRDj7D3AQ@5_a`lM=AT4>9ZXNEDfA0UmV6_d0qJPO>>c9d
bg<N]>niLY7dgkFU7G[3m3LeGSfTGo29kFPN8Fi]L\OLqi3H0NVZGabc?Jf`lTbI
h<e7k4XSmBTl5W[;Da8W31hBNmlBW>LCGCSk4?R[Mlc[OiCkcHh:;ObIW4eD0j7I
3i767KagLKcE19[\EUg=4_^dIJJ6?SHPO6SqeWLDb8YD;BU]TIjPoi4<7:M80E;>
\ggc?GDSii;NiAjDgOXOJJeI;mHH8`XQ4bDMeoo\jbKUNBdBm<3JFT6UPg^I94Aj
IU0l7GLVWQ<><RBJbIQQ=:bU>hp<I?a4ZMl8@c?PKi]WEJOAHVS9L]K[aP7[c<S8
0m\Ve=1L=D@8]R>AjL1Y>LSSQTA<B7^b2@HW@ZnY67aJGSbZb3KelnEjbn3Nci4E
UMl?mj1C^0na=d9Qmq0MJ2IJ2jSWAh0]``2K0l=]2`iV0@C<mSn`T?f0;WMfe2]C
\^N@H`=2@>]7kaMD2b0ZJ\ABGCLW8OcMjl>3`J;aqk54<E6Ji?>OeUCffcB<PQ9l
6Y8lIK`<o41_l\5n9o;1>Mo`]SNUO\9j9>knEB5MokFm^iVaWScFb:k8mVX65e>4
kWXo]P4iC`1e9W[M^nn8DkUKLS:9=<Bq11i97ec`hlJm2gC1gY:TLdH452lioKBM
>PHZFYYGZg7UXY0MWE1>SWPhXHeDL0:h1l5GaDGlKh[2S2M9JUWO909lm8ILJ2F2
DPAid6\kORm2b\9]H\6ZY6p><gSFG@Q7168BU40lL^QC83225;@=IKoh22Woa]IR
Ijc>WHc;KT=;f6m03ebk6=O>5kXM:PM^4=U7iKlU3o82RFXa<L;_=nio22BXXQ=j
nI]>D`235?NB1qn^L7f0N1jaI:naUJhbI4f_>a:12CI^U46U;;1@dZP5i=oP^i6]
<eWgFOdg`@ee]nnfM:V9`ZkP@LcM0hVBmD3mqC=86@hhQAc16F:a16j__5KJph:o
kMf?h24]:i>gc[cdA88XfBU1IFd:JeYOl:[7::3ZT?^M13dn:[7n668nXgZ`;hgh
glNU97S<LeJL7kXl9L7h^;LBmI`SnRY:JNLeBG1[N0`lb_S=<\>q^a02T2n;VIX8
7n`8?;oUU:l]Z]TBJL<Q8R2P`RGG0Hg05M[@@4UI^AN>4>E@6Ra_^YkG3mikBhba
U9^@NNc=YUkCa1i]EAJ1mRW@_[o\=C>Z]fX^8MiQQ[qoS13`4921V[8[l=C1hGlg
C@5jVFPY[1f4FRD6QA`MU?mB?]36AfD@NgY?f^2<<3Aof1;`l21;9=1oGlUNNeHG
c8WkBbIoO8[TFZD;dB<4fT5GJGHcC7JDBplSN3@C2SDkIZ9;:>cbLZZ>0PK`8@Oh
;ifBQ6631>n4D1M_jQ9Mf3KoRYiBM6FOTolEbCk9Zi7DkZ6CWhIgiDG_p[_2i6Ik
_=?j5kE8o01fXBl<hc=:JF^;C0TWP6]_a2FWDPPHP\@7pgmlXQCqi92U??C$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MOAI1H(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
S8W[USQH5DT^<h=`7m>\Tnp?4[Mho9iE4KZaC10>fKjDQ=;SQiPL]Li5KPAJ34VP
71j_jA^Z[b[n\H5c=JCEed7JC<iqhaC9ALZf5^`>KiTE^NE2Q]6hG]ZH0lR6g[e9
hhVb;T1abgO0L@pH@^CZmqmO?;n5j5EH?cbR;>l\nHWB6C[CiQjJJOV?p6\mWT6[
JkT1U`:`D21HUcSE<05n@;>bTXmqo213iBN]9E_V8b^c`UWdS04NFW9KlO\Cq;ZS
k`Dkp^mF3U:[H8P5o9fgHP:30oajW5_HZQ5:LC4c6C\]QUPbUFHQE8A9__1<9Ih>
B12nfq1Wh8hnq9]PJ^[JKH<lfA^]kPR>3i;^Sd5SN<JcHb5Y48dMGl`4fl=DdXSL
1V6]BPl?aCWJ09dV?T_=_d<f]`O8e3T@`KY8=A0QTUBi3l5>T5CJ_Qa?aJe6R]<H
Ogkp3mOU??`UU\oMma@PUHF?A95h59RAFCc@DkR8]Za8]h:R?^n;[;cQ\X:kS^[j
LP3h3bClef7X>\U>SELJ0kZV8a;C1H2XU^;g^kd122fFCP\Z_nacXVUXb2qF3UUd
`B[:aXHCamn[E5Goo:k5D442J3F54XV=kQC:OkDOZfkHLZ51YTXcFoCagG3F[\]o
Vg5=a6JSS7P?S:C7NJ=6NQmR7SMR4i<gDFhJP9`5m5EJ@bFklqCc[32W_;KnDVFb
W3<VGcL^\<FYH52fbVaHl=I\P_mE=79fNE`LL8DERiBboRe[_NCFN9K_`c_nO2J`
:A36NN1YqfcnV0e=`MU`WW0o[:;LKo;a=7>f;9d@^;aH9Ice9\;NlEcA=hBOV<NM
WW=a27A;Hf;dV1O>oFU\fX]XP3<LI;_dkM\>;SnUAQa\jj>0Qcfl:m4a^?;jkDbp
Ua4KJCAK9^EaAg>F4nRBkD8iDmCObRl00nOQJo]_VN\=8IeXI4EO5Q\Dem;4naSe
Uk5n>5<9L^i8MfL?G4gcALQL<=J`5\gD3nf:GWNN>DiPVkX8D3i\nBpHmB[nB?D7
]=\=Hn[hbQNOg[2Db`11`h4]Ud8Q<M^]P_1HFS65ESCP0C2F83kJ6^DH98OnkUl[
]`bK<BLC83Y@>\5G[6h@DH^GUO6A\Y;;UaKPokBQWCP5aqF_=K=hW\LEGkoKaJb;
<aQFmDCcV9EnfO6aaSCNJ^QP]Wa`;egg4OWKE[5:ad<6T1FXml_2c[ZEiEA1WiWj
h1HUq7ciRX9PD4MPcWjS`anmVGScYF2Be\4<1;O4]X^V\8E77q:9:5e3]8K>kJ[7
1k:PNnTL2>H6TMEehFcQeKeg:D^^B[cCAb`W5G@[;<mfA4XRbG:6C5WeLGI2g1@]
aPJ2iNR?dPZn0Z^4Hf0QC?Hl@BgdM:DZh\[dSk<>qZTi3R7]d<3B;AJ08JCd;5?n
Vk;D0hlie@8DegVUmaHQEJU5l0?2RkU>aMgFnHX?KZmlDA`EUTVMLi?WXIHAMNeE
X_a>OdK@6\8FE1DLQmEafE>lR354jinpBe>[\OJBODFd_=2@d0:VW>G2TU>fUK2`
@ldC60?669YiN^CS6fgLRdK_gVSR:o=YBJJ13D5od_]2L\@4^la1=JHebgab\6l=
ClB@oXP[N3bNM:Lk>Ca8JTpmMU;95kM;Ikn`1fg>OIeJGD49=T;8K2kK]=QHbZWj
__fC7dME_M[OnH_0WZ?MXURm^@5c_^lOJ6dcIaW8j\fA1qf;S:ePUEgT=^JcI1m\
HfDnJJ1]I73eGY3==2`R3>m]eWje[DBmIVTj`JFZOe6l0LfYcHDX]_?_fga\bfQT
l5G6KA>]fjSR;2f=^1IK>mIcg]jP66JM:KeKqOB8b>okXTIWPnaG4d@BnI:0NP=h
9^`m=1ZXoUS=pF@Y]RLohlS:]SXhbAj=2haBDWd03;@a^C1DMZ:NU\h:HcWLA8fR
J0_NfMl`<=B_YF<2ca_0FM\>;SI@_7aT8j>0QcdG<mEB`51BXH6@ZaNAlge_TH?5
fC1pN`7bnaeVUbmNFm?E1?P`Qg1ObC6TgD8]8@<QXh\:0Ya\KjNM]NoGMNdj_^AO
kIZZNcVY7^AJSUc@Zaf\NS;=HGNO5[?KUiX]e@jDbHOK:IX^4Q69<=\V2hpgeO4V
fn=>e9QnH_4_d>mAhW8Ca1eY2:=;HR59MoNoeDk7[7RMAC6cDAn>VUM\NWWg5O`U
]?NQHNo>N46>Bkod0p[\hFfoq1Fd_TGb$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MOAI1HP(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
3GIV^SQd5DT^<N6H:BgV`RJnAHgXAh0^o>4pgdcL;64>kb;SeN0MEBGggU6Fm5_]
`=Odh5H?9LlafPMNq6e0eTRS<K4B4a=almaV0^EVTqX;XSg2paBVW:4`jS2h;=>D
EI8J`@RaOR<b7AA=A8OqJ\VQ=K`7]O0d;gVDElNaeY`FHAGib9^XD0p@Mm<[`V6A
O^dE9aCWa[e9a1POFSF[K@8q6jHbdn:q;eRYRlpaGEfOfM@`86M0f>f=MFB3`g94
l34RXoGA:MCQnE9?jqNS=RU5D\XjPK6R9b3bF9_hCm24XVmOhN7]TF43UHdXD;Wc
`jjOlRhLT:Ph2iUY[FN86C0A3CVjdQPO:1:^R`XlQK^Qkm=KJ5U]78[M5^II^maC
Tm_J9e=Wq0@Sgi;WjnAX@C8O_5kUm_7XP@2?5F>hVG[dgk48ZYW]S>22jfaaEfFF
k3MoR[?bl0?YhLXED>ACOU37d:3mngVn?gMH;YK3P_[njRcSnA=18eVn`DR=c]Bq
cWheB\k^Iek4_CYi6`>KY;H\dlM32Z_mXUe5K?7J6^88]6iSckPmX]FcSoPdGNTe
cShZXf]\KeEQT4P>DN2ikgK]^Hk9YdMg0Uen]9?HlgN:9B4\<I6LK6pY3UX9Mm0a
A>S6\Xi=Mf;i>@<9Za;Z2Qj0mhiXiLND[CBVMeCoGKdQlYH=FV_@>GeYi1GS2oU^
AcO\>j;I10_RApPFf]\m@]b:S;3f]DIR9IoUh@Hmnhe74PICJT3X:39Mo\eSM\G:
1>TZ=?90O7Dg<nPW?kUE?_O:4P]6UVHi9U>Dl541HESX\g`C^gM@iPH5bVWP<N2L
dPB1q<n]nmV=2<Jj<7Rjh98V\2Ia7W7eSRj@77f8bV1B\VV8NdO2B8L;MV3IdL32
bdf4J<M0hjco3dJHGR0^oCT^G>Ni:AR\>VQnD=fLgdZnSJUH=ai@93g<T]6plm:Q
UWoN3IX1OH_RMl8SmcbfF6K_0Ti^JXkqc`9LYE@>^RRdcbCe4@TMILLjUdkG\N]_
K@VH6<cAW1N<nQdANO8CS3]>dH>HnWfDcH]g53[aBR5MPVFA_AO4=bY0=MBaZgeU
<@PA`CBjFF3Q2YEfC^L2ddqV:gTQ_AK=<iXLjZieBF3bdf[MYQPOJDE5^8C6J1C_
Ii\:3h?MZXae:;A1Ke5CNO]V;9f594?K<S:VCQJ8^PIClpKb`l_j3VT334:b6SKW
bkPIZe<\jlEeW7`eZoTOP4NQO:fWfCNljg5ee?78>^j?RMKhBl0e?o5\bM`KQfk@
>^fcQNO4:JgUMUJe21n9_a:34RH4hJ`HI24AqadRd9DK4K_:dg0CAi^R?7M=lIK^
7j0LQdUnn@6U30:o`L?]58T6W[TChcCibEII:anYl5]Ll=E[If<jmSn5Td[Ed4P3
Lgb8F1UGEoW;Gi]EPCB5V6K=Vm8q]oY2^D\76jSMJE]hiMcYn[g^Bm59]d>T`i[B
d5BF_=Tn\=EjV6\dgNU@I2\b3Y7F]l2:@^Co9GfEB=5\^6P4@J8UH6aMOj41CiU4
^7l3IQAkQdhZJTmiVMpkbbTWI_>GX_UQl]>`m=c\[I1<c2\ZOU>_JX<R64KlanVG
fJ5@V[;3f<_DKeh9Nndkc9ZBaNEdlof7R8<MDHj\=q^T5dALG4K6LEbkS6gN\M:j
BDe9MKQ:Jelm>M^`gRBVFjdc7nM[Tba7q^[Jn;Fn_OCKlPEmOYZ6aM3PB\A]`FW_
M:g8=;2@SEC2IN44@jR]ikJ8Lm<fHJlMM^>?g=KCaUe?XEkC=KCSb5R6i9oKdg7\
]Eg4[1Yb6Ng;>0dW9_7ijO2q00\@`F6]S4_RWC_EDK]e>F6c`>EeSjZ59d1VTe>i
jSm1=BPg^BWA3eC91ann2Q>o0X?I>C^A:Tlk<?ZMoK;ZboI@AeNkoP<l^dg4G<fN
UZi?fYom0dcFAmp5hWOAYh:Y01[1kGCM?_e;jdCNOCkB6Y1LGF;X86SP1:Y[`hfd
\WdPGJ:8LlZCc`350J3O?WiTN3URXo5<HP<U88a94Ge=Kh6WG>9HRXU<Z]Z?9LTl
eKkVEp>D=B>IgGY8cSlV1SIc=]CMma7Y5SiZa9>VU8gB\BQN]lm@^2KEIb_EZ?KZ
@5RKH?>j0oXo18fM613oBnFLUSZnpH;Dc;=pL9T;^JH$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MOAI1HT(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
b4U^7SQH5DT^<5kH>h7;RVW7MbeKW3GOCG4F6OW2X\i??B4Iq[]WEXFXoKjnQ3\o
Fnh1=VgTN;BVl^N8KUlGoSUClp@SEPO[MOEmL0C2q^AJW\0pgS\]_TcUS4>Q=GKd
\0AkXO[8QdId1X9gcXpeeJ_OKfZHNKKe3UH:9@hXMJ]?1H8@67n8@p7c_l2hUEZm
[j];j?D2m_;]90bmhI5J7GpET[g>XaqhAJl:?pOCOgPJ9ZWXG1>AT=THD7XnB9D`
DW<=jaaW;Q=ha31YYLV3dG3gLXZ;n=dDP7Jh[WOP[:k7N1gX_mMbmZYjMoW;AN=9
UEARF`JWZAVGX0H0CBb?SUa=oeN=pP4mG9Q5TX[hAiMi2MOe[j3A\cFECOhio^]H
XBeF4haDhb1`]JCWPMO`B4@cJg[4LPLGH=XEGk[W:N>UVZk0eTmC=jE0\n2bX8]H
B>2][f\OWS[]1ETkIa7pO6J;hjHdK2XQ`WFMU=6RM=]?9M?h>Ge;O@<cTO1kb=6f
Scb6;SiZ7B8h]VAZDX^ZO9o?iX@Jl2M`2Ej:I;\:fOWW@a6IQN8;H@H\C:S1mW_K
__AM6D[iASpEk9<fhF]H`JY_XR9bQQoCFbbd_H3pb>CI`ll@neZlNnPkaK4MPD7J
PRBTE4Z_?8dQh\CKH1maN_Fj8Ik^MdeA72g>H8MdbA<S6W==`e7KcgOZ^nn_k5q0
OP:5kffOj6YSAU=8FK]bllcM[ZUR5P@O]c4IWUg=Gi:k[cm_O<cPJB3[[RliEPk0
PE?BXcS;j^YL\<LE[K[cG`H3KlFgccIM]Dkcac@iYmH=3=:HI5ag0qXiD2Rh50CE
oXbCaXagP_ZAPJGMD8]<ZfbPNjiB9Xl:@H@9U\GI[BJc^W:_nL\SkgXL2g]09_fE
@=J6[7>SJ`QcV@_RYF5>S<6P8m<KWkgIW:nQRRQLkO3Bp;>KMiL3nU;@B3o:1HlR
@22;SSh=lKb\7W:O3db>TD=2PVBPC;>ON=WL5mP469jf[;DcXd>=:b;dIASa?A9:
aQl6Y_FN=eTKTi:NP:ek8<mDacjg?_Sja7QpTFV2Zfj?TJcF<4hc7[F^m6`Djg6>
b<EgaZ0R;cB[0^W@DKJek\0Wc:22CGGHBlUET\6eQQWHYJ]F=PMQ\fT8P=qn?Q1I
5\]aM^R_;D61?hHj[A_`IlhHl8Qb`2GS;NJ;ZCKio`;0D0N^^HjkKRFYWo7nfP;D
JHglC>XjCT7_Hf^JOE1V3X0eT6HS`jj7jK5jI5Zn[C^kNHL0=pca7CBPGRUW9L^`
h4]`8KRj`45j:NHg:SLWZ76SK5@8d6=]hMjKFj4V<X:lKX0h>7ceXPPWnKWP>VY^
[8U3dS<[9?fa40=TG2^W?C_eB]Lcb\Oe8;JO8mbmq?=EXU>]^l:K6Uc44W^EA4=Q
pGM]^1aT;;IXFTY]_8\U\GGhUB<b5Un5;ccE=hA_H^9ML5KncgUDPmPc:;2Qo:9M
iG@B7HcY9\S438cCR4>WT8e`@EY2g;fco>cG1CBHoC=XE>[8[aTU=e@p2fc\O>3L
9=iDPbi0C[^lhi6nbSJ;CTin73[3_NI0RKV5EUgH7;Z6n1:B8=NP@6J[2[07@]NV
1IJDIK;81a``3Dpn8<AA?o0mPUWfZVBkfe?obM:@U9\D9GKR>O@7O5QGBMnM39BR
l]mWbak2:Uo>_X3ne@e?nVjA0Jdf3Y21g>f69lkUHl\2TS^E>GVhGjd:QC\a<EgJ
JYckXqjh9MH2\BEHQd7Nk<>kRXRPMg_c@n\ld=9RWF_Rb3\L:1Lgg_N`:hUNL=WR
HUD>=Hj:kZ\<iK_h]5@Hl7YVEA7nk\W7NO51_JQR?OU9bVSR^1PZZk3\dkH9q^@6
hCI4CZmYAMiM4FgFVM\6]RCH`MIe3W2Z>7XZRGCQ5@5Ak9E]Wb_DR@W6lR^J^^c:
3O2?[CnjFY4aE\>;DY=H=3X060PV`32ZXBfnG>3<NA\LJY6S_lBpdFJUI2RH\adF
3TTfPbON[>c^QB94fR=BgjRLgF[NYmN0cM5hndNPbVXg2^U\LkL6d8kTij7lSG>c
=VXZXCQ;lbqalV4Y4qJaP4Cmnf8NceKHPfWP;4dV2\=J1_YN^OPmblp2kNT>`W$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MOAI1S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
P]6kDSQ:5DT^<Wa:3aaf9A`Z0J`9`>KW@Bnod]C`567S[575@D7<Ejo4GBn>JopA
hCB_9S:\?Q\:25Y7fZ7UoGe9`LSqEGmTj2eQb>GRS6VYUD3MV?l:Y5T2CB^U4^X?
:N>PF1:4G\9lk<eV\b;gc\FSd?@pB`<I``pENBd]hc1??AmBCa:ekMcY56_S[1<=
DkSOXqGGJJQZY6caCnN_SN`Xd9d]X1k4eZ;WcS0Cq7h7U9Ajaj_dMh[K:WNbFXfj
<Dm6oil5Xq0S[Z?`@qD6`a]dpU3ZhA:JA3ORcgdPC]gPa^hg@`WU2^aWD6__DmXZ
3?6FlP5KAcI\la[OT[O9iH8\TUkeGO;N66?dXMX^U9S\=1?g;\hLl;Wj<n_Z2_GU
a;Ok?gB;@G_hk8Wq\B]ZK_mboOc8G=aSFb:Q;\CP<G`]d`gb6U1SW4fNS9neKUIY
R]SHBkk_fA9DJ^OC\K_4>CTkIQjW9Gb6UJSC1:nFN1Cf@Fc1QU<50V<91@mk>LU<
eNLR\bqnc6aMXOS3Hf<e:\8`dB37=`S?2Ga=1Y4HfN<4=QPMUR4jMeI=\GfaL9:;
DU2hnFknh8A01n@`khD`?SP?cGX_K=N@2>5[^?g]f7lHj2b<;XjMg?e=9d1beqO;
Q8Bl<ZUT<9\]LZYaJ[`emgSa<:H4nT5LoTW6qcMM^JU>DRE;<c]khE<]?XdIn]ZB
TH=nI59MBOHaLknZ_QcdfT]3k6]@immkm6ZVkc]GF3>Lm3:fR75^C7TebI6qCIJf
8]TA9FICBc@k@fI2@niE4<l`LA1=6LZP]@ZLeahGf1?gPge5gI<G\5A0LcG_Cf6:
H1bPWbl:c8Imi]Dm^RMG5`a94OaS9L_;EX;G:I\2@8GL_1T9mjq^6?LBn;A]U1bH
Q^hC_e7A`gmhWh4;2oSD?^jg;S>JVnJPjX:i=CjSed\2ZY>DieA^d5^o9IEj;`cS
k]SY_ESILNQDi<RDP:hB?^9mdU@<e?\WAYMHo@9clqdGd@oWe8_BDD3LXeG<h3;n
O<_4pWW8O79W\493ZF6oaa20Jb38_^g_B:C4R86BlNBk<8gmc3Eij1^n_<2<[Sj\
XllT6Wi^hU8ZERFJAGIm3aVd16[i6XfUIm[P;D6QiBHbV^J`;8VGWQaj]>^p>o?K
d1QCEY6ThFKgc;k]Oe:QF4dAD=:f6f9M\X7;1Z<`@fOBVlVPkImmA>DIDhVV>A1K
`3eW;T\>831Nc:IP::pJ]A8BmhOkil:XD8d><4PgTmO>_mal4D6[T8e`O7J441jm
Lm4eE0>FCjd7_l>^mimJTRb_?i7VPNGjiN6KWAGDLO0;P6E@<aWJT1PO9WKcn?G2
_4ZWgKHE2pNYARZB`=IjZVTn]U?8ERnDepXHF0\J0O0MiMYi2kgGcFBm4]^f:;^S
gjA`^`b0?35f^;XcmJ]SC8\@W?F2YO^k^CXB9lcobKOggjmFjbY;3<2bH<LS[L6F
MdV`^C=;UO4@0iSZWM3[af17p@?01bGDSQ>L\61Q^^cY`7bM\2i8:J;Vlk8d4@j<
K[bSF3MWoJMn^U:2Ql1L:F8oD@7[_aSC\NC<eP=O\SmM[g3D]UiZ\P?6mo8WODIM
cW[M^9kNhG6@DoMqGOmOE7m8@;K1[oCLJCh>c_IlG2:GhK9oThcdlF=L]d9e49Ye
_^k:I>;[a<mT30=aGj1>7;K0ISoQ5[JXTh64=lqDmW0:c3Q]`;Dg8Nn8V_JWKOSF
?@FLMQ`RUZER1\UWmc\bdi:TWPQ:W<X>6Zh36KeDoSBRHc?Snd2hT@MDZDje=@UJ
`FD1\TI^UE@ZRHUESG99Vm8Wo9XVmpM?LFmYQ0TD4oJj]7flVnfk>gnG85dfLdSV
eVmRR]C;4^R2T_3D374^R01T20_bUhM>3Jo27eGT4=a8n01VPXLMd:l0>\:0Vl]V
1h5N:gVDJaI6EU;So^9DqTTGHI?@kMRRKbk1]QIFeZKTXnOLBPJS_]EWhZmo`e:N
J3o_p02^jeGI<8>OjPB_nnn`U=oDeB64[:^ZdD9EOjckKJQ2HKjHTK5_4fOJ;Kno
a0=Hf011?k>6Rg`4_Cg>3B;_L9Lm2n6>DW\M8c9QY<VIkHGaKIEJ3oJ8C?cqM?Li
ED[:<2KEAa_G^SG=f@W7WEPjXYjUZTOW6kiSnMg<61gBJi`4USeaR`W0Ab?_MnNb
=9VYij`M_GW:@_i\5Xpj=1m6\pO54bL[4$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MULBE(S, M, Z, M0, M1, M2);
   output S, M, Z;
   input M0, M1, M2;

//Function Block
`protected
JKlCbSQV5DT^<YMl50D56d2A@0>=_nH\m<FQmfbnfOJS9RWa3DV\D?oRh`XaUa1`
NVGbiD0E_^7>pR[hWagLjA^i55eSE6c?Jo>dL[i=c<^?]\]Ih;^<RdGDXM0:Z@<\
J=<\HkcUk8L_oDme<<Yq24b47^nKM^FOmK^:1NXo2N5^d_kH_ITDjNhC8^?oVS=Y
fadhTRLF_7S2<lf[Amp8T:_6QpINBU4?q`^eb=@pMd;GT@pi]nR7DQV69P6WZTUm
eG8DG6OQell]OdBAOpX0Z_jC9mPBI^N`I1gEDcB4AkLjpIH74Y`8X746Xi\A11j5
9m@@T17Bkm`pcdTLQ6NOi1CW26`o@bh>=Z`aU\P:pdV^62gYHAn=M^FCI2DmIW;b
i;i1;qOZiem45o9YW;D<mOCjTP4W2JL>bdpO?Yf@?bTZ^LM]_034W\P7l?Y\gZ03
Kj5C7L<qDiSWj2T\QTU5J;OI?UF>]dS1KQnnPBSZ9D<4?9lXg3S]ba4eKhKNhP>g
poBW7n0nK2^F`RGG7\XV0:Nf?U@n1SQ:Up^09QkflZPC[I@;KaU]5\Qnaa6mfFDh
_:Nap3dcAaR`>;iQ<bl5=^gin[TSQASA56H2R4mp43OHlO^pLeF2R=pi^WVV5F\=
=W]F>C5[EWnUHi8K9ZM2VnSf]Z\5=:lCDnmTaei[E8Q`9_`[RT>B_Z>iR:@8Q6[N
E25336UN@1]I`[b7ijeB_8o5]9DAgTA4:IZH<II1nMRIbpH?c6[<33Z21hcl?[5A
kROQ;1Q[?A]?PRoCPBjEFQ`<QThBULBB?=eG]laBZCQ;D1HjWC@]HC5P=fEm];15
_lm:4bPH\iRk]l4CISQR5AE[m`EU^;XAdl`WpCH9_BfboJFo6;WWGnAmQQ_Q9=Ao
H=A4]FhZR9cmATT]e1]bP=W\2ACGPihoYWhUmC?l?ZJ;?DA3K<j\R9n3S[KUagFh
A2oZQRhBFIHmLJEg7YhNDMdNm`^p3VbbCHoNTC3;dUMMWalq_g@[;_`OClK;=Ica
naBS@_;E]A??ijOa20WYnJD[el`IJ1;gD;ZPL9G?DLDB[XlK_Bo1EnmAfWBJb7JY
llGYE=pd8<WVDZ`F`bW]GQ;`d:55hBfQ<Zk?gD=>GKeZf^d9P`MfIloNJD3LTkKd
bMMH2g@dQEAi8e^e`aB]bg9DT8YnjIBLn20o9[J>G:Z@mJa^0D_kS7GNDKGZBqFG
4F:PenG=7`Demc`:GcT:<_0YX?idehOFUk?@9bNO3U>aDThdEZSb=eZ3kdaRXnFn
Yf42Ecg=fUEaioLobUKfbio7iTYc[GgFUn2I8KE1mYI?M`:fQJ:dqUC8[e6JGRYO
PHWoLlDQnkD2h_fAXY[7kCFnH8]UfkmO>ngW2OTk4QjkMFVHJiZQlULN3]YmJ<YQ
9aK1M0dG=KX6:HJj`<f_M6FZBkTVIi8YMI[`W2PMc^Tq7]LFJKE9j\4o=QJ4n9ZN
BOm28?nC4iUCJ:ZH@MNiCiZQa5Ok6d0E=NA1Anhj;02g70RbIERiL\b1V[CBGCea
ZQqBUeFCoZ^LmS=@aNT^W`0N5cV^BG7[KOf5\B:jgg@kRPImaQ:OLUXj<WSBgbh\
o=VPeG6pY5^j_P]mf1m>@Xi3iZKN\OQRa[0@jJ;D@S^^Sl<hl]AQC\F<77bg5mOj
S=EY3SAB01[4dcDbcS<oN`nYXfTWZDa=W[XZPWG;eEIlg<FAZA95J2q@^ToKH3NT
9?LkJkDYjP908QcILNoS5No4PN6=_?n48ak429fM>8_3@Te33HdV5_^@7<QUMLaP
l[o:QWmCc>Lm@TRf>oHm9N_di8M1Hp_M6RR_HKU`bM749nS4ni@3O^KWPINoOW4h
d`LklZCh[OV23WV=NB9hiGDX>L;K<f_7kO>`KS0Mc4C@=`M^\<`SpINkcE6:N0`Q
?MO_AhbSVkb`n7FF1q2]oICNcbNNUS8DLEnOJWKFb_3`l^Il`8SDkK[:9GZ^nH>h
T:ZOjmP=[FiMDjNQUScQ]KoOJg69MI:=mGR5_ig^O`X`U=`72?=Zo7\`dM__d^VU
qj4P23c]P5nX=gc7NBc[^jAA7_fPiBb3Ab6Hj9ngIQMeX8;hEML31Z:l?CaWAd\b
_jnO7h7CFcXeg0Y2jjH?9?9AEEmmj<h31S1BJl9q21@ERWH;N=<UQ6P0SMh1c3]G
J_gMNc^VAco5SXd3?C13fnaR@GmT0<oUOhKm5mi_2jQD742MciR39n?IRebG_Yp6
TRb]mq[TcW:<T7f>n2oWA]9iNgNNPbJGJO8`18WK3?Na`nfTcM3jGodEXn^533U4
MfVUPJjIWnA0;mdlVo6Ek049`@HPi\V0OpZ\_Y;4ZY5fbQK@Ph7mKUlfTjd\VCkX
`G1T^B@M;CH=aLc2o<2M[IdQd^KCkVTXUeKkC;QGFTmJX0UHKVgo^:Y5]Y5K3q6@
1EGX[bTXA4lRT?\C08\e=0`N8aR@ZX`IH^[_EM<G2hnG4dMlMdnMPj?YJSd70M6S
mET6HfUGo[BGLOj1<pGSLR2@>CDb]5Q?kJ7XVVB=K9oH7afXg`\jU>OM5h>lT8D6
Y@SJlH9QY=Fke:edKiGTF1HcVN<TdmO8=4im\q:8VJGJ`$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MULBEP(S, M, Z, M0, M1, M2);
   output S, M, Z;
   input M0, M1, M2;

//Function Block
`protected
NQ>EUSQ:5DT^<47RDoMO`7dIB5D2[=q05kAQ7Y8cI;RG\O<3fT^5C55HmIRhoe0J
I<h41fQdB<`O0eQnNnj0RpdZPQmkeA022WF[2Pj[VGV:[S20qSHo6P2pToAWNcpO
mBfEnp=;1VS4qdh0Bb;Zdj\g_h@?jE?fRVSo]g?0CRG>^01pM0gG;ZO:OJ<a`DQV
bKDbn4hi\Qq1]IZb_A=e`7cWjmHljA3\]4]R\Cfp8D:<c_c60MaW\ZNIeiZnN]LB
LSoAq[D^gI]B;^TGOQA]=JN_]OLe2JM?\qYlDDW0[F9g1jlh]P9g3V1HfVgc:WEG
npGCI`HG<Vi1oCg]\T?QFYbOKjFfDL^7Za2<8iplm4`nI0[c8l2aa1\?IfQOW5:E
IIBMjdPpaUe8>WlBD^Y;kZ[iMBiKiNcciXFGgX`5UJp>QUR]d@C2BZNfDaeQ228P
>WnlIPomAjLEXpC6`AM71pOm_:8a48EQdg1o:ihYhg<F>]bg3_dnGe^HlYI7h5Df
31pdl0jDhpIko81Q9Ta2=f]OZ>`2IPFJggNM[lEY?9HgJKg;A1O2;4Nl0ZE3[kM<
Sc6g<1ZHNGaiDK`=]GNeIIB7UeE5MZ[Qe6c_m:fSOnCDUM8;3[e<EVSD\kghXIBa
GmcGqC=8BX\B2QZQA81@f3knVfmCdOhGC6m>U:1fQOU^lQd>]8ZX\2PN205e3ohc
eMWk77I:iMU[9eCNmR77L=2^bUV=d\?QnnchFRNU_nU@AMlRoc;c8XVPYU]JWPWp
9eeVRLJhF^WeE0hnOcnH4H@LV<Q[\EZoi;E\IX0JFePLgZD=Sd[aTPl?]BXgbI4=
G?=Zl^_f`48Xgh>^@l]lZKcV:nBnf^EU5\h?nX9@oNa5fAd]JU6YNQhNNbq7lUMV
aXo]FU5jIp:4n^NQ8Anf`3X>@j4L4E_bI^en2e>K9L<C[Uk6Nh9aGKFog25NBX7H
k6YeY=d[\EO45WeSWg>?9MFS9j^FAJZfl:_GqPld@@LTBjZ:mcDTY_H9V5BWG>N>
l1VU`:H6ReDCI1K@XRo5SBO@Bn?loa9YiR_cmPoh]65[_g8_KhGg2jPGVQR4aWV:
68giQ`H6UfC`;IM]^DP`BZ75<B?qkOFm3_`AERbdkBf>e0<BCQYc[LegXSUlWQJ>
D32Dgfo5_CW=CL4MFW_kon5;_CohknQ4I?JO89_=H1=BW]gR1LH9HdY2V_bOBQEL
8gAdBjC7HG6FfeTR^[qoT1=i0NIAg5`]6_XhcV1gIZlOPW0\K2RakASf_RHGMmDn
b?ecI`i^doVUGQXV^?:oe<BNEglMSgYVX=^lUV7SX_mUcJ[LE=e>kbSZ52aW1;fl
j4MD=3k71p`eSo8YWKCm8W:Snil54Q?Z_[7H;dh]WB6bV9VEjTl[5G1?NBSU3WPB
M?>mXWQhLWJNUaqJjWNnci>;<PiDjDWJi`c2jQ;fY;ESB4;A@TJaiVQ<>a`_?XYP
naNj@lD8]5Pn:iLJOm^BDmQjUEP_lTELO1:O?pY^[O]4>7:bja?>4^XRh;@9C1\D
RoaPXoY7dS_PJUNfdfQ2X=Gk7KX79n=V7dANAWL4N\WFWnXbTWg^9jUMfAB4cWCD
;gEkDVI8NDdSSJYiNAo2p[@Ng?NG\3P8X[E7<mcFI@<Z5ZRT?B`4f70hKccIf[n?
Sg7]>@JL?N`6L9jI2JhWMCe_X8_eCLncR^F:YV<VUEM1=TRRRP[JL1?\P>0gUG52
iG?pJ@jhd]MBF7@KeX_llmhRTT8ZRKe9EnLIAC4miTQjEQ>;:FCcVB4FO8@AOoc4
A4[UHVM@0LCMYLQbT^PCP_LV17[c8iTREmp@@U^Ib5diIM4@Vi1J5Y=@K1j8FB?X
Y=dR37`XkQ<mDGocPDYGP9aOd]iib^_SYEldi;P<3?maXgaD0Ye==f03B<LTFgkZ
hJmD]c`\;N9;]]6c=pW:SlAYnimHR9ID=5NB3od\GO8VHDVagd_F>_cOPA<lichc
N<_Yod3402^QdC`ekMlP1::9DCb7HnUF];3B9?;n@=7VKYebO_D2<clCMoRmj_=c
pGBKaEneh>WU==WhVZ_SH?b0Db@V;Jg3=AnPckJI6cb61?P^^Q\>32lhWg<8j[`4
MaR>M3Cb\WckofT<QB_[4I82?[AB];>p@MJB@:8Q``YQk[jRq;EooDNqPUY6CbfT
K;aoOATCMn_>3:]QK6EhWoT42<7b4[eHiUE1eBg>>K<Jgn^SZPgQ5=7W5]o05eOg
hXH_=i>M_kfX<hGB\43pFYF6LfoSWa[Z`?F:EMkPk>b4iWX=DnTY\nUdYT]WNlPP
X3`YOLTYQ0Kl]a8S8akCaH5Pbn0X=4Cn>6CdP77l3hUl]QKpWNfHDJ:hT6=4RR8?
HH<k`3Lf4c8ShW:C];53UTQTE2J[[ZoKELTLPW:2J8c63PQ8LJL[0?>mb5l<>jh9
`M^DFP@qXb>CDIaI1=^]5V3la1H7g_OTVJkVg9Oe8@g2oFi<j8PoC2ekFMI?A1Cb
WPP1X]>:`K2n?R_[>3]i_\26`B[Y71YqBLl=KNj$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MULBET(S, M, Z, M0, M1, M2);
   output S, M, Z;
   input M0, M1, M2;

//Function Block
`protected
`3TO:SQH5DT^<TfK_Q\PPYG@1WEVH469O[JcIdP5`fop9PXBFLahZmYH1]mQ[co;
HS:6Ieb>gAIP2U[]54ZqIZcEM0J\3;DWTa>40Cf58EH[EiP`23TcVOKcNWS8le_A
e3D[7b:0jQpol@3bDpHcCoFbqL59Hh`qm\bY8Lp1Q^XT`oQZYJJBcF<hN>InL1kB
EU;ggZJ=8q9aJkYm@?L3\NngWE@:Cp5adakM]Y;n6cd@4a0bLA=X7F^lp?j;L1CC
A<_ZJ]fKLEA6_Q]gB8E@FqJDAW]BJl:DR9mnDD[ZMiiGW@1BPDqJeY]6WmOjI`M@
eeKDX;oALOGX5KWq;>[=YMDB5ic^NC_pT;2i@F_;UWHG3UJh=mFhk;oGaLLD6eVf
daccqG?]59oDMlBSW6S5^k0[m9l3Y31?@[;\:p1F`h23MC0HV]Sil3ba?UFVK3gU
GhP@WNf2qU9a0Xg^U>2\Uml[mPNOSKZhdA<:1_^n0g`qYj[8YX\qELmnhlqRHaD1
T0Co6c]L2=og=0j`GM[A^8hOgH2=VeI`ThR6eFDd[fc`1]ki91TO485BNM:n<LMO
Ve709iehEB:oD5OSj62n^8iHW`FK\BLTYMfoCKVAVb`n>WVV7616jLiMTq;AkQhU
_=E?QEPfob]^i\:@GGCBVKaNIhd<qi3H0NP[\aN3:S;dbDTGne4YSa;MWCVV\[XW
7kPW\^FajnFEiKM<S\Jh]Y]>37dZj2?06dhS8OgNW4ZZYiI;Ibf\C?;UWIcB09F^
U8g_E_oaLNjdNXnk@FbkOS[5eaaq>V1mG\mO4h<@58d\NFm@U>`Y@_kSoGdD1IM<
a3K7[nmBm::bc]kgcle27e9il9>TU3`Z;EI^C]HJ718:>S1O3:VJS_]Q8?34oRW6
W8QJHOV5ELo;Y759G<Tck7[db`p7ElS\d@\E]?V?Ymbd;@D\^6YKn3_M6n\a:9FS
^lA66E=RZQZGiSKkj@gN\>oRCDg\Rd;g]Fe@`:fH`G4V1DDfXaAL7FOc3qN\gNcT
\j?KZ?@cQHDGj33^onmYGg>TJDL`XRkG3X1ajiXUZ09?B58FFSkGR2SZPXNFJ1\9
9jnJId<8kCnckgFNkh>jT?FmNEK`Fnl<No^j8G@IE1RD>1YUpUiB[]458LL<PA=K
\SUQXPDV:[eFT]7b>CVEEkd>Bn<N5V2bKZl@;`7\RkoAT]ZRoUc\Md`=0m[KWOS\
^hW00GQl[1<gYR^Ic7VCTb;6bL<<3>L;`9M6m2np41cWc96g?@=>L_eN[O2leciX
GKK]o0\?UbT7D]Hg`gCOiWE4nd;S0nF:o\KY7EHo4^PSU5:95\KS2:bW9k2CTVNZ
Uahf8:2X:bE5AP?OQED`RiU:A[oceeqaPXa2Hj:d9Pk_ca5m6gT;[M0FV9dHc:U3
S96B3VAXkZh03ZkE=PG<Q=1\jJ8`[7<a_X<>Ga5gL8K8O``<J<f1bpiognUm@MX`
ZFDa=:A=SHmoInTjOYMIK[XBg^`oRG6W92n;e0m0T4UTP@Z77pmbgJZTgZRMRi7b
LmnL^=UZZ8jA@OLA5OR2R09jgW>c`dhE7CCR<^VXYj;P3W6?F]33`e9mGYPZK3_C
5aPW0WMNn=6AA\Q5_DcNNPnYd^eX<EOmq19L<?7KMA_OnPSN6gi2@[n^5i]:kMCA
JZ9lZEnA^O4ij=h5ElYZC]R;SMfBWa7VKiOX[G4g1TVZ^il1oCiBW^2e_Z]T7Dh\
f9IM1UmC?GZW<3Pp6jblSO8hka5U88kI[cOcQE>Yhi0Y_2Md=gRnK;IODUl]I]Ji
0NOF2QYe4?E9f7;bKcVVm1KHHEOT7T[Zb4fR;[QUJCT>`TqOP;B_<Uh8NTm83QpV
B4Dej@7keag[:>Wm?EFd<X<\kI=fmDj0CBR2RCT1^dHV=2L19hb?D[?CPk]Rnd2Q
J7lXM_GOFVMUFC0AB827d7iak3hREKLRG0hgWO=`19N]<p22l=O@lGYi8idV[e<H
T\MUGR^RNTnl_4MK\]:V^UY>Am5WEM<[2h;Ib0l3O?c_8^nSod4[QLHT^Ra?CQ=E
6M2aQLARCR;@hfNY0TT\\JiX:gP9qhb706VCMBe=KWg4ZNIg077XZSC8X5WC?7?N
AfWd9YTK7l?E>4aDA`3SW`cY<@B\P_EcSM]<d05gVKdT`SdkYUHmKbW;Ua5p0c4X
h6qLO=lomhKMOQ=kh[^PN5VFNbobF1Z`DkD:bcb=@K?T_@mOalAgWWAC6`0j\^MA
SIZ>[H_3`kDD_;F^0YVifP=Vm^S12Bp=]_iUG0gJk<Y^gIbl3M8jB>7hjbMQLQ<2
`bnV:YjnERlSAfG@>mc?g>IcM_Ydjk7:V4Z8W]8EVc<B<X6\7TJSEiko;=pT@S\n
7[ZBaJLnh7L3OhCV1G?aGNoZX\GdOA2J0oX;RggN9AUS35Bagp7>0YGOo2JaM0UW
ejkDmB=9n_7SE5c;9UE]DEWgc46[_<IfkiC<Wm=NfX_P:`C@6Dmkm^;dOEHkaA5P
40MlkNAKX=XJ>p<mjViL;IdN`ghEgeCoZA_<__ag5V0d9iELll7fFEk:R90FZDk0
6E3Y3Z096=>SD:2o`676[YjJaD2b?5aoH_LZOcDAop<OUM`SQ$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MULPA(P, S, M, Z, M0, M1);
   output P;
   input S, M, Z, M1, M0;

//Function Block
`protected
A9]1GSQV5DT^<FTK^CLhL13Xb86=lO`MSZMRH88Po]jO_llEWe<f4di=pNI4`FG=
m?]IQCLB`<g]7h_jWB`kYMSNJfh:5iC`6WY0j@LcWSU\R3@h_qF;NEn9^gMef?Go
LKBUg\M0gM@N?QLebg`<:5^GGO\:UL]oJcTge\XGF6G>i4ZI9>Rnpg@Km:7pbF1g
CHp_g@[DBWGC8eMb7eVffHDeTb3_dpOc_FiA=CbIdC9E510_g0[d]4Clpo:o;EXA
D:8[TbQoelfeWfXbe91p1BcM`4iSmDMcF@i>dDcc9I^IDL03qWm]:0?:4[e2fdUT
Y_kDjmgnGmAg1q4X=BFEIG^_jS=99[ZY644mdnI`8cDF?TkR`qA_PY9X^Vfg8A9F
odT7oIIdET@Hj6oY]Q?U5EEi9q\_Nhn@=SbHQ]@<E@Jl_^6NKWDK[d`b29BP;kpd
QQaC=Adnng[QSdXT8cLjPQID3<2nZm[:bO9d<p]Pi[1F[=3O6TDJX@5J\Fj_JQA4
k3?n^ObHGq3EQHJCf`SaoWdi9RYe_3Z:9E5_<B_4I7g9Pp6BN<gnBHHC_bc0Vn7i
0D]k[jH@9bc_boD2KNp02^j1]cECLNjkoN2mW91io__37e;U9Z<1;fHahqn3HWdj
GZ\5eWobYLTeHH6feQnC2jTY7ofAnbp<0V;<8Gee_AZh1UaiGcgF=cjUn3>cPG1G
:RqXYKhOF[qM5?oK7B?Ihc_5S2<TBI;Og9o_N^nimo?6DODBLK_iC87e2SnTce`i
B<]f`bW@@^d>hT2qL0I^N<qC>BACFc=A=9L1<IRH0jI;OfkeRc`==263b4TcI2_h
\QNCE@AUjLMj58HOE_i;6[m2_c0cCTXF=ZU=aPni=b\i=5hGcKVVHkM33GXj:j7Q
F9:A=l0hH3\N_GX`gCoS=>kPJMM;CE:BeHFFaJml]S\[=5Z;lpEiRo>=04:>X>JJ
n2DG<;mJ0NLe2UM6cIl8S<LPR\^^T]eD0@95COa`\`4Ok5`oiGC?\T5N1937iPCa
E[HWmVTQk_\QjIZ6_1l7doE4=liX@jH0\aiSm_d6;D35YfZIdohIF1?NB9aL_Ila
D?JX>5jQ_0WdqnoELme2hKXJ<4>lUg;Mf38HF_3]WMKh[<43<lCGa]hW`<]UQ;@C
FFoQS6XfXBA7^cEglW]kj^d5`T?I>Iln:]Kkk^ETmD>OH<S[G5dCLhERaGU3032]
e9UPEJ^n7IDfREKGjo]W?kCB47?V0l=c`]KCfF^qjQ^9@Q6V;EYocS8U]a?Ebc^T
<Q;WN8PkkI_gLbESJaVf3a08aA5N3gOEEPG4HV:i9\Kn>MS1[3A@oBL;1fhj>3Lg
QjOSMJ\Fk708HSgA5@oZCJQ\]`UoMiRc^G;c35oO61:dCM>==G7AhB0=^d0123l4
aepe83T24fb>;Kb2;?mY<3C>:ke5iXZ=D<2Kgi8PjIZ<c[R6eZ8Zg0aRnT\7bLm1
G^l<^Z?omW@fKSPB<NEBB[L8XcY`Q_nTcOFKWj3LXLh>Y28mnG?NAjEPMS5Y2\MP
05gO9nl`mc;3QR]5<ZSnYd^eXEU5mpVg[<iJ;hCm\1S7JL_1_T?jQGLBYoJ9S\9i
[>cHRVl=Sl`b[U@kY_M2K@YCcS:0bHXd0hn4jQH[^U:FRGA<8J82]7@ooaYKYY9@
@FokdcB6\Hl7h\amBO1[I0L?QAF10;Y]WC24ljW3;0VF^EVbeFo2fFD^pNf8Hf@S
FKO1nNU:UJ9cQAWY=Z;RHc>ZNeNUfE2^LjZO7mLFC24no?4UHW0Oe52AHDY<i5lN
<aJ^[YHSCLl[HQHU_kX1<VWW=eKl[==3mLW^V`0cGXX5>E=TRRcN`noXWJhlVMlK
_=>3j=HY9>ZoZGHcLn1pXd=4]JH7I07nAnkBOmlieJlBP9?h6ZbPkRl^jEmc=Q<l
BS^2O_0`0UK<QDcGDcgj4<b8T4?Ul;UMfc@680^GfV<S6K1Cb7_hkU7\Ll_E206H
^kSnf5W_9h9f`BIOaQBQTLHC24W2^hhiic]J2N?L;V_f]Wp3^9R\G7<iU7k5BCmH
UA[LK=PSMF0bHmUie=YDi`59KZ_3LbFAJGUTiq\ZjKI]@c0j8[UN7V;GNTPiY5J^
;KED8aH123;P>]W\NVVVje6DeDD8mT7J]:i4@_Dd2DdSHf89_873k_o^Ejn`>gNc
deqYK1KQk0AFKhPbL7OWClT1Z7eLb^GGlBGZ=PRAJVR\39WbIY\N5D95h6B;:W=L
nLHk`;Wf2=:eO_Ja17fOd]4LCJeC^@RODE8ZIglQV[<UV2RX@Jb9?jL6:5A]LbGW
[ia;GiRl2cOX01E91?H9?_e1C<D@NpE?m2\04TdP6bi@>KKef?FSFN`<^`0PkQ`7
kjX:b:>l\InBI]29W8d7hQSaBAoOH;J=g^DGhi`AJXHMXZE]cS16F_VG\\M_[]`0
7MEiP88lGS6Cf7l=RP:Xdi6iAoHU8E>E045GZ_LW6@DM]KRoYoE6deO1q_0FCTd9
H8_[@M9U>I0KIRQ18WmK0[T[a^\1VfBeP^hl2g`C=OMUCEhEmYJHQE`l_lHMXGOJ
J2YF9m3G;]ak[1M>L7@8F7KJe^n[3BLCiM?4F20CTgeJMKChNc6TDYD6?LIkbJO@
>4eKIS328l_bS=M5ELUpD;b6C62hbk1TbF2Q56Ca]2^RM`C@>@NP@ZV4cY_f[7KR
a5m:4^c?E2_enehnlRIJQS7g7\D`5;oOL3P@P\TkNGfM[CLV?>?_@5FA1_Z0\VQW
E=`Kc>>YZ1@7jZPo\NMEQd:AQ\<Ld76`O3l4XAX\RGn\Zeq[HRT9UQ9\SBZb=8HJ
2B14n7=OUJeWmX@fLEG8ic:KK[ii6Bnb<6C]mKf^:Q9nLFD^^mi\?BeWSO>KK;3[
EaFS<0WWeKMa3H6f`<7Vf6b9Lk7:]iMNMICPe1kUAmGaKbQU_n59?Zi2kJBMKB?X
G1?S<@@B9qQRnY4PZjV2]lAhW8gF1VICM7nHan?MY9=SF^e[YDP:aofjJ0[d<b3Q
d8B9hcFfa8IA9R<J3JR54?4?Pco=ZY98ZXUa777BNB=\gR0dGiYQFG0PPB73cP_7
m3X<j@L511f4?@]J`J>chWe?38nX43Y8laGoqRb=ASZC2Ie\Pi55mp@fe[UEhn=h
Y8ELelhJ64?Ol;A;8NQFlJPMP2OPa6j4Af@Qj6\NP=D7NIY_@>@n3biB^]=Ld8:n
4<7cLINT_ciOAccImL8SENPf]Fe9h]D5G[_G:^CD]9aDbY9eS6kQ;n0>liFLQ1O1
Egmc`Ff2IO[O<a@?pd;kNl8V^88gB8NQMkk?@G^:TCDeLU0bH?@eZgXP6mjZ4mO\
H6mGe==0Lom[GHY=833Kg;ZLY5N4Y`<1J:?jgQjJfTa6W9hPE?ggSILf3X0U3\@M
73b;W8XLle0jd]ZO;YJJJPZ5k`f3lV<EM]76fgj[VHVqDoRTED2TV_V;X`@IDRg9
K<Hce6ZSjY:BT5Sa:ifTC1KD`iF3T3KFjG72k9VgfT5;8<0k]Oh=5>NYaN8Mk[Ik
::<HKkUAqUl;\SEBD9cPeiVoZ@lO4o5?m7=@@?nO?X1o2ikTdG1eF4>Z8n]3=T8I
>>m[aFBFUTDo8E47XHS]aa3__3f2?R4WoX=C;FA?k@[fUL9lO0m=NYCje4[2P4EC
PjC0TAe^6gIdKja=IdOCqg^Ab0YNf=k;UQ<Q60fnFJJZc^9Fi2Pnm0bH\8VFlNYJ
UK<52\26BZIRo<W3L0^kNeFQ5XhR:6hVe11[_AB5m^<EX29Yf4TR`VLdLIiJm^MJ
^dcD>X`_iWf3cJ;BIQiAS>A5XXkg]b1hpXJKDWSgQi>RH8_39M19:3=J9Y48NP>l
9CiA>?ijQqeHTW57\90BEN;T:@h:_Pl`78h2]E0imTXERj6Cf;RTAB?b]mAj0W?V
\[Ud9j\OPD7c[mQ3f?ST?Qm>DiZko^K4AN?2@1>YiUAR8dTIVgUnci`Y9jKgEHSU
]_JA?7hJ9ge1OmX9Dc<lIpRi2]XGADDnElFG`HEMY6309e>;iY>=Ml;g1FIC>i=F
@kI\][o8GSKKSJX:?O>RJZfIY]^k^CXBXTcobKOgFlmFjbY;3<2bH<LfDG6FMdV`
@M=;UO4\[6dOW]h3G:@P0YDMGYfFff6i@qNCfdJLjGcbg?6O27CHGNNjG@?hh40X
Ra]DEL_UO3@1Ci471>[hGUNen0IOh`3AGlMhX:ILBb1a<\VKF;YY?e0f]C\6ET<a
q1]_O1bkI1FLoSDD@S:\0QWm3deTL]0<OE^?:4D6QA^l[gF@K7iQ564f9EaCe\_R
k1K36m26oM>Z;f]j\YCkN1n6jdle0jP<dbc6c7TM:mCMXIGn]1BO6Ff3>>DVQT_H
9a4O1B2AA7c37E]Hk3\poggMk[Ko:7VVK9e7iTl`5Ind8OhMp>TlOo[LboPSPn0R
QWaF79ei:Q8`VO3Cmfg9aa6:?^^57f=Qm5<DC\RbS@f<h50^a>k>B6NGDk=MO>a8
_W4U1ab82QX:@ENClQ?@F3_UBh\]V_FZVfNnQEJT@22K580QR=:AZeN>\A;Cb2aE
7gipfUk5KJfB6UbbEM<olESKa4_LaI8hRgg=3fl]WZ:[Xb`jkI^\[;dC05;lb:\?
O^f;f:DRiW0<YPfIIZ8C7L=A<I@Xa<TdiSg<<fnKH:B:5S7I2>QSHGE4FZ3OT^jA
N^_Z2\GJRWm[Al4[KZeP7bp_Bd6Y:[lAOi]3a`=CZ\J9ElAI`1`;]NSTPjM:h1gR
OJUU7S6A@X;^mF:M5;=C1jR_<B`Ao3UX1`ENZ@PcPEma2eHIR:GB?Nhg9Xl4b?JI
di62NdX19ae9QO2HPX7Q1GUh37b?oRE3>nLVZG@RTp2QVfDaMHlWP<oX^Ji<Fo6n
CRF6H8BS[gdYnPGGJ1U<PimY1c0[G1^aY\`G6`g]4V2m6@C;b<?RDkA[QB5a_`pC
YRF=ZM3LfW]6FGjE:g04:J?Y:dnQ:Aj:U0WF6CA]Bj:_HS_]oh[R\:<XZBc:=3S]
0<BSV3_;R\AlPf_g:_iL6obR::;6L13=4DRIMCm]7gZPlcT2XLP3W>:]TZgN3W7G
?9NGKlPU0;p3O3_HBoiWh6fIlH;\75e87k4RbIJ=46iW4[M1FT8;;[03>7n70XI`
;8@RHELW_l2obNXSgMamEgEdBYQb_n4Tf^1Yb@SHo>TEK91hl8V=DQHQdo^=Xi2\
\H2=?HOdK4RK>JOgS@aN_2p^@[]bPS;=9A4;FMBfaZ02hB15n\3\A4XOE0BZS9Gn
>@9ENFVN_2:1_2[WAFjGjjMWP9XTDRheB?XXk1JaaP6EJZh0nWC4C:W?kY8DKb2A
YKAn1i]UX5eZ<S[267adoQDWDclISnbaijpNAaooYn^8WOOH?bS>URXSMMNXk`]I
LY[iPDOR6mCV0kN\dEI]3PdV3H920]BmfGgciDD8hV@;7QA=4cbeWb^Jo70lk\:;
VlagNMS<Mg[TY\?2PFQ?W?FJ4kScFjl]PF^T_7o^?c7Ojeq0[61oe;AolTPleoZ?
oOm2GG]Eh7No6eN@Pgl2UVM1;<kZcU9U2_7D4RTI\PD4ITflJmLKOQFMT_9VH@OQ
m5bcRk\n=b:=QpEcc`M?ilN4I9?G0cW=ddNLLD]X_GP6LIT69A0GSekZ5HFK5UXU
cEo5O5q7]TiinpPQ]9jS^$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MULPAP(P, S, M, Z, M0, M1);
   output P;
   input S, M, Z, M1, M0;

//Function Block
`protected
T]c>2SQd5DT^<5=bg6[o>@;[cXh[C<TdD9Fn];<0<BDCoK>J<UMRE:aB3cmHa<EH
^aFI7AplQg5C7_Ol;[8n1IEMiGZDAU9ecnTfXiJ<0bIbH^X7\>JQbFUoApeHB16J
3@nU?5FehpMXdXEnpYnC\h4qWCYbSk<k2iI`j6moOfNZGb_e>mpG^WFiOL]b>kFD
^mUPLIdeU?0dQpPV`m:bohf:l1R5:Li2ig`3UI:bk:3<Y`CF20UO4FX9a\?M3^o<
eUAjpm_dVR<Xm^8eRcMl>RU][FQ=dZgq=7`0__;j2?38W`cHV@B>8E5:FXnnp0MJ
2K9dOLnViU\^07PHT4WV^V[Unp@L\hQOTbPJa[?JAXRAM9cl2m6IF8iC@oG]apEC
3U2I7BGS@X\T8\Xe8BIV;QH0V[`8S`O^_Sqj5cG<CUJ6H_ocHoQIY^WR`iOD>7JX
`g6O@8@<hqH>5jo@>9db_E7S>S>N=4CA`II>PiTDMn:=?4CDSo1Wj9PV8N5^0>nc
R>P7h1A4`pV3I6Qe=AWEX1@nBNO`KPnN_:bnc4]?8QFgOp:KD^\6VXaU5FHJ?]a6
b7@e_][j4E75bib3=q;R[h^UN]KI1:1cij5TRocdG_PlXON>?8ieUnpnR>[cJ9Z_
hPIa^Zndo1HbIY0F@N6YMh2@]UQFXpPTT_D=nlC32N4IkNB`L:m2ZiRK>7<bQRA0
K2q?<?g5BfPF5\:4]Q>08CWH>WU=4dSe>;BhWGqd312TZOq8O@B^Wp[N9V:8=h6d
cf`A4FUFDfJCPhP=JWONQoC723@59hA?I10QHTfbjI6IE;4>DPS]hHSI0MnjV\?f
5^A2=@2imRPIS7m9e1T945CXTYXVIPOg0Wa<e3G9<K<Rh3Ff>;^X?`6D8NYjQL=6
hLJ2<`XR=dEIYHMnpZf^;hC\\K>lZ1F9AWhJi6Ijgfib[^\hoHZSSNZcT41q6a_g
IiFk]9686:55femP<EENFcTJ;5_I=SAGOTUFMYeB2L7XOE=kgD>L\f`1`[XFfnCM
C?MWE_20knLA^fKdAH9lHX^d4Ma:=V<hXZ^ahC`\fKP@\^NBJOS0kNYOk8V=@\BR
O?jM@57I0nnA@@Mb^HP_mlq>>_YS;2_68jZIh:aIjeiK[MULo];gWGf_=n8aQci\
?:3G9FT9cLnKH=Z[2;PHgcESBIKUbjo2jNnOkS5VkiI^1`CPDba]en`_V_@_jLV3
alKPj3dI5Se]bXUQo0\^bHU@TbY6bTaIi2[WkJ6Aj`;71Rf<CpkYdnhbGVk5Ia9k
R[?QS5ahB4P]nVfCN6bN6m<[lO>6O\hF;0T_N3Mlcfod12AUEVCIL0DnHm=g?U@k
k8b4>Wj4UefFP@H\dlbkgICNUe62OBN@Gj`FJi`aaWPb1Q`P6;Z2Q0Nnko:__LOk
6XHL0oG4:O:6q[d]]iHTXKDcNgZ`>Vk@jTU]Sli:LHdT5nB^ol^L6N]UN>dAI2O\
2EoBR93UI[1>;j9YmPb^7;`mmb6AA;6j6U;76Y21I[km>nPOoc2eQK2L=Mh6i:_V
kfg_7UOUR>ac30QGRCb9:`00J868_m:n\T;Ce0Tp`aiSj]:UNVGnPVAUH1kAk7oK
@jApTS<\Wm6^0HAi9VefPXcAGB^;Lm1T6_lJ354dTC9Te3@Z<1ANk2llnTkTQb6i
;@eEgJ@>:IkCjd:l\A_SNbDb7j5l5;4l?;2l3MGj92aV7_GVQbOQNKIe11HnAgSk
fk0WoNW1RIbYWL4o^AT\e2LI1j3SHlqJX4lJSWNW>B_Ol;6bVC0jgD]5fWW@^g]_
RZai48mLgc2_76XLe4Y`?97FmEUB9P<h:P^MZh=a@`eb<=ZX:oegeogSiTg3NKM_
GECYYlLU>JJ0LWiJlBT4aM<n00F<DO\e>@NgZH3:neIc<Jnoj1`Xe]h<Dpc;lViD
UDWY]`9Q?V\?6NEObC9@J8LHn`=ZU=>WX2B:Xg5Ea79A[IaHoocbTVTSDZ^5e`OT
DZ=92OIZl:k9<UTiJ5OA>?Uiln=cl2ES=TgOX^mo8j3ig9jQVgkZ0LNFi:dSUC2T
X1A`>:YZVH?Gdk9ial=Jq7l_OeLYZ5mHU1lpj:1oQ>5RnjM:;j2@b:DU[lcUJCD_
oJLKJMXEgefKh?l05dQ9nF0n];^P7\>8EGVM8Q_GRSc2AHHM=aYZNnAea<3\SZU^
pQBIGnamZU5BIS>FimSUgZ<cWE`[2m;bodIk2`3]d[U9DXj=RMV8hdko`0:VY[cQ
\R;Zg=8SBL7@\JV?[V2160EWI]6b4[M?GdRU?`fVjW<Xn0T^agY9hR8XCT<6JJn8
eb@QY>8_j>JX12VS60I>ASE1TX2p2B5I[d0YcC[a@QL@hCV1_65o=o<8hFCoX^DR
;GiW=g?TG0kINTh8Gk>80:o`iW]8jVlITd;A:BFiLI^caZad_]L`Edl\P:jMX[6B
X_nRmJckAlL8\M9i3MPLO[OOS`5:`?6Cbd5@A4V4?IgEgUH4j][iF6pAmgBE`iPd
kSa?dGo4G@[K7449ie8b?NAF3T<i^:l<Y;1CMMC;6PdT:Wm[>`FJW]:Lnb^WPV\=
B9YTWC>e`dYLn@F49@7m[=iF<nHeUmfUOBA`:ZonBYjbYceFGfRf1a9Jl=gCP`n[
^CTKW3BVYE^3n]deUpZe=9<?IE5>6<k3Ze?8nUY7]oJG]7@0iVYS\Ucg:XDHkM0N
\^Gba\Of7EboSffJRVkj9PR[TKIgOGVcnC`M5BARDO4eh8<cj\YX;UmB4a9CCHo:
@bEF^1_CU@U0mcFHYeNMe=T[H6MXP4=c6`dX1?MRn>lGp_e=AmjG]Z_KZeg4`32?
7=OKanlZjQeEO]U1HfV[n0V;E26M\QhLTIIebg7k9EoaF?V\XBb4>[D:i:H`P9AN
NBe2519i5M5I5]AB93i>8Q`29`naQL^OMQY_K97a3RUHDHLJDhbdJbIY8CHk>[QP
29en8Phpl^>Lh`9Q8\eG\MiS0\KaoSYDcQRe]T1@PKPW`N@14@cYpo<aNh0EWc?;
:0fW1k_L18?4dOflW5a7dRcXiliGGbj^T`o0WWk;HAdn0JXL@V7<ZQSSa8RdEHHa
a;55ILkCM<hJThm?J39FWRn:_Zo^E`j;LiHMdR1;C3MO>h79<BIkM<cU^@Rob8dP
JF5FWnmIXch_X^Qq^D6YPS7H@mX?;7i;2To09:Z@D3:_Xll\>666a>oIN:j\]JJ=
6[i:14JZVLeoh_6d?l89HEd>40m0lH`@9a4:4dQfP?7loUYb>hIUE?N:;YL3NlaJ
aQ]cY\Q2o@gNlW2em<d@<EP=M2S`GHS5Eg?]2dV7Z7qnC:7:ZVb8X[W=`UN;9aCU
d]:=ca^d@h2UQ6]=TiUD25:>i=[?8o1i1@J9aDFbdDc<=IeEPON]bY7?n]Go<GYH
MW=l3_VUF=VUAN\1oH[;SJNi80U1o]oL16LB8A2c6dXYe_0FPXaRodG_nRH^`kF0
MeI=DpZS`@I5_9d@Q:1CIB2JG=J@K`NFgAhNB^2dg0YQPYK0SI4E:mJgoW[FRoCY
d[I2Z;[=511Ko>FE7O04\CHB4eA44ek8B1pagXITNJIe\gb[f6HIlVkN1o?488L7
M:`<LO?96FAGodjn^i\kDE=c`ejcklaXlgJnBlW]fTc0onnQ][[0eVgdHNLg82lo
LKP[196dW<]NTd;TeWQREm?;jAQ^eM:W`]3dUFlYKQJkRTqhIOd]`27Wckck?T<B
AEBj0XB4Ne<nH]^ML?SJESSL67iBJK2HfZqIR\SaUj?\Y;bU<R2TcA;KR`lm912l
<SZ^?K`dm7Aah:?hYWJZXbmEPng<ge:SH:949jl>0SBDM2b4>\C3nZg9<1^T9[4n
gM^?lT@Z_Fb]i[<lA9c\nEe9aR8o0A<Cg`TBOXcP<ghh5?p7kj\jM5n`L9InJcZD
N1YL<1F6n@Xie>B7?7@]>R9]4SfU]]GGAjR6YS=e78MG7eFnk]:XW74jO;b:`_SN
NUWiP_Kln1?I=>jkiG7[KH4X3JCeTdkQS9f2>FE_@e`T;W3\7L]j:Ia_f<qZIo<G
dnG4h\@ml?TSFk9AXST\o0NNA:n7aJ5YGhHo`Qg<o`N>UYjVhkbikF7BB9SV`ZC1
SG1PA\Ao7a;;QQ`MoJ9joAKCP7Vf:YJl\KX]4<\1@180Y3LLVcS5[dEd^88iEbL_
@=9NP8pkeAg1V>[QO1Td`\YeOo262TgjGfC\J:ATFE427AMLJMdI>4W_Y[JfMm_@
Xi3=SKLQOQSMV4`TNC5EO\F\diJH45jbHona1qEH<Re\SCQ4>9hfNTPXjJ]A@^JL
ejD5C@<haNNB_SO^@nV7432l]?aC[e4NeLYW`7EB[\AFG8n?i2PJYL7:5:I9_jnS
o]PJC6Ig?OZ?U0k9m4bUL3TJ\52o@73JT[cW03YKSMhF:o>3kW5JlSooq@MM6CQ\
B`GTC5I5\KaJh;C=ch>RKY5=:69ToXY97M?^Y:7kJBX=i<if_T>07EDWZ4BmgBaK
CqHKS>PmEi9109fgJ;\=:F4ca`PRG01\m=@@flhV9>IRABfG34\5^`6<\MRj\W[A
[8JE_W@555iUUYOJ31j7P8oM_WhHX40>]K\8fD<jSb@AT?L`gG^4_hROH[Pk6\Ph
Lg\EHVHOCoFUA:GD\<l7[8A8q0o3\L\_^5=aAk;QeA4QLlQ]S:@:7lD7<hT_^fDZ
4;>;j=`UNL9abU9K^liV1FQ8jS[YY1kS2L^KAiV]kn^H4oQP[T@N?JaNRnV_7:H:
m]Rd]oN[0o\ke\SZC<Gj6Y]=ML[<:NgHHB^EnQL0En^ZHaKqVU8Ve8WOhia]3@LT
hFUeWjWb2iX6fFb>9TXUX5oIV_lS^XPPjBlbaZ2>TD\`_km]V1\fi?cHPCd:^>QS
8QJnhkR4U14R1Fb<B0iR`5`ZfI?J59=jARoJRFHAc[Mghk0d6i3IF?;\g1MYQ>=9
M=qcEEZmaa<kXfDBko;OkZMN45GRaHj>W7ZZ4UX9afT2;J\PP5A`EB;SJV9STh]3
31fcM<76conC7iF8_MnAk9HpVOEchE`oB5f3gl[c8Q]S4hZlHk6MMU\SW=bl5e92
aM406>7]f>U8X@ULJ8_N`j_CNSO3j3FTS^Bc4Sh?HVibcJ;5?k>P7TU]WRUO;SIF
FX;a7kK=J8[^`Q^TLKN]KIY`V\m3>dYK`C0q]ZlEUC\3=`K\`nE_[BMdY]3AW\cl
blOL4C^K9ii2]Y_7K17YFI<FY=j73<B@WQDR2?PAGHAcgkb<kAL9:DH]6K[Ba\cM
^c6\EMfOcAb`16Q\H<LSa]mWhf_WjUAbQ[RaManG7G24Xa\p]>5\V\STaB8G5>NB
9Takc[Q:cGMn7eohVkM?UB@53W;lenZGdNdW`<VdACm:h48mPka[G@ZQMcSBWn3I
^3fn[:4gGGf_6MnNL@^TM2W]54oJ_PbGgKK\Fh@K^=?b56<oL4YPJ3P?7JZqQY@m
;UjPY075NBXW4N4QPX?37@MMngiUEGEhF]@XTJ6A7d\AncYWT`9@3bgKD1?Y06`q
M_6<CSHaTiU^OlWRLhT^8njGiXm4dJ?l5;X<>0X_^UE26fnIY<^;8HSnOKW_;T6a
c9b6GjJSRgPY\j[X7W6B_>YFQXm45jU`AAV;ccX?6Rc\;STdlAI^9@Uih>hoFMfP
K=l8[ohTF9hqiOn]ibVI_^fG5mm]3C`GJWAi0IXAhEd:Q87lQ0]WR8U3S_fT^lbi
j7=TPFIeP0?mCBB5eHTm@BhPKaR<lo^R<m6oH>J<f^qjjcg;ep__3k2k9$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MULPAT(P, S, M, Z, M0, M1);
   output P;
   input S, M, Z, M1, M0;

//Function Block
`protected
NR7=ESQd5DT^<`NiL^OdY^CDq@nNoTjaRj:oZ1Y5R<>ff9OP:F5`ZL?3a3HI^mB>
8OLD1oCDh2KpBBKXZ3>dMA:=?h2jiednp3E2XdkpEoUR5QpQUQ=3ORU9[UQ23]UE
U^WiT?8]6qf79?S]H2KHBkOFI`4LRTAAF?UMqgQOj^W<kE?O?NmVfUj[mBH9Ja^q
V8HU6Kg3aNMJ]aBfV:<i_3Ll>o92phZF4h3M?IgMc52Rc7iZLMK7pgi`a3EKKi13
^T_f`1FYBV6ibeOPapFa9C8XcKF9abh2c=YOWc;QdbHm1JedHd?\hqa<j<CWm\m>
SZPaA4L=5PMVNTJPMj2=WP=m\;qcbUh>=DclUdkJTUO4QAqI3953akPcYbS[OoaQ
c0TU\_Qml1IjPD5YOH9@Dq?PNFc<f5@??PFY?bRVk=j^7kVaYkC?ll2`;pQhOi<?
1jnOfEUJUg7fDVCV7AoNXHKANe7C[pWWE<LJC5cAPh5g==NZW[7e^_mQNWg4;f8<
6bqn1KkX4[igEle6;Xk<jXH?QmP_J1iA8B6G^WGjDq>E?:]8WB;k0a:N?B;\\]:^
]i;9MlWc48h8cWpb\DgieD6J=NTjgkj=8:`Mi=eU8?W@X;WCE?q^OdZjfeq=>`jJ
\L<?NBRQo@09gKnE81COkd:liVOARJe\CR9qaQofACq?>JYMcbj916]TGN9Gmn`5
90g5K\XT>Y4>@mg?mLiBV6mLUBAb3n`647I:aec]Ggo^m;Mn1G>k@_7Ln>5GngP\
]4ebh^hB2`EPiQPn_c9nB_f7H;E@YZ[A5N]?6JJa]m4E@[271^jRHiDjnWR3PUkS
]<SFRpT?ZZUR2:DLP<n1OiQh?F^2g[MUfQYCQ1ndnk]9U4@\156b=_;J^nCjB?EO
UBaWmeH[LZRVhYUU778:YX:Pm7RPV=DE?l?KUiec_j59?C>:k?>MKl6<BjT><OI1
]J__bTD:M?AViK<R;J]:GX69e5JPYW=Xq_a`TN@S<hkVFiiL>V?lK@CcKW9a\072
FbmjZ]F4204O2Ym_Ug0X7ond6L2FdGokF29?2SS41R__lZdEU\?@4We6OJNeXbQ`
1bNDSYC_Hee^<D>gTEUJPDc2Cn9jJ3OI\gK[jVSNm>9PJcdO2c61XeeT7mTpT;2i
TWAC09D]<5GU5A9Q2lOKl]8L@Ea:Vf\OoH^D^BTi4Io^\:QdJDWL=6kT\UPgFYg7
d[A8E_L^S;jo^3K1oSJ;8SS06PJDTHhU^NeZ>HFNgRRnB^\Z6abd^44HP?QfYm9P
8[=89?lfY;]f=;nS:SI361qMBnZ^`g3iV1M`RNU]VUUYG1mHRU[ZSg5B<GheQBI^
83;bI4<BXZ\9ciVhQGPgUQB:;gGOL0732F8`X``A>V<_bY1Wf?J1b0jgH]Aaj0MS
jHC`M_bHI1I:ZL:1N4k1?m8TNRDBLGLgNoOjXQTUnmBPbTI\1p:_fK_Eg9hefX2j
9aBWf?;J4jKQ8e?\CV>im9ZK]Sn7fL?[iBU6FTYi=njNTXKK8DQ3icG`e@oeg]c3
lj2F<mlZJMK=2YDbG<_G?gS9M=]jlX_MJMb@]>=E3ADZF>2^g>fgY:H`S<Mj7<O3
neLnHB@ZQoSbq4FTOcgbbjd[g>NDcNX\nLPLO89\AVN=?Kf33GINB[=XF]R`:ElP
OJk7P675VDQ06>nS5?44EBJ7h^o5]JgSnT4XAZA[_83MHW[cR`g^adhJn8hij@[L
>dUM0Jc?[cTkC?]0HQ4W6iFaDUo95khd4J4=N=Yq?c2Z2=V`hg\RH;H>kF5>I_T;
W;gcGh8@cj]_:TREWFk=`FORaVMQN3gF6H5=?3DXc@[WjWGH_Yb[dBX;;1j\mQV\
@n[UAeABa8UEFR9J5<H0=97J]lVL4<WGE]G4>?JSRH<ORWdkWgPF3Bf@i2EG9Q=`
18poI60c_BAMNA9[EgZfB6d?Rf4gjRn[B<[i\a7NW]LpkY]8HV1K69k9201iG^Tl
EUW?D7T]k@bPdgFgKPhFQ6S7N^QX1SLJ2ZlGHHAo0WZi7NU8do@KUO`EN95H;iY=
bN]H9I1_p6?1EI9_bbXHhoO105PQ0]fK8ZL_W4T45aI60gUX^IOFdePH[RD5IeeW
B6cGD_oW2kVjFDc54I8e`D5XCK_okZ^B1mTnJfRkgaR2<mm=YR]7R1Lk`NL9MFZ[
fWELYS@OU1jE:]cSO>NOJI5]oAPWiD^o1f?pOh2>Of9`S9:1=GN`do0N4;nN4kXo
1Vd\N?G0AVfAI5;Nc0<aRXlW5FH?09fT;3DU9ZokWgMVRIM4WL^>;9DnjnLlQY?6
9[SXYO8TVEEOcDMFDPNe2:G=MQ0>_DV]XdN207Z`Jg\in:b9[L@jAXlgbnRl;0qe
j8aKkRfMM8\XA;9?dFFgLM>B2<X`D4YHY=[;\4_8D1YEY_nhW_eoH:VYLjEjT;U^
:Xi:ND9<Q_^@idW1F]AnX;WNe[fILPedKY[RPLVm18d`];UBK3>nJ_5b6;bQm4lV
7c0:NTQ[DOgWi=aWjK^@X]YbQpb`[j<j_Ino=PiZFmCjlDXVM>LmP6R<F1o0j`kS
ERCj?KH]@cVMT4=]fhjQY]Zden\;?[f:UV?RWGIPHg]2CS\:e<90\YI_S<b[IUCn
8Vc5^1UOmRo0\n?VYfP>aoNR86WKH?G:34YKfQlPT[a=bbH:JL=Bq[8LfY43XGcJ
b2M1kXea490cYojUciJN3C^=I>`NF`Q15TGFkH8G=AP0\c1FZLMJJTAZ\^dSNP2k
21^K9iKC@<LU89_PV4375>Uf@_IInn1:QG<N=TQPZlW=5Xg8d:f0;2VK]\dOoDVj
l4^faPKG5LL126AqCcCU8>i[P]iDO@3IgMXdi;U?[f9Z@WC5H07>UD08FK0:CkPO
T:9jMMh0V=0gd>3Z1C[;U37c3]\5\Df0T9i<HfRTlbK7BSU=_?0W:B@GDPm3:YFO
`QneTn=>A[Q>MXR@:NKdn3[aKU52CDb0Q0>Qef<CfWqZ[_:mUT2UiV<NQk^0@NH<
VA2WQi;J0JYnYp=b<:leeNZC2H:W^:`=^?c;fRJnTc?jEB5;3oHZ0FXh\\C=AG\o
ZKD58Jk^C5:hl_T\SOVgMRDi>F:km=;X;IfPNmQUE_mLoT`Ni=<Cl7nD\N?jdRD9
GABn2P^Pd2ZWJd`NOB?go?<hL_@k>7@]NHkPeOBMpbE1T:1RXWZ:`Z6I7=XI8n5X
XbL@M1UnA9;>fYfMQ0[FcC1nDAh>9Ua[\CgQ\;GHLXFnHT@?8A[PPGE<X^^8fTT@
aOUdPW^lGQN113joUe1anD]MgVLGjb9aGjSajgEEe9Qgg6@V1;l3[>E;m>X2\]T;
6Kmq\gE<m@i4i];D[BlBhY?[g\7caY[Eb`JB5hedRN[g?m<400EN8_:j_bXMSG5X
;R3hR6`6Y9FJGanfiBhP0k\>DG:WdIUjp>F1M=\9lcVUJ[jA_[OKbO?TL>09GG_k
fa2eb_3DkN^IkV=efTaWK=ISUfBA79920nJX3C`fDJdnD:;C9lhQF`RHDE0?i1>M
[8@BU3SemAW^aS@5[><ZW@?@bYbLf=6V3Aldm[bJocU1pm:;USP3VVU3FC1Y\n`e
TTQWok5AW>`kSi6TAJIlJ4C4`S<\@RS[l[_i5i;H?\_`?ndi6mhS4_`H^e_<7h>n
A\b\E55bB\1k2@14K[i5?^ONG>9\FPdAg2fLe?[QW@MCoYeljO?\<LK5p`8LoXSo
5[=TSRWC5@VWKjmY59OT:ThlMYJi1ElYAY`d?OW?AKm`Pa1Q`BIn@PYMMA=Anj5[
:3kJ3<S]=^:b7fnEJIObIjY2dZ2h3mH<nCKPEBZUeObQdgo1U>ULmOTeM>4l6<ih
5S^7qBQjYk>J_9FIS1[3mI2GA6CD4O<9FFbN]WMccZ[4kjGGehgeIOBn>8c>^ge`
mW]FR@i\L9_;43CNlh<gHiVW02fY0<<ReA0G1ZdMb>bmF;oXbkIJJ];>F:8I>DM[
4H;hc_]fEhRKfIo`q=`YnZ?@mmhDC[Bnool4OACI5JAQThcnk0<jj<f5G?Z;O?fM
K9^c`l[O:V4U@SI?:R`_6\12kHQeTD=4M9<D3CXAlRm@IO1qI4gmVPieg:c[c1VB
l?V8lJGCI2PnN7c1Kg21aKin>eMFa:ek6k2aJJZS4\KE]]7Z3cVUaKm6>I:4TE@1
_9`@950ECdPkWB:YKcC4cdl`7BWgNZMa>9^^7X5RSm4l8\>JEMJOSK1b5=ofHEDc
Q=Q9A5mT8hpC73:N>fbQ[B5DcLUQ0mRjOLo2g6oL3L67Mk1>E:GVl^AfcWS1>pIW
F>AhFjIcA]m:G<L82>Ci[UI5XiK`=iSe][C>VcQd?fAi[mc]gV7EkngdNFc7gB\a
ig6=Dm5[Rh2_\Kd50aak3Ke[N9ZXe1S:^n1M78Pe5ISCM:?ndGVfQ2ME[llE>iQ0
?Oh=14aKn@@_B>JVdobkkQnBqVb<jKGo`cbkDIS7=9jXeXgBj1hKSOjZ4;ObT`:n
aok1EQ2jZ4?BoJS[UcZ`2VN4HhWeFJ>>QEol;o9nX71D=9kIGLI`mGZi\;c>G>[c
MYFQ`@lb751FkZ3dcN99]34h0J5lAi>EHJOn\j9HXM^Pf1kEG7Rpl7?a=Z`PaJNf
m\HaCPD?2CMclgI]j[hMIfWeNN7DY7V]0\C=[FhWFZF@;H=8o`GGUcg1@gUmDcKN
C6@N_o1ALP?83hRjmT[;IbBKkZ;dg5E=MNSmA4Q17^e9GT\2H>^_n_8KLgOh7JXK
S6>6hR8GLPgoY4p0^Li7g\jEJWOd0FVld@>B?\MKo^OPM\8RjjULX;^N3TgfAPG3
?I>8M<MZlB5o2VO@QmDR<SK]>VUE;Z=93K9cCl\A54_q<JY=8Zk@>bDccCEK:hKe
nRPLh17TXR8k8N?Q00XR^_ge<H[BPV<S5]9o87bXYHIP[28=VMmi20iR?QLc\RlI
\C=e[18J=??;SjPBn05nlIliZ@=H2KT29VA7`CXMAB?=6o;Ka29;Je:qRCLnRc=[
b`P<fea?5]ob8K]ST4QVK8XHho77>E\41<YKm13??=3XaL@3ROSUT@ThFf\I`7R;
S7?Qh1\gAX@Q0gQg;4=7CbF1XW\Xml]=kf^jnFM>AR4TP\KD`D\@XLlRiiZ3m369
nHjpg2Qf:_c4;K`I0iRLnT;^mYC\KlNJCCRQoVoZ@XjmZD6Xonn=WKaL7?XepJ]F
FH1;G5n7d48mfPaGZ5Xd_A^F\KFd05?4e?BG73`0QmMZ@lgI\T?Wg0WjGFA`OZoJ
9n3N3Xgd?m58MED2B85GGJ^b:o:8<d000NOh5go\ahLnPkc6=b@>PTNJc:^GJRbS
oEh[eA[Up;odO<;jT@o_Zl72B^MR<Cl?@kbXP>e\74PT9801YVM?i8g6k`=;jB]j
Hh\oCE6EeU92b8J\SFd9446VdHX2moSBPRbI:oF3>N94`9_C>anQj[>1SQCX7;Tg
8CM@8dSb?AQb8SNnAbW:qP:T4XmNEReGWVV?lSQnH7\NFeHk8klX?EPJW4:;2e[o
3aG=lf>]6MkE@V`^DKnLF0=]hT_bSn\TA8MVKRkiIF7ELD>?HT=pP?GE\:p]=G56
m9$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX2(O, S, A, B);
   input A, B, S;
   output O;

//Function Block
`protected
>RjjcSQH5DT^<@H1R_PG7kE>kWP?DVj@3Fn]SPpaCh87He`2Jl_mYY<2XQP=D@;c
al?<;GU]k]fGbIOc7?mMf;BCKZ=Il6>19oVqJlQ:Ne0gFfhIAb7SahRAQFb1C6k7
[EKn=KEj]\]Tmc=<Vg9S@9MmgFQhQ@@<M5\`pCl<X``pNAaoL6c3?[TRF=VT^d^C
@S?^Cgm16Z]c@>i=Ufa;7Io[1CpK<bBD]Cq@<F:Ag`4:oS7?RX]A66jgJSMmoVXi
QJ@0<XCKj=0h03Ukl_qO;h`d^q6FWAUS<R3C1ggk^Mg=5CoUfl;R9T:\IGK:2`Jl
=FmK?i\f[?S]=^DQSXIKo_cUQc6\gP448LX5GD@Xn8Oe\NSP0Ah7A>d:IN;ampIO
HWJgo<?iTPE>_Kikk2oHTkZfMH2K@`5Xj^nj3e[AXMID@kcf1ihSKAU3927d8cIj
SMT3>jUEKAYH1MmPWB[@Lf]8]9JV@ADf:pjEB>6nMjoHBFC[Q:]OSTMoFcjKeh4g
I3:Q3^4TWe[cON7_K8^o5BkO:iSZGi^XBjjjbB:\<;FF[l55C[;ZH;pZ`GfPTF28
S:OWh69aPZABX\=^FCMd5nTYR86D;A9B6l=kBpUZmSen\?OLM<QOD6gf@2ljOH:0
K?l>;TP[<RLXLXNDfeaLij2;YV@8WeV4R[KoP5U\2:nC8L9:?eVB]MAcjSH0@Jm`
P]Q4>h;^3n7A@5J:_BXFhe1@q7KKD_Dl]6?koLfd4He2ok?AH<8^N1egS:VTYlPV
V?M4?7E7;<_g`EKXeRDcPUDPZ7IYjEnDSQl=R[lS=kdmoPH]KU_jl?]C<;4B226c
Eh9iKJmDTf1p\IAIU6O2O?O2?n7C^kP4;YAnnDLgMjU5\B2HjKOe8oAE]TlH?OnN
c3Xjjho6Rkfa\b8ZS=]mW0\7Zk2mbejdq[6B[6f_@K;HTkBh`X1eN5aS_nbl210>
?JXjG?O0=VXVR8POE]@]hX6HFgT\[Bb4>[DHR:H`P9=N8Be251li5M5I5T_Wd3V>
<mCXp`o4\O`SPQUAf@IK6IT3m`gKj6oW_gn;e;SQ@D3K91EU^VSnb4\0N\7i4Uf:
KH6fF`dBD5k0XVOXT407C5hWTie?k5a7Ko8;Xe[4p9U;k=oC5H4M\Fc=79>gH>MC
nOB:FGfGIa747E^KS7TjKL^eUi]3S\bC4Kb6\HNZ[9Xb_Vfmb;;R:TUQ;2RW8pab
7[RUq7SVBnVa?H9T`>Ui[_\>3`XRV`ma9@YY1WG04]8?T2_>G4TmC0T>pdX7h0i?
$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX2F(O, S, A, B);
   input A, B, S;
   output O;

//Function Block
`protected
K`=c0SQV5DT^<70M=e?D6^6iZVHjWcYNh@847h;KK1B7>YV;Ah4pfAgWDeLeNSRn
[3OafWUNe\732KLGMoQ<CbT]U4D4N6ZGjNS_Eme`l\Ti=IJ7A6pVL[=<ILWG=CkJ
E?nOX^c[<b:LSWKo97Pg2ol<NCLM4mT>5_j14PE>^O3=EjY;[3W@J9Le^4pnVL>g
HqFM3c>NYi7CJ7CSJhP9CPnB=ODR^;_L3j=f6K1C:RVC:;B4qK?eXY^hqM6`>]dp
D>T=W8d52F[_aai:]Z?8aB\lF[KP=29Pl:TZ1MbDcJIM:_>I;o78_=H3fSD1eahn
i=1M054B4e>fo;=>6]SEjcokn68]KFVbDK^Z`4bkK<mp=fDiU@LSEddDV5`d4DHb
XF1aO4AK?Vi]2_bVQMD7<2oCM2YPc`X8TJkOoW[4o3nR^kGSfdkO95=`SkmC<T?7
?OcoQOEoUdGR`@Z8IG]=gCIpZ9RRTAlVoWaGkQI[?1JVcjg:5`jRYLie2FT3B4_K
hPlh?4b]bjMo?YR1h_AT3fTB\IP_N364O^\O0<N4DUBdlRaLBTYlqXic2^DJJVg<
1P[LDfL]67YLEMFiT<g7b@5JF>IOd=ebg9ogMPBQIZnj6=_L?Tg@mRNIX4h?mWn9
KRAA@mEk1[CGb]8o0e3EJchJCNeV<=FFNRRJoX0nRdbVAQIq3^NA_O447R\4f:W?
4<YgW=JRh2HOnN;YUfd7:W8n\l]K2[h3^cP3@Ma8C3YES07hfK;EE;6`<\4\6E5i
RH0@ekcYA]?Njo:c=Wd]e419bf^H_^KA[\E69M?S]6p7eD>34kaWAL^TN@i2]>_D
MTcSBk1QV_3242l6G6SPY5^UH@n=gNHAn]n43qQd9:OYTmW1HE2F7FX^jWGVYTeM
K0A@YTJG1U7P><OFaVKbS>bbZfIUTN9C1Wi0o[<J7Hm?;kN?cogJ:Ym3imW^PR7=
2mqo1YVKa:K8a_egoJLb[?oYdYP740>N_C\FgBLZcR6h553\aW[baAP1oE6OgA^A
JmWJ04^3@THZb[h_HCHPH;g4>=mYF;nAIBA=AFihaD`Fm4pm@l0Qk@@=[eeiZi^Z
gi@2cNkf^I8MaE=Pf:CUoofh:4k@JXk?FAO_m7]1mYXj^[Qb[KMh1;nnW4bU_BlU
S<5Hl;OaZaXNAA9APCh55ggbCfpfD_DN;LbGY1\]87QH;HbN>LXbOQZVKKZI50X=
jJ?CAiE5Wl0I8>KZDQi;f362@OL]Q@4\H]]:hk_0f49PjG]=bP4:nh5pTVeO_UpY
km]P`g$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX2P(O, S, A, B);
   input A, B, S;
   output O;

//Function Block
`protected
Ok>aZSQ:5DT^<`A1QSnCn@jK6]bITaTU>gb9PGgQ`9QUZNhUQYFe\3n:RbMB7fFD
qMblVcU9N:_OZijSS:HPK2Jo0[=k4ahL\GH:=:0`1=V5eHlAo9AMlE0Qahi@qT[@
mdY64Wk4?:bOcH=FZbLg^D94]qOFLAgTpEN7XeNbj1;PC6oZE6]mmXK;[<:hCe=I
Of=o7V1Fgf[QJcYp^eFK8OUq`eRJRlq1F4`8D<R1nmahA2K\\ZId0FVF\@7l`chZ
o9M?MaCSIAhAi6=>7V3BJmP_\QkHMQL1RGQ268I0`1^R<G8V^92T9XfT]7nTKcRh
f>piOe5R2[<C6doJ_fd^Gg4L:RJU?@8Om]CQEB[QN_Hn>mP5cZO_NEk3M2^16Y]A
>D^i::3GTKTFFIcSHlEc9`j1;XROUD:2j]m8AWqlQ_9k:d=2LU<Y`>DojKY6PnU^
SJcjVOb`iPdD[0hB2LA]FDfLQU>@DaGRAeFfaNh6^MpA[=on5SG>HIa?8B0i=4kL
mgRnaYeWkSiaSMjB7AJ`Z@SO43Sgdf4NPARNlm5X2kSAULfOoZdb92?OlnljQ>0q
TR:]nZQ]>KWo3Dmk2=M6XHGVk?d]j]hecg[<j3O46hjK9H0Odo5df]G`d=a4^DXe
hX`_KG]Bg9>6BcH^PcAg3ZPa`deBRRh54PmDnYOMSl^^Ye8>DcDcFoqbAjQ4X?V:
RYS5^>bTf]7;6YcF_fJfoR8f88fX>HASE[:UgcfnWVgB1cmJBN;:3PSRi]K1>3SS
DPK3ZOC5LGWF6[T=9D08d1cinmISkJ<;HfMfedjoNNJHJpQGOo8FOT]_WY9nX><M
N`^[D^K1``k_M@jF=hf72_a^lHhUHl:MGbQ?Se=`:MeIP4W\<X]VeDM@C`0V3LRG
CY]OobqP^86Ub8;DdffeUcMa^^58hhclNRdVn\`GR0bY9^=9>\[mT94TAZgbB4i1
>H=JHmWIbP3bUlon\NWHgBc\FCC]]iE^3]JYHVXYH0Z;:lqYN7J<iZ[T317AYEj^
W0FCS__nELd`R_VSND:OWgJ;gc`bmRUD][XWa1MWJ@kTWCUBYW6W\bFG;I\XQJUJ
gan_SQ_=>58>m[XU]DE6egqK^]GH0FPZSVnAJbgbm14UEPNbHPddcNH`a>DQFj8B
?alHX8gIk11OEC]H8G28@O5a>5DRQAmm@A^JhCX\Z3HWgLEpL6Abk2qN<@5k5^o\
;1KB@HRWD3\b1Mg^maGW>>]9dbdNem0E1XENT:h0F34jSpKI2D7KN$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX2S(O, S, A, B);
   input A, B, S;
   output O;

//Function Block
`protected
V2L^3SQV5DT^<45RlSYR9Bd\W5J2XdBeX?\Q=K7E2Lao4J@]o;enbnj`0dEDh6@U
IF[RgeFCB;\k@FWqf0@QDGG;5eH3_>BbOc2KaB3b2cib<iMqCjCLd8GI2aS@h\e8
nXcV;YeTSS<:<6bd?ofU>>PqKW>Qh`pA\k^Dgb:j;7A=m6;;iQ<VCB>EB?3AgcBf
6\PEBDbfajD:lq23:oNiiqf3IjdlqEb?E8[L3InXH@=[^fL4Q``Hfhhd49Ok4Q55
_Cg?:iefH?=:05XQJ=mZG\@iQm2K`EF]5e]IiD9nOXkd8f?2YX:^DK]j7`6k95I[
peDOgeYePdQS<@c>XY;FW?kSF<5>VbA:p60D@M=Z@CoN2CWKiPDDk@K\h6MEF05X
:amG>]QM5h@3FAU[TYAUh@_]hUUT:M6jl66JRkNfCedW5_ZiWKc]m>aa8M^[Ck7X
H3VCpZ\j=N?fW4KPe^mmM<1Q;kPn[DBoZiRP7aNdL__VSjCXG9Tom;ej8:g_]eTi
:Whc=ZF[lh29cHDOCcKk58fIIq<6S8^QNcPWCOMIeK\iQKl4?dBQmh8HcX;=4MnR
Wlbk10Pj2mK<bkEC0N3=VJaY15<cfnaGX_a]2UdX<fff@TED7m3=KV;T@4gcIma`
SOXVK7<N:]b>p0:NB\CQMN;J@HSNbffFR2Y2SNK:akPH1SdKDJCm7RheQ1<@=Ll@
eC`VW26AN`J`D0<G3N>i4eOY1P>44>F3n[j[ak5^T\COO:]9=J??gNbaYm1mn_eq
]gZhM:We`QI55oE^2dIQE=QVKfGm:]mMne9dBH_CjQY]99e^6VaB<jDInhTeVP>B
]h]kM:l\HJfiH[;1Qd_nq_1nU1gfFFCb76G=GQIO<NjRMe`El\13A6aSLN^hg0YM
=O^<2j89_8g39lHfYU`V:_0FT;0[i[<7H`[WHl3oW3gcJC>T1nG3_`ejpNT?l6UT
=1Zf=4\:3H0Bl0E]7MDKc<[SNdKMnBeGaDEO4W_aha^k>Y\_?Ph>0O3?mNf`\GHj
NYi[\Vd2D\3`F^nde?DM647Sm7jIp\FMH]lWMD`o\NkP;d4KVW36>7da6lUVKQA\
?6_^k9oR3HY44??WT>m]<U6VfQ9]N6<4q>MSZ5I]Cck?7cmJTcQd@h@3F5?[N7Af
X_Lo:F:OI;;90Oh6TB2>C_oDOX1j^f@ic>^B3\W08k`HUZ4Yn>cL?pD7bnk2q3Jl
YV7Z$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX2T(O, S, A, B);
   input A, B, S;
   output O;

//Function Block
`protected
jQH8LSQ:5DT^<<FhNX[g^^MT>UlQR\=gq7TO`^[UE@n6H1F:761[FD`S=4\jQAJY
?1a>`8mTB`Y:Z[bIFSeJ?4aUK2=nf:F^p_O=d=e9=3cXMDoESqTf3Pg2plJ3cB04
a_P=6`CZ2:k=T\ZV:o8ZO]gQF@bEafJJo^A>dJ0pERPVFi0pZ[=eB`q8:H]hY8?]
KgL2ioGACUECKkcN80hV0MHX^aK;3kGT`aaej;8eh8WV0I@YDOhcgGR84YI`e``C
>mfDEFkA[1;62<m1K\ib0M;aWhqDdZ3l]MBn?fAi?mkKQ5eC?;j7OiJVQkn:1AO?
E97g`>mgb7\<EMPnM@jR<06fbmcDe<`A8cn\_oalMKQXICaYYjOke7b8MkbFn2qG
QBE=B@8ESDCfBoA;XaB8Fg=jO8VQCS6>c6mWVO@1cMT<NHgfPUC5=NNGV1YEIUDG
GKk72gLLM;kRDC_4AbEp3B]\\R>Hg`=U?iea@MeN=?838_:2T>5K^9LZ_aY1m`in
6>`U>`JfRQaj?KMmde@6RW9:8CciP?gSW?G5_KAMnjAln4j3B=5WL2O;GLP_k9c[
4K8KeQ`c6=pI?<JBZDiJ9@MiM8<5HE>mh7W<`gnefS6FW71JdoT[dYRAhmXClGcO
1[;n[SA_?7;q=^TfR4M\QcnKo;c5N`Zo7CF?[;NZVi_@4gLh16Q9Q>KS\Q=LC:B[
ZcIdA\8HC;^8L;[BkG4Hfe^_X7mm3ncIjC1en2FL^>?gVHUX9fBHBAaCPMV8`Wl\
kAp8\`AcaWe^]Qk71WBb80D\5cV=m0ac@;nec;YYg]?SSJ?Jo^4Yo@da[Lmk<oG8
;?RYC=P2A@?`n7j2@PJEe8_nY>Np`MAH8EJoELBaZ`YBaNbjo3;3=f8SFU\9<UeS
MW<O>nfR>o`7B6D:U3[5@EIM4fN9KY`7?3G4:J_ZVIf9G=<HG@U\fEgd9;2[8YeH
]Xjq8lE;Xk7>=ER7RfgR2Z4;Wa?_ShI`8aOQ2NF<UXA[ClgnO5X9j5K^j;F`U>`e
C]R5_U1X5<[o32MCY?nOaTI3;a?HL>BhX:m@G`Fo@6Np[l?\3e_nA5NA@CkG5bbc
U3VU6UA\LhR\CI;Xi:TFpA\k^?D>Oh\bZnPG]0`55D2bH5X\[io>22=ATUT9EcFC
ShNXV<`]0h2BJP@:7T_ejT4J\kllaZ1^Q=9:T2i8QUEFoqJlE3?7p]SgmlD9$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX3(O, S0, S1, A, B, C);
   reg flag; // Notifier flag
   input A, B, C, S0, S1;
   output O;

//Function Block
`protected
\8HFfSQ:5DT^<X=hMdajEPb`H5?IOoaiB0=2\C\FTSZl]IpfPVhIEgVCHJ^KgnO=
;FjjQq2NJNl9K@dioe^>?52V;Opao]mZ=q3:dBShPiYmM9JMTeJFg_5;7U2S[hhi
MlHh8[L=n=^k>5d7<LdEhb@JTViKGp;m_IFL>pc^^THmq\j<f<7YC>gQQ??k[miO
Y:giHhb26faGIFI1L=]hGRAm1RdM@[YS9JIeGX`33<?gdSA67I8BUU4AaWi`;lGj
kL[\a^n<^GN8c@<1Qa<P_i8SdPc5a3iVXn::Vc1qU]TIoKEgK=kLhRM\2WiADQfM
`SfUaO_lFldF_BUgM3k<7g5_Eba_oDle@GoV[jO^Q88=RFd0?D0m2^2L=LEEn1R<
`Xol6cIUENd[TaVFShPW0Se=6W3@2hI]WCqPk<^EFVml3leP^aNodH9R;9cFifNh
m944l4HNj<MOAKoRL7XG@U0i9=8iGlL1A\cdD_IRb:[XElhOkoj;ZY^>VI7G5^o2
o4Y3[40ico@L^Y81:[8a^Xc\\5YXDpX^RhHXS41jj9BKcnmlKjNY]]?Tm]fdA:RJ
GWl8RWlE`:P`fPBT6kCJ^<4eJJYB5lVP7`EH?_TKjSJgS^19AM8haZ\\W>0Q[dUh
GiXIJkF:XPoFLQR<go25O46SqY:QXnCd:;TL<F2;YnSZlFVaPd>PK1b1D[=25c8A
Hkb0R0=HkffZNf_`5`:Ai8PE0G`<U?NTKB9VNKM80l5a2HlkkV]N]qg2@\PgW3Mg
DTIWcoGNf3g8nNQE]\g;:\33_cZH6_U`?h6DNIcYH\3:UNMjGZ\QaQV\U4qcWheB
6aBI9kF_C5iB`1nY;H\S_M92Z_BXUe5a?<N6^88]>i44kPjX]=cSVPdGNTecShZX
f]\Kd[gT4P>DN2ikgK]^M=^C>_40@IJO6X[<VXEkUBWF3FEFIG<l\j0lR7\9`RlP
NJNWYoAN=OVh0pMD_I<5aU6iIEnR]=YPSTX913:2ac[1=hT\iO=\5;P<c16O<4^h
ege70]hia]^>4SMdlI9kUIiFW6\abEhT=l[oXL2M?c59=jAEo\RFHAJ[M5hk0dei
3?F?33gW^_H@LYT>nlh>>41ODb6>EmOIq=f5X3Jkdm\9dMKWmJX6D8aUGZ^[[KkK
IJF7h\amWmZljX?D@3g@kPN0ZMk_Y2J<Y=oi2G8Q@h=V096WGI2W9nfJ`<ZBd6eK
LTEgiV=0a3DBPBJST1^h17ml3@@Ukh87QT91CPD^X>U1ASa5Cf\qZ1PeVL4Oe;_=
D:GpR?nBeR6IV`3@0<52fIfbab6DEGVKf3jDFYEkSYFXU@[NMW1CBLUIY^Cf9L:f
GGgDR<mkV9>76hTTDB9iGk^NBXH:WhEXAjjS_5^B8ZSCG0RE3L1@<B0oJGQi_[kA
\0To1@6OZ4UTVeKG9]g8OYp[dQ_fN]DJCQadC2^;_TSIFF;hUkmbB7^e2g4DMCPI
2>A886Z@ABU]c=ih4b2Y7H7[jNALRZUmeOIT@Of?^6=COQ_L<R0i17WaY:gDo6^_
CKVEC@IL[i8Hfa_>5mRXcMl4OBdmA<GbNZ\FHJ3;Yq_ZAB>6ZO4cZJR01h7YlgjJ
=gi2c0]^9ACE<M;mCX3cHi^nl;D:IikkT<kg[8jWGH_Yo[dBX;;?JYl[hUh;=ceB
jCHjUhFR9J5MHa=97JdSNf]4<FkL5<eb5Ob:Rf[ThXXRVjMGf`i2EG9QZ`Inq>=G
S>^QS?^40:N6Y`DE2<7nC3R4W4Alb^N>BeCSXl65`f8I_Va7hEEol2k_J=VdU>?j
3\:6hKiWBm=bN^:7I^3:cg:neeUl::SB2mIm:PmF9nd3JCiPL:`0nLl9U>VIB:Mk
?dCbiPA_A?U10]<qTj[7j:K>cb0`JPB@Ef3>?^cdCYE_2bWX<Io87OkAM_d^<2;k
MofU6ZM^4F9Og70aTS[c^2\92Se4@2?oG9o=RL:n=c=EIiWVi4HGA:<iXF9U0F:b
KK2>C\Xamna^PU?bea_NblRKUF:Sa\cSQEqlY1OSK\PABV^`d5?q@6ZbKLlS7K3b
h1\11_5\a1K:Gkl>a`o9lU1[AkOMeO?Endgb1`1j@=5LK>\WGTI`@TT2@9TH4LRJ
Bkc_RbF4[7q0mhU:Qg^fB_Y2i0g1G>2V@LJPgbL76C19JC4DH?n8DAJc;Mg>hk1O
VBEn3g`4_oE[:=EdW=T7lkbU4]E6G`W2c?^7gj?ic1HUhQh`ISgC8ETUli2Q5_24
Xm^HVMKQ;;??hBhDWJhcBpkBf3]SThGk4hD8?:IY2^Oeb>TgL>T4GG=WGDI96m4M
BO1Dg2Ul4]J?gT9C<OD^?FLhjLO[_1M5N785QVJ?bm?oFM^Fe1SU4`7]G0RL@BOU
O43fZdgTW<>;HJF5ib?2D[JhlEG=p9>OYo8VcM?HW4W2@f:WJA6YF:>@JPAVC5Vb
O]e6je_i5Lc:X=L0OeM=mcaH]CU_>Rh[T9RgEVH\l9^VXF:LmXg_6\>kdK^6UIn5
C_NnocCa0m=[7C1W7GO?iTCFA\Q]6A[\?MRCEf8pXSD_VH82mFcR3T282WdGHmi>
NAk:YL`0dJb=OPBA9K3075]9VVV?kTF2C9C[3AEYGBk91VGF4;h<iNE7[N\`nSN:
[nSE;f9TiHbE@Qo4UEX4Ie5<@Ya5o25oPPB5UmHoOB1iACpI;=>Vd=`n8KQMn5K^
1BYPJDUBA7<5RQ<ZE5k_`eKd;I=:H];;Cl?8_E_dja3:dXMiOPc:_6>LN;M6Hd\R
93:0S@Q8Rqi32=O`AmT6<XG@DgkahC^0OV@[F=FiLSYJmPW:\Dh8aCNenH=Whl5E
?2`BfLoTbIilAAY_kb9g8Q36UWIifgEdTnUncFWF4oL\>;UamES`m?a2jlE\e0[b
=0fjU?IT_?QOpL2JXH5=OlDPXTH;hgV=9lRhOM1W[WUI2>CHF7h1O`Xmib\>]nO5
YFoOFmAY50;kbLah?:Pe2B6WDAZC0Q\AeACll0V3>CDbk3Oda@CoWmmTFndff<h;
=L9[DAi\2L;^X81pJ^EQjnfd0g:@T7bCAi>a[10Oq;TUeffTY^bOHA9PU4EZUado
9o5B2Z_]92;1Bm3FGC_:=[C:QGkW;hW@8b\M_WC3h;3L;S_R5HZ83F99dGJj`VZZ
N_>G?JKHhZiaU<PJSdbKIk?Nm`nlo=Jah@e[8:Cj?[5p\UcX;HFmhlT=@Vh6C?lc
QQ_L7`a5AFTcB4VXRP]Y?I_^eY__L:5?7;Xma3c03Cf^\5YZFgg7dYoeLZNF[jG4
BSk6\>X:>j[oR?b`EJ3?FB33hE969=lEEX2eRMI0kCSScNq4BeV>R7GPUgOlf_RM
@cn?EN8NG]@6RbnJG?l]]iGZng5Sl5i0kJ9=Q@0cVb8d8Ah4<AWjcIWNAC[LKRN5
EQRJX70\ng<[^_;H[d?a0BojOBRhj<6[6bZAFnTU@I?_8=_KNq@N^?AVYOlkaJYg
73bo4e9CS=S]C8FRUC>lET8j:FX9;>h]4nNIo>c3Llb3o50A9M@DS?TH`S`1;FIj
;XNHFZBHP[_W`l\e>73l7MlA7h8en@iVV><6PXfJ@4WNeomAUTaIqA1c9C]VZ4c`
_?P5?Je4Z:Zb:COLE;<iY0KQ^jcDj9b><\SWn:Q:Sic;m\EH:U^>1AUG[i?8hBjf
F5e5ZPI@D]@1mdGk4H]m9Q:Dn^_4K3A[Lkc>29;BSR59<PX@_5^>;\`q3M0[Q^C3
8X7=ljlKHN:e?:e\W:HS>TJSHPUbB77J?;MJL<1SQX:?XHCO3B_?d0`k3L;Z50b5
6OeV;_hIbYoGbL]K^X780mn4a4B2im>R`o8_XN7ERmD=b]\1e]l1e0Z<T^p^l30e
YK=I0O:hh:M`:T^k=U;0R5D?49FIKBk\>?HhHPnP\:W:^hjgQ:SSEmk=KXn^<o?>
l<4aL]V8^;_CJjVpec<P:HUAJXFFW5nOf5e8jFnk\?j3\QmfVoXfNhK_<QhP<P?h
22gamQacg=`L;OY3B<DHGS;[OVG^5WU60hFCM<HELE75FFmc`>XmgIZaVdm6BiaW
??ddl`SR62phHAF`4kRkl2dk>Cj^2OcQ9<JlhDNZYml=AoY6NV_[W;J]7D>lXEL9
81An<N5F2bY?>3eP<S9I`2@_ZSnU^^[9`I0<LT34:\P\?o4cQVTi60jU^Zo?eF68
;_RIapROd[3ihT2HifeeN=QMdMOen>XgKSfbR4FkF9@TlmLLYT`<:W0:4qaL]UB_
J0Mj:7CC8fO9N9RgbDFNNfg4508UcFX6<jChQM`]UgK@kEN[>C3[Zk66i6AO_UgN
h8d=ZHNTW^lV^d80f]jo`_GK_Q@2c`1PcG:W?\g5Z3J3dNjgGdb0pKR@5@Cb`M`4
6QRdQ6JPNHfR6G@UAPXTHG8T=`;A>2[70gSZ>@3:J]GAh6k]P>E966Oh6o:QW9WU
^<1SoK1_nW2bf;7EYL;[4M4T;Z4Lf<IY`n6h60]hV<Rm`V4q9i<DAT:kBe4n_aHN
3;Ci<VP\?98nN_Mo4`:i\IAH18A1aFI^eG3cc8cRn<CSFdNj`Qf52iI@:05;87eN
[gYDObMm12Hiqn@E1emq3YNdS\K$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX3P(O, S0, S1, A, B, C);
   reg flag; // Notifier flag
   input A, B, C, S0, S1;
   output O;

//Function Block
`protected
ijLc9SQ:5DT^<hbD0B@hTYDc`iD7O:50gbiZn>`0jE[afLi@>of5CZJ9h^mp\\\f
=lJ0\=1`<9Wc5_gCaR\`=0J]90:5I4_BcYA7^UXghXI?]d2BpF<RVJMSKbRiKW_A
=DR1eTgYbq11F:Fbp4iX15Zn1Ek_06e_3hF[QCQ\o_5AMn;0l6[ob4e5=\P:`hP3
N21=HV2Oa[m<q5^HYa]Yqe=:I?OqnZP344U?NC]:0YM=VK<M[joO^P3[:4;kSCAn
SnU2HKdScC4@D`4oKHnaNjRMC7E^A4`:KeV4YCnb;V?C@^dhjKna8m1UEACV4cAd
J7F8R06lZV3P35lJXWWDC9qe@]E`X?49a9@L]Z\0WngRKY[MKNTM7\O8@`BNX8H3
VQAB1X^TT7Xbg2L9\]n6?K4;36P3adCe54FJ2M7[0CPb3mHo9@Z7^Um1E`7=^oWS
M17ad04ZenQ6;WAEcq^OKQbLmM_\`i`eJJDo:OZXo<5?CO6WUkWW9BU7R:WlTpc<
XUbab3bHkiKo=C6`kgRc=3R>S6Z[`QZ8OhUUD9iIWA6kbCBFbEUcfO@Ja=BOIX7H
N6_GYHIC3?GXiJFX@i<gjLV^8iH9mF^9O>YE14k[eT1mCGPY<0:RdBG1q6U2X<^L
BX8?b;E8\aUioJiFmm<T5ih7T5djoG9ZAUT_:VdM;cBVn>91jCnIjK\15^D35:d4
:eUh4YlegP<5[iWn<T8C3cCGfM;jhVWN40JJBK\RiN=5MRPLcTaplh>h`Y7l2=2D
6:cl8BEmje]lDOM;kMO12B7>HdeP`Jn<<f>VTmnX[[81@_ZV[KA^YZ_S;P4<?R;_
5P^Y0aIDHPM\2<8[q;aSK`?lOe`2UYH^d28QAHEd9_[2jQK@M`[ZRiH06obEDOg[
2^E`X9`<17\B_egRBdXI0cfE>EW:Yg7Gh=@YMc6NO4O<=;6A\[[ZU^iX2Y]fd5am
5FmL\\3h\j`E<Y\0Z;QaP<lbhO\X\k;]3;^K0>cp^7R@[SDi<@OR6V`TV9LHQW\m
F5]EV`:_0V_Ge_nJaG[6n3=U^CAdo>fIh1h84Klm;LnO;_IFPH[UK6lQmQngEn]7
bA=^=:`]k3S4;cRmX]O9h?VKfo[Hn6FI8dO2]H@\^6PcjAFHZT@3Lj@e7l[D32q9
9^JoRZ<MFnGXeqE4;kH2>0gHQ@I=Z12b7]0be<dn7AO2_b;OPiGQn7`NFi[HiAS>
B[N_S1W0QfBTBX98c0D<hMJ7:4CH`6<jTm<NE2Cdi[f3j:1aPZ8aAef^PYJVK;fA
;9j\>6QoT3NiJOEQ`kJW>@I`mlG_3LUh4KQ<p^G:\W`S5kmCGF`4d^]FU02B?X^Z
6k10Iedmh?bf@DADo?gVH20lPgKQRlY;SJXeEbn=`m]oi1\9AZ3n;9EKjC2HI`1n
KG1`dloDREdeP?P_N8G23bg0mRjQ=H[ao8H2[^X2>Lh8<XVWD]h988APe22qfJ4<
4;CEo>S:eog=nQ1]W03\PkYHIO\DJanjY@D3b7R>ej6<Kl0FeX;XiL6A8SHX9]GU
k1hCVcmE]?5?]4`m4JmFLNmXjo=CQhn8JWgPQ4ko<2leM2FWc5UZ^;?53eOBfEOZ
`SgDImV`<Ij93oVQG?pWgSAV8NVEMa3ln6UP6lUin`39[6DAbk0WS;F1dLjci2gD
4^6lEJW1V?>?@;nBX\kQ?M:72AGIh1UjG^W1X8WaD[DS:HHifO:oE\O4^\jlVWEl
_ZcKObSl6[?oSKA=NnIWiBRmj4g]D@Z77XXG`\>b[pa5QK`6BaRQ6?E`akjg8L24
q0@bPejZM?]aMkc8Eg^oGb;mm6heeGB?[`JY<\d0]mCj6C9j@4nAIo?@7B]b2Z67
AOeLUDL\@=3O1_9]gYCN5jWPQ<cXbM3>cYNY0UUXm1\@Y<So=<JGe2INWK`D1j]e
B0m:9\jhKn81KFD76ne5]UIpT?ZZU2FOD8SUJo:lZ;T\17EH@V7FCNUl9X6=O<KC
@boK32A?kh^1HMgRloK5DW19K8CUXD8S><od=iG369e5nQ7o[;4T?>DK?5n[0@`S
Y@InkKK]M[KFE5<]GDWo2aaATk2ITVNZUa0_8k\6F]U^T]q9SN1mE<m\nmQaN41@
dKOeN9^AU1lIo2WcI24<e@nH7l`@TGJSd>l;m=_kWC0^7A1>F]88nK9812na5_dG
9967djN\Mq^:hD5<oJMO`Z[h<5KUWVY=n@4IeHOShc60f03GDB<Gaded`2\9S]iB
bP;B6RWJ`gk><PY246N408=X<b51c;Bg\fQI\5M94?F0J=BEhgH_`gj3b?mgLZUg
;W=ebPUU`DUWeTJ2N0O4pYFLGjDh3V0lVmA^>`iFF\1?Q_]Z<BY^><>L_@l=h`T^
AM0W7QUTNA^oZ9@BSldXL3DL1FE^TDa[T1\Na?PV;WhJX2]l@:g4?D[OJ@BB<8]n
ON5`c4WSl6JAWMA3`>X<>[U5VoEDDiCpnhLDU17SDJ1_i^O2Wo;nbER1O>o;onAd
Whm9Bk?b@cL9O5g1iL5Wc\;>j=o<UgmF\:UZO4:Qg7PLDPh2VOlVjf\d;>o;Kh?;
>8V7:kP6oSg8ckR8X\J2hcK11Z<S1S0]d6Z@Z4?59bq875Boh;2J0PaNN;OoOhUK
`5E4d[]<@NfE^h@L2FNRj@KUa0<1kX]<ON6p=_V6TP]gSm>1:e0IC]fXk4\7bDb@
=TXCmU]iXa6Wb<EU>gh?Nk`IVM8HmWK=`SDi]\l1GB:6Pa=eJo=GmXW\f9CkJDQc
3;jJ7<<@f\6DM9[nE=gb]T][LHMliTWK[Y7hl20EIBcej2qalDdjTJVFSk<k:N<E
S?ejh?ahLOSBF1[;B6Q22;41BMSD>=SjaHX]cGE;TSH0ImjDXY]SkgCA`ClFkgY8
6Lm1VH1Dg]7E^qK0bD@\cA>9aLmmajAbH?U1^3PYHYU3:l<3H=:j:G8YMW8PIIRK
FiONJDabf45>eAc321BM\[H>oJ5VR`fncX81=\DC9_fU^0W^k5N22[[C`0U1OKZ[
7Y_CP58nREALPZ;3N>5^p\k[_nCdH;Q<iVLWX:m2i_<UBfKEHd?^?l`V>mNLmRWh
i];4nKbLfm<DWKIFLkn?`_>K0Ql989b3C_MTm0KePleDBem4e1MY1R1n:cf5kEal
36=ONa<9NRlmodi4iBPYdJ>MJ^=pYje^33QhV=`ZlNF9jPRgjCWn9Y1g:`alMPTW
hcHSk2=I7;_k]LKFl\J1OM4Pa]?LOdX06R=4QICJ9mXAMSOn>bhaQo=YBWgCH_on
66b:S=3:oJk<F90eQ6EAHXOhoSBPMdRQ\XqGjG<j?f36hN?PnDjp@PkU6b4bV1QW
_6F3df;UJ7NRa;\H:hT3b[el]l6Zf`PcL_8J`X?0eAU@C\mdBbW=6De`c`O9AY^D
K8lKI<;Hf7i3d:RX[nk52F1K6ak;MZ29lQBLeMYIeKB`mWLh9WIb`DbahWqiPS1L
QcbGO4;RL84ZUgVHf>T6\;l8Mdk1h=kOb[E7k`J;NN0nbBn_Ze[3fPkR3;X2c>Ib
6gJl>MmYIfh92@9jf0>9<jAU=W<Hj@F9[A3;lYd5I@M?JEa7jh_IYK8J;i\:cM7B
6p5mTikdRANdbb>_P0Mho\oiFA`Id0ENioeo=dMl7[`[i?3=YZ_8=i0^CEB0nn=d
bS4jIK0S]=1=<dF8b?fKh1Kc`1]J7[=JPnZ]kme<E@AM]b[Rof0Gfd6MnNLN\HMe
jZ?jAWNZpNYAhmS[\oaKG;NN0KZBnOmJaDQYdKH`a<Omf2Mc^n1]fRL84:4gQIf0
Gca\LkX4=2joTI43N]lXdXMCC7Tgj:`YgImF4JliMdc^GGC857>VJhbWeK2m?06P
H9JdD[YWm4j:907p^UIaNO\D2U:fOPKG9M0dF]CIP703fE^AAd;j1?\Y:Bn>gKo`
1PMU_SII34Ri2a7QHG5lmb0:[gJB`E@dUn8mM]e2fk<WaeSCZT8aOD9gHTZ32AAC
oDhkJ5@ae[oJk>]bDG]ESeqQ62WIa[YOaCJH=mjNRkg02XL`cj6FdXQFnnA3@\BV
K27@TiE[7jUFDD`JH^>cT87S`eNZ]RTUId<o33WokRXldo8p90iWh;M1dGQ7JaSG
]?VZ4ci;9n]g\dJHb>eQkAke0@Bn@PKCBWAE8F4ZBU]@a??ho[beZNj@Sjf8W4Q\
>GI1cNRXP6]nDfhnkneDHjl=Nn[LX\_>jiSb\8mXEeqQh?<U]MT:FZG7S5A0icVc
_P6gLe_E`0bYFJ8iSUndWgViLQ`e][m7>oGZAM?3GCJmg5aRL2A2F6cM=i1SAaY2
]3in2EdNK[\L?JhGiMSdYle^ShDfZ6=kM3cKIpLAAbM`Pge4O4jkeXP;6iOcj2f>
gKXQB>R0QQNRTBno<ZiAPR3nYN0?:q8IiVT\T9a0BH:@]]nMnWk[Pi^T0?NS?bdP
J9MFnDQohQUM@iML6akJAXPfb1?JS>a;fUg24[j1K:ZBW]D;=Y>D5L2H?QJ6oUCV
J\;dEPQC:Jd`4im<SR2fKoojqA0eNLG>^9833a[>9W5m^mEH35CJ36hAP[5eT8WH
E\Z`iM6chG=He6aokK=nAI:;GWBMdZB^NA6DoWSI5>hb;:e0b^d_G:nJV;1eKg\9
`36?POZ_QeOR`G@aU^CpL7mfgCH:?h@cL]FbY>f8E;862@Pia5dF3Vc<<i0T6^H9
<\]R_7f:6kn`fnXb_\W7d5NfocDReC>o^:C;56R8dOkmEPT?q[Ja\]Bp`M1C@RYY
_jYD47iG4]7ea06X:[DE5>qIKm`5HB$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX3S(O, S0, S1, A, B, C);
   reg flag; // Notifier flag
   input A, B, C, S0, S1;
   output O;

//Function Block
`protected
<SfalSQd5DT^<FQ:WN_QYSjm;NZe2e?laI2P:5D^J7An@a^EfWXC=d8R:I>RU[Nm
`JhaJeQPogpPjCh3Ed>9>OYXGZh6]Hi3bf0IQ?bbOY1dbkaLfLh6]0leIAJkYP0Z
I]K6JGgZdZlImhp8;a`JIFoMkAG<W?K=Y:DSP61PUggdQ[5nOH5U;hBiX8DY;^?E
ZplM;>CHpj9N1_]g=8G]YfKEngH[EOB2?YT_jh?BNOUT]gFWEGHGiQgF<;KI76<U
NJ3Wp4lI^Q6Ypj7jId^q9h^L7Y^iga@o2FGSlY5IVn;^E1:?BLVK`=lN2IA0FARB
SOS3L7A^2SXJD6kVpL3Qc6c6CIHCV_Jo[<6Di42=Yl<@o=O_aWe>bfmT:UH0=JlJ
_FRfG?YL>X9>Sdc?a8aK0h]P:C_Pd97UPHdBjY<50F@?GH9622m]I]dJ9QLK[Whg
F<CLJmWpM0?Yco;SVPh<<HTd>oCU5=dZ6X3c]2PFhjCUa5A2ckVHLQkEYfGbaJZ<
eA:AEOYb1Lkbh23WR2d8_5i=eU`c^=iZ9EB<Njg`MlA9h`^8jAi`bi<Whn1Z][pc
J5k^L;B]7_?dA`E0;>62B\_3Un_?>3H9Y@Y:9emD^f\EN^LVDi@e]5\i[eRdhj4f
^>imJA1e=?R2?9ORW2OPBb\Z>XP_XQL0G\J[m8NG0]TR;BY6nC^:>qOa3GKI7BSC
`C0Y0Wnhf4C2Ak`BZKGhEmAPS\fQW>J95QBOm2\mn:ii2RlAae2eQAch1mLUXQ56
O;SC_Ic`bBTlK27IQZKDX4a5L9^5CkoConmmU092V2e7qe997<Q0UHjPWO2OMVnW
gKRR`b\:J^bpJ;@ic>N^SMeTD^Ue?4Ua:JCBDA399>J@T40M_O:A8MDTB2]HHL:?
1fDna[EJ`J3\kG21ooFIjle?U?ILa>d`d_<[pa2D[XSlMDcKTnlT:<ei1ck:e9m\
E3KAVO2VT_@Ig]:6e3oc56^e>GiAk_YmR=;3Zabc[[e7WSOD5Oo4g3:PD<GI33fQ
=GUALlg_6m9oLQ]_9G5k9VTH@M`7\VbDJ[CKoJHc39Ze8lXUPcUj@W[pQGC4MVDX
n>=P]4lWbRja@kKc8ge:>5meeFNP_;T[Mo:Be8GVa[675]lHYggjTGO\Qk9OVS=R
K380bc0RUaM8a[R`DKbEYamBTJLf<@O?Ejc6iRSDBLk_GecQ8kH5ZIEeaP\j_Z^e
;53A>O<h>Cq_2M3YA\kljAOj996Tf72A@6978E?kL4?BOmO5E`SL`UgB9khL^0a=
P0Z0O:R2g<c_fgka=O3dMA>d?IcAPbXlGR0KkQKg^4Q:[B1YHh=b4MY2J69n<J]R
3M8Qa1kIHfTOY^>`ZgKo\Ofi9U2JlqW1<\ih<CLPjeAgZga^Y3@ShnVRael3bae@
GWSncZTAb\jjN2X=4AJW>@@>]5\8j`WmD93\FnODPR>aTa[;Y5@L>I@I:1T^b>eB
o2bS@mZ:C?Ief3JlKYKSCVCK7HoYE=i5cDCK[94^Ooc\9^IMpf1_6;1W<[_FijnO
3\DTp0?6JcQdhM87?<1HN2`FC]8hhO_FmhlRbEmMkoNWO\C8L5Kgk]3OLSGKHk7i
f\I`:0YK[G]PJF6M7MI^W5Se2;IUlKcYadRR`3g]IK1UO`c;RX5Pm3MJN<`;DS2F
oF=ih\7;D3mhU>cU[SL;gX?qhb_m3ZN1UWe90XGJUd2MKA7hKW1c@fKQ62;FeT>i
kX8YOi<D?>LJNnHE40mTHge8hajGF[kU9XfVY5Ila6L<:\lcZbalmOKM:@20d59[
id0cMde@fDn>R>8;Pj;DaaX5iPlFS:Ea8^Y[an:ni?pdhYIZh282MEJ;o9IgXgO:
MMG9mLGBlIcO10V0]VgaLdTD::7^L5H^dGDHhMQFc`<d5?jn1W[ad:Ii<B:fbc=3
7TY7g9]9MI]PH;eGRemEQY:^4V3[B5kHh>a4M6nJ6]R<J8N3;E3g47^gjlTOPq`?
RMg?9mol`i0Fia^ol2\Eo1B`547MaAZHTE2H=A:fiKAVC^DOb`9>gcg^jE_26i`8
Y=:BeT8X?:fgP\JM?a6KXjQM7PLhaL:gDHS1A5dO@BXCOl?>:m:HA9QPjZ_=6=JO
EaMVh6@=KB8TG`^XqK_hALagKoUoNV3m6UHMj4]4]:^N`0T`i8[E[YmaSZR1JhWO
03GJA<DAb`f>Gj4I?K>i6_1103^M8dCQ9D[i]26pV44J:=]_1BV46^=m113lbKhI
W]oOYh\BHAo1o:WG?;79FmVS1ZdP?N]X:O?:hCQ;CDR`BBDP`C8BP:oAT_`0O>E7
OO8?O:FBAOQJ0Ugh8^?]7Z<3PZcN>G1E[@<R_V3OXDj2U2q>DY^bH8FX2kgeHL11
be]YlQSfF4;@<E@305O=06?_[IVj=5[[kn?BCSUmXkjR2_LK:cL_k;9d`YccZ6gl
bO_XH\FLCeSNeQU2758ZA[W3E\S`4@XS49^nD^d;WmIC^PLK:9JQHpnU<kCOnVO:
[RkR<SCY9GkZKm:;MK=jbH6A2l3G1jg2iZB]Da;6<F1Lj]?eBS?8Qc7k=B7a=AYV
0N;bk?;_T@7f`>_`B]d\JD:\8I6UT;`SfhZ59ZFKUXP\3?o@J4G2>mWkkSKDqOQ;
HinSbU42Nf[;a3fR]NPIfkCA_6iICkDglbA3UkXOMB\;p6c=3lXbUTcXJB[0SMCP
oIQ`PU8HoOJgUjJ]C_fa;XQ0TckWT3gG3XUC4F;m_M_6ERNY;;7_afSWV<YYQ:VO
BU8fT>\8HX4nJlU];fCk7hB>M=j:2f`NJ@5>Kn`c:n0eo6NEF[lp4I:Ajn_W5^F^
?dRVN^Z@HcRYJo6QNO>jokWji=IM3nI1bA2_oGd2VB@W_FDmIXI;91MOmHGo1f]e
U]aYCi=KS_V6nopJ7B19hhcD7D@mdXSUEI>MMQi_UXbUOg2a]AIR7k7RVT:`RGf=
go2><[gT7cTYmJBJ\6LX:m<IYKA5cAU>\8ae[4M29^MT^Qo5;Bd:oKmNh6gSYV]>
M4P`\PA74>OlmGCgEpC@B_=P5d:1<Z^kf53RFj25dE;D`?I1j3;SjHm2^QjoRJU=
nhLO5U6dNb@GjC>4iQCRMOJmX^hO4Ojm^7e<eUZeo;ecF=PPgo^aoA^P9:fg26\2
81dUS1Y8iUI1A;:4?`W1qOW[bU0g0YM@^>1jW\C^W0V5<C8mQ2cBQK;ll64jK9<Q
mI\8BJLl=0KFRFM?JaCY<O2R\FMnX\9dl@32bUTGDchMD4bbLl[RYLX:mGL@7Gaj
Y4So;A`MZeHf]PWbo:CJ331pU=B3Enhio1;81\OSCkWP?XKQoRnWa[]b;33i;W[Y
BZc@LHF>^bI;\23kAJDYWld3U]f3Lm_X^_gB7F1Bnk:fOF<>RDL_7Flcb_bAl;Qi
?EDj1P_FoY[YBKP@[QXkSlPI<BpIc@W^N_0d9;2_IncdN7dX\L?[aGBDVK5GjQ5J
@`X7ADM3ddU40\@4bmT]?6dI6H1:=qFZ6<O?NEcSAbVk;\ONCm:BK17@N:JXD`U>
NfiNZn_Lb[RG7N5UfoJ1?0GhK3W0KSFTRd><2U2JMWX;GHYiGIKmINf`TGk^@:JP
m5hRhR`5RVjY]U6eiMgU0`OBe@;0[A=KqA`I<J;oZ]Ae83H:VdDh=IP`5Fg6Qo0C
P3T=Jh4M@i:6fZfCPd[C_fdlLQZB\@oX7AXAfU:MLgoQ3eAneCMjN7CcUkUPllO_
A7B>EE0lG<X8@Q9IBWoe8`A^iPeOe8o[^`oqIQ5fV95HIH08kN?43hMiWgVfZe=a
XUeDSJegXIRle5O\gEE:E?@7[[=Oa8C_VDI:I5i_K350bMKA@^MeBm9Fecdo<cN1
AFUg;k=`hbK8inc8OfEIOReQFA@V<[4oFDlhW6pfSU2DihHc_9e1iTI@5Ya_=Tnb
dE^d670bK@mMS`G>HYOlmV8GMoFMCjScn?6IioEfIQ=^7l[6\haZ6NEX68fIdLQo
mhBlT=f`T94NnUFNYc:]:5^8^ea9XbEB=5\_i?WQmpiMAa0_1CI2hhf_6e=DWTgR
^J`_5njB[S7oLK0eY\:k>Cb<J3koOBFZdXUlV4kFILi4_[2RVHdm0oTY8K>;CApW
UQCUa4I9o3EE=f1aOUPe<U^Q>BGZ[D[n>_IFFlMEILL:eV@F<Ik58;9lTDoRAd\U
VaaB[7XAUP5PToi\Y9ABg<@H<<YO45hZVm^M4aT9e_<;SPGdI]Wkhqeb1Bn4W9h;
i3BD=6BJ@gbdg29M4;3SmRmB_X2:Z9VS@VJZ_\=l1XW]D]E3LFo\;97F9B9VZiPY
N[\;6<BFo>Sd6Q3QPYb8C>Sm>0Ykl]\AIA[QXkSlaI[aqlLonaTLELB`ZQZ^5M8e
6cmNi9GQ:fhS=7<]Ymc3\5CBVL4_OQNS?MjUI^0:7@]IO9hXWkZ8>\X@nXT5fg>U
a50d=3CkVdXXDCf5:eKQO?8gQ]\NZ7j@Fmbq]j:j7?em`MK?@f5PlUH1O5p:B5lO
PY7YFN5ChI36Cb?E_Ab1KjF]T[WPFd[>92o5>g^eGIVbC`fT7j:E:3D@;77UmbJN
f=:@0?847;0J2`a<_^IeIe1eUchfkS?6YGWP2:R0Hk9k1Y3>Sq?VKRb4DZ?8GNU1
0CSVmSgk`HISgcn>KUENLcdV<GUVX2WAFj__jCC7`0bBMT=fFMOk^aaGE0ETKJ9]
Ll@C5^?AH]pJ4gMKMp=HZoJDY$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX3T(O, S0, S1, A, B, C);
   reg flag; // Notifier flag
   input A, B, C, S0, S1;
   output O;

//Function Block
`protected
koVHCSQH5DT^<biRga36glT:29NpRd0cMPaof7T0hHGg[T3PA\?E6_hdNG_M3NMi
A0[9M_`Oc]=DcKp[LQc0cUa:hUo^WT:p=T:gnJpF`YhRY0k;dG@D[Q[9XQY[a6^j
0Z[gnN\f\@7?EWGQ6eAm7ho?Em2XOUa=doqnC?hUm:qo4W_b?pl_l82O9TDBN^cQ
X9\j26L_G2N2neC2g?<BmM1ZJ3EFR\^UG<>8AeVZI^_n40\BWWRmL;A]?HG?^O@L
ZN>m2I;lfBE?FmHLMOM3mo?miH`5U54hR;9T`Fm=1lj?qDO[H1d:>VLgEXI?M>D0
\WN@Pb90NCDfMT5c@h>eK?G14mNF]F7;6h[Cf>Qa4P:a>3>S3gcThc8X98KoL:i1
1UJ\]Gmg9:Lh_?Lc_aSYI?4e?VoScfn^]Ng<Km2pK7FIOi;IQHFPBmjW1kH<XXR>
Qj>k_EcdKWmEB8PCKgoXBi9M;RhVCl;^D6S<W3?9g<XOgk`Glc8n0GH@WG6b3:<n
doX@DRl_CMm1PUA=:`cNeGi;b]@3l>dM1[pDL;1m<2d57nG2jb\;j5@laF8ZZZ0W
XNBX`a\Kcb4KC;QWE<>WjUJG4RIe64c:2VolnOHL9?P;S?HmJ]>]m2JiWI\5<f1c
\BEkGa`OJGTK\Pii?1T@_Q:hTm;35pc[`VjQMQlV@PmTk3d8DFb<7:mLeH9Hd`^o
8Z\9B;Q[hS7VkOhg6BhlC`?^eb6mElBIi`S>>9HG>^V45A\jRGlA6J1?Tdp?R[6A
JjDhmXY>bnB0QpjEB>6e\CogGb^iRXXP^hne>jklD[]g2;BlOVdJk6P:[>=deTlc
dFfoMP8?^IM>3L;OMRWZ_4=^cEeFCKGk]51T6AlgBZ7G_de\Of3=mT=cb^OFGmmi
2M=0<o2AdQGXMZja:@K\@kFdmdE=gV=C0`YDqJPdS[B_`[6jI??TdK[mdc1gb_2B
0d?\aSeK8cGCmJa>c6M\Po\YSZLZF1hN`en:T`^U4S?3KF98J;be^iE2P<_bCi2B
mLfZ9eB7F[NW`]^[?AYM9fIo7_^FWbnli4f1CZ=iDdojUi^MDEOmhRR69S>3Jakp
5g@?mGJYWILP3[D]EE:5XF6d;L?0E[mOda`YgY^Y4bOJ?ghdmoB5P0`b;U@32G[@
WCdC_FAK4Xdj<WbeKREgV`oSK:Gie6?`J>`1Y@Qg=k=L`dUg@gi_N>o5Yeo_NiL>
50MW1XT<a?SGH1Ug`k:S6Ip8<1_Oma^;^n\ESHmlY_AMS^oQ25[2b@IT<Y0U=K[K
bchCEj9oQ7Uj4nMm1_XfUEGBK8^9>8\L8dZP?N[EeX\YT\oL25d<MeIE5iL_bl>L
4<7M\[eRjk>bl[CnA[cgMHUQbOP:Lc9BeH[HACCQ70\9GmC:aqI13T8f1]2CGSRM
R8G_^UNP=>g10QZ?R8iCA99B\>jD?hJM;\XoDlm[:k;\G63XQGK8\@aMg];Rg`[D
JAON1NGMmbm9WQRCCkXXA`0OB[^NiIJ9MlQO\D5DFM2A>INHObIVbV<?hC@in\Zj
KDF@k_?@plXVR`7AoBUbG5MinRoS=B8CRPbl;RWZ=@g7[CS<2?>nB2T=2X4Oc00N
N@?:k42?XIABPdLFm=j6]IMW^]eMaZXUHWblJ>E1njTWDN6WhN0NjGFlSoY5EgPG
MmI;\[9P;EB:5m;DEHh3GWP2nPFh^IliC@nq[L[f0m>oh8:9GJUASB[c859M7K49
9G0M<S\B@SHDRa\3U>2EcKaFLnXbVCb]TR=BJC:16Y<>TWB_]KQA?:eSn7BF=NZ:
DLIdfd\Z@o`4FR=B04UoM6bnB6S=Z5300_J2[@J?Kn>NU\mK^n7aCcRFBJp^b<ii
Vl3cGPhZh_H\iFiMB0`@Iffb=VBa1>IEPhDon\Oj=7Q]4oU]ejN42I`?30@X3b6B
\ek3Ub9@\ciFUR@gW>FgIffEf`VcDPX0?94b7`1TjmVH5@8]Bin[CQeiR[D4SUNm
Yj4aLMd22^DC`DUMWaXIhph8mL7Hk[`Yi9@1=R]SU27?iNBgmGF_0HWc3hcgLmZo
fD3k]H5H_78UXSUagM0iec?1I?5h9@I1GUYPnh0\6gHH1=?ZQXKopVbdTc7ILK6T
EV?EA_;f@>Mjn[3MS3B8F2imo1OFhK:>8KiRH_nql=go0>4:cdQOnF;?U^0HjK1\
NCHAVFQkA0X3g91k;`Rja6lF7A]0o<AFVDbD<ed;LXHjQ2:@]Z;M4gf]D:3QP;TM
@CjG^2^^NbmOV=;LU1:1OR\3PCNb39RD6afhe;o\5TUl82MB>4qUAXf8FGV;<0;h
=oUck6fGLm8JLHI=]U@PXUDIYDj4BQ58>]c4JL5oJS>eog=0l1[;03UfNL:j@;E=
JfG1cOE6Jk10L4Jf2RQH@in\AoS>a6;fQm?fHSB<c7Z@_j9So>I\U7=8Na:`Bq:7
9RCNVZF7?Q\]7e>l?FjSCc:?DPBJhJIYN2f1IIk?Th9\_?`IjXF23K>YAjB^cWa_
`UegMg33[1WmFUCa2]U1FdQ?[;O04nAf?Nk`PJ]fCKoKbQ252J:jag84UCX8=Q:8
Ng=gKDB^pCo^o4_X1DUc_U?La[2fCMMY9ChR4IcIEJj^VO5<\VlMY]Pfh^YWYS`K
@H26JYgEIM9j^1Y066X<CkmV82b;M9YoBQh:24mk:`geC=;N3c>4indC7bQMFa^5
KbHk?2A3LbcJVUYVacJqjocB^KdlbYF2@TiEQ7jU83i5X\KE0TX<KTb^KDhXG8UG
gYin`Fdofd[bBOaShnD=C[`1N\k6dVabY=`Yf3\Y^H9_G4:EMhqnZQ?5^BA5no9^
i;H>F>^o7XDLNJcBB1[MV7R0m0MNUl?9<eGi7>IJUT3P_1S??7=dlO7X6p6RA_PF
3fK4g<Fn<<H5:?>H]5ZD`K:6:G]bYaAS0WPO_lFllD13g:@4a;fdWd0TnDnH7ZEe
DBk8?lMSOah]@V8ZiISlX2=_cg_5YM@A5:?II3bUEMnaVebAa]lSPG7V]3<ADDke
4WBap<X[8UOV5mXJ:La_=P1M@Y?HcW7neTZHEobPR\Q`fTFnh^mE0EjWH2II6FWf
7S`WIEmjOoN0`bX6E5EQa0>=;di2iO?c]ea`\^XP\EH\b1b>d9n4bDUh9IeaK[<U
>[VUdG]=KCNI52MpHo6jFk7mbgU\\=F=54M]e4@eVo2n07[]AT2=o4Fi]JaE?0I;
YDg8;1k@jXC;XQoC`RRU0@;_Fh8GNg\8P5S68hOkM6fU^=`HHR2KW>Kl_a752;\R
B49HedkUc=TmddgBJ2Db4@GCl`qfK26:Eg`_4:jiW^5SkiAkQ`9EfP0OdWRNS[EQ
:K46n0i79<[H8^VVBkGe7B5]f9M^`h[OO[9OfJZL\5ia;CY<YgK:TcHHa[6e[[\>
e;TjnL>V0UJh4B?6XkQne`RBX[>RaCEQOH@N8pfcI1Q=Q4^_^LHoXB=1F\A1VBMW
a18HT9Tc^cKl\2PMBFg=^bjG;<BYLMQ4HljP_]b?kkm>@BZQg;HOd\JYk08@]9J8
ZV7K>hIc^jALI>Y]Yo93JIJ:1@mGLlI>XVlG=IdDVU2>:o;Np73`hgg4@3E[1Zin
E;1XhPOfH7?GOZV_oCd1EMo];b[Ycjlj\;O>2c5JF7]Kk;7PgFA<49khP@``AIM2
F>2>\4\F`YFQ`@lb7hC1`OQ@6L[W83X8<768@]1J7\Af;1C`UM^Pf1k7J<bpZlX_
Oh>\k4b;onpCP_<IYPb`l_E>54lKT42RGe7^=QKR_NAN\3SC8EdeCl\glNA`_`Qh
bUfn1fj<]cIZc5\`UQDV23E9P[RTEg;`RTmPb8nTf8Dg@329]>KB5CI60454Wa2c
Y8V5?H7G8dd0ZDO\Uc`:2qHcgDBGd_2XQfgHTIEGVDihP@BP?U>\NVVVm`=D<L^J
mG>TCF5blb2?=nA^4L@Q:F4GP;KG3UV=\B8BJ^7gn3HkRWlOPSN8F\2ZmdQhL?7F
L;^HfK3[W]\lCnRScO8JTP7E48bGZiZWqkEa9LUB66lkI^ghTlg;dAOiZ5W[o\Jj
:3cc5PT:IdSnB?=GkNH7IPbX6TG8\DNIk4De2A0[>V><3g;9E6PbCm`XcWJVfqa9
lebbm^QUmPJ9GRl4hj<7<dOkTTZf8ZlLE\U70RGnfO?Jg0>A]MSj?N`YP:<d>@\:
hTb:k\3ei7;3SLSMXSeUEbkeKJC?8MO]E_Ic:5MG65D@>SOok5elAGAcq0Q;6cLB
oR8[PQLfMJ83<NJ[l5aJ3c\Gj@U>nQcFNU<?Wa\0f0@HGkV5lk]m?Yahc2hYW\\Z
G]n[3bn?DmU1B=I<\MMifc\L<I4>P0396nCS2SfO]DZgm]?M4W1qLAZ^=>5`TmSP
LkDXSf0m_=N0;`8lCib@1\nBlm5MA^Lbf;cJWQ`4gE?`18e3`Cd@G=Z>cG0iIbbb
W:4;6L^\0?2dW7WTUMoDX8nPaDE>6G2G6_0G8m2]QAODM>p8^F7BS5CC`eY\0WcM
UfTahLDFHT`<KOYff5e7O>5a9GG7@mni5kW80:]<?5j@9_=5QW1OO_P:W519P;<T
n72R2Zc5ZO?Qc0TP758S8Ri@UdgO\RU\ZjUoC`iE@qlI033@H2SiGEFW`FN]6id_
>Np:lIh<=:@F5FdKENVNMPC3]RVDGaY<=8H>@lO3d0G?mAi>`V;_V0WGk6WI?8EG
CoE>VUm?ejiH3:nQTOX7\gK1W_l1E@1p=_PkD2p]7:aa0P$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX4(O, S0, S1, A, B, C, D);
   reg flag; // Notifier flag
   output O;
   input S0, S1, A, B, C, D;

//Function Block
`protected
WMgd^SQV5DT^<A4i8ggJM:P[R<oW00@<mOHnf:8OqRGJem\2J2MQfn6EDXRZ3ZM6
[FHVl_Rj:\Rm<OJ4]lk>:VNYGUCJ_:RRpm`]ICRCMch:nY>elSaYZ@E]^Bm=gd:2
\p1OQ`Hmpd@e8i1gdlg?K^HGJFM9o5S=8AQT`8G>D:egf=[OZ8QRD;V>lc8VR^QH
ZfOR8oMUfq<BVoO^4p\8GU;1ph]]9g=ST<OYjn?RDZ`A?mJXCC8[G?km=KH>GkB]
?mm2KAI2Gi:8I3=9oX0I5Pobj05cIH`bZX\G9Kg\PLL<ENhJf9KRFS7?6^3>NCNT
`ldhol:K4Nc[UA:2SRSAlCTMAQce;KBe`pU0fl1g9LQDgbQ0iAn:NIkKSED7S2m]
XQV>X_D\ZX]V<YgPQEb`ZjYU9mAlHhY7<QL2Gc6HJkh>oEZmRY_?3Hn5ZL;SekM_
Y\9iX[MO89`9X_9l8DWEW8me9`P:LVKA8;GUf7]n_cqLY_>Qhi]O7]31>6;E94e_
QXk1MoVRk_>BE27DiClJWEdB27W2oC]98>]AgiH6LUZXbM>31eP:WTK2kW1i2mPD
f6@kIeoClbEm^23ai_VcEJTkGTJdIEY__Qa2>h4lBMkJ7:Ko9CnqPAU0N=B50FiN
QI`0HS<PQo25Q@VDccNgZU8^BPb?WANm7FS4EkjK7ljM7=ZX5VEP]_FhIeJ8HO\l
5S<i^a0h[hbbQe>U_RY11682:8Aj`Of\koEP_YA\9[TH^fkHW0keAlL;R>?aq5TN
=QnOV0l3`V?NCmG6glmq7nJVT1:1YF?>35^GI91@2oMQhkNQ8nhgfCULoljPaVNL
[]d<hDEY3Je<8j8\L0AHeR3b[XBVS<e?KZdaL?`UK:>mS]FhW1I@k]UQNQh@ACS0
b9Q_aOn6JleFQ@9nB@;ffQc?R@I@qX]STT3UPFgc5PAQEDWbN1P0AR`k<`>X>45c
?UE]TU@44QedN]M=m6=VKm]eWk>[;ZYk?Wo<j^F2a1l9Mf1Q<gXY1o^N_^Mb@>@c
g_6J[W1M@MR2n\l?^g9V`>W>nlB`OTMBl=3\Fq7KKD_9?_6GB0<nPfhLgTYLDL7@
b@?;Hno7BiIN6=76077;D`_cd:TTc]7@DM>HloMg1S5n<CQi:=Ol;jGCO;`>AG1R
hlY^g9W2B0b6SELGiLBm`ehbEY@Z42fj4`g6QAL1T2:S5Pp9VKcGn44^1Mh_:@F3
1MV8`_5dijBTaEWccd9c@^]2m056;?Bjlih5jYYjT9AcijaMT1Il\nHe16mQkgB=
JY7Gnb@lROY?SFoH]d:B730ZCVhOGd`;:cLbeYGOI6TON2=j?CdH;lhqb_G2P_Za
SG^c90RUkEe=14`>K1e]5VRN^IZOCG@O45b2DY5;=F7fUieKg:aLZ7DkoLa>0NW;
C;F[0nb]RC]B47;4:f1jphd3c:aH?OiM3l;W8`ZI7jnPM]SS_O<NnH4kb3OSIIhP
4HSE^`bfb50bdZ@G0ddTGh0jG8X=M_VVnTdkNoB<Foi\J?N]Rk?N`<Phb`1Hn7VB
hSC4=6f[Gf_;^b<6<o0?lQk]550f:_R`M4PD?XA74B:0=E73\kHcjpa]nPnOleej
E<d0M>cjPNYNC<ZDXi;a^]d5`UnSIQfHmnqR04Cce\9VHD:`6I\OG7KIR?kX2BB1
a:<YEfY=GgjFL2L4N`Qh0?UV_aAL06Z8<YVRlJPW4lj=2kmHaPlNkF^j?A6V7_ea
l:`4mj2ia1B8WCbOmHeKTR]2?HhaX5RWZ10>cm4DAbg=7]OOlZkK:lYE>V6WXRFa
XTmqchE>HQT?SYb`>in?GTl;@JlL:UBH\;kjibN\Q?Kf65nE6CAe`omG2N<MPn:o
C3QOc\270ZC>MOImR`]H:APgPIg1a9NZWYkP;bJfcITm6Wg<A@iRm9R2?d;iFA6R
k][efUgKD3kbMn^L]>:CX[I8b9:1aef>WjY8q5=XO2[YiM[ggQPXnY82Klo>?En^
g77D]gC2egB74Q9l6aIl5m`jISJc]@eB=NekK5KI4R:jOEEZ=dB@1TC2XP=^XR23
fScDUTmTePe7W?h:6ACC^_8<ah3O8L[JonMnK01kW\bn^EKE[RNb@9m`n5\c[>V^
]S7Z1p75J30hBO]8GV<a365fB^DKj[Om4B5FQZ<VLB8m=L_n44KYJ_Z:>ZHYI8EE
nKc=nV7@X3LUT=:iX6I_k9_GG[e`TWU_0A4<QC7`NlPLN;9aT?<6:9GHj<\kG0Rh
i2kPWJ]X[0X85I:G>a50d=3CkViJ[EhfKJ4fkNpJ9O[PjJk7HMI28HMZ@h]V_2^h
NnC\Lh>[Wgicl7iZSqf6I6D]C[iYH\Kd9S8H=mYE6;lhi7:oU6ZHC^VS<;lZBloa
6kNEVMJSQaJe^9;kcjfZBLf03OE]GD1@WacJ:M:gm0b5d51NU>mbK03kTC_725CL
OD7iDVS4PG=nLQ@>RWIHYOh7T5E@3ja@lO4?S_CVPWRiUW1cHcqT6XE95VNTXBV?
2G:fZf3[04ddD5d^flLKES;:m_Z7A?dglBYc9A42UQcCQFlUdd^TWkQ_D1^VTGWB
3JV>FlU>J_AbOFm@8lUh2>]M2JVO@oRdG]mQb9i_;P?TmPSb[P4L9Y^?F^`Vfme[
L[G5Z3`6?3bk]DO@4V[p^8;NBm;_6C9D@XJSHSSY\bY^B4A^:j[0=2Z8L\]TGmEk
jhYOTKILj232aiP>BTZ=^?8oA8EoEanLH;`@h[_W;=hlZK2CS0[FA1JA7<GEFVgA
?Pcj]KJ5hCbY6Y1?K5lUSPCbQIiCESUL8Ld:8aBRm0a@Y`PGS]\[q3g=K05ZXMW\
VeI?GC3B^@>A_d<F29j2^l9Ml3L2cGXTCMOBaB02?LEf2\J[?[eE^3fX_>Z\J0XS
O5n_ZcIbeSo_`Z`6Y[\2D@V40@W<QCbo1k2j:3P2OXQ<V40Nal4_F?n1]^8>X0V;
XLF]nTKV\Z\7H?lhL[aa;p70gnKD>86^i3nKV;b=993[ef^SGK46fMHcdHdllF0>
2Ib><J?YiL]cHoWNb<9Jm]782S@l^`=BmHdFBnaCaQ03KQX7Xc4iffAUHL2HcZ0k
9AckR?edCMll\;5A9Baim>:=VEI6\D=<<[:VRHE@gT[>_QXOf744=XqOc?63cME=
_m3QgIJ]gRo\]<en7VhN7lHI:iC@=mEEKVK0oS@VY?H^;6Z_IRHF]_HObcK6@j5h
?KLYo___SnZ<[GF=cB;V\lfI4m4fi:R\g[5WbY]4RPn3`6eR99aHF6SgfIoGY^hh
Gen9AZhbfJ^P2C=4gDIV>Dep4CX6l@G4`WjCEje\2]HFS_>NeNCZSPIb?^pSE9V3
V59>caU;7KZBXD4542KY6>Y[n?72c_?N1Y2QGU=f;D0RbZU?2U[YCKi^9^KSGS7]
=eD0V?QhAmmaK_8>3QGHaZ@mm?RMMOg2^fS<VZLXUF=CSin2e2RRcfMf=i==TQL:
2iS0S0Qj`>llnE]P;hR:DWDmUeCpm1f@>k1BC8D:WDIc]goRSSVYDF[SKl7Vi<DN
geic<=A6ekPGiR1h7^^Ko6c;lnc[m^CRi6;3O8gPPJPdkWkE^l^Z>_Mk>=7Z>CBP
KW_5oKbNhQYH=2jmFGE:NEY32NAlh\c5>nJ2OlJP\mnGA:SI:_W5=VC5>WHWpTE\
Z:kIH19m_F69??85^`DHM`EMh?:nmYGTa3mYJUITn24^AX]]0GLM`6TRFV>29TTP
Z?V4Gjmn1eY_>o<YaAc\km@m6_hn>_ZBmk97f:h95E0oB^TVLb1Y2DC>0N<AeNMb
@70\Pj4I5m1D@cWEeWmhKSGD`_]IeqYB3EOmfcflJHXm1ZXK5i8322EdG[@nDQOL
g5m\:X>iNRTilGgDMTIEL]X9^7GY=NYRPKNOkUVMDI57gLU\?EXDET<30O<4DcFC
]TFT[iX?<`O<fF<5Mo;?jhZ4U9KK5YK1ec3AMeVPQg08hgh?9n?QgfJ>[:<Mo_q4
Y6T[V[MTBn?7H`OUSiiE@43j\^T]1E\o_J_D[DYRCOXd]6WCFUb@TCg8Y0N0hdl4
?RdBkIldeG@i8bL37i4]l4Cachd^=EF6V8WgU=P=Wl3:X2ki=i1nZJ^lSXJ=]mZ7
HnY3CCOdA=FI7bjSUnfm?E?KCFF^j0FqhYE^Wfo35]0cmceZ@1\kDR9hnc7;QEV;
\=6WJc2YK6C]nk>3QTp<cO2_JT703_RDbLOfeHheZZdQhXLhQlLQF;^dB@Jf>VZY
R25eUiQ5cJ=k1n4nDDc<m^gh;2Ne[nLiK_N8a@C?Bq7]LFJ4=bj]Kjj=AXMmFFG7
K4WLDFbAcGjBohEhdn4=fCDHI;ggbAek65FiKajjALc@QNn<`iA5<HdQaBU=ofOb
EG;2hRkKHj0ioM3iG?OEkKVWcIL6D@2:WT:`?a?0SH7B;]eEViL63Jd9CBK6AFZH
U7WnaNlY3Y0U[bpoai>5Y_g?n\=ci`VMJ0ED1Mk41kZE?U81RhWE4aH;:m5Q557o
2PTX^h@FBHOS3?Lkodlb8ne<5eJ<EdoKDf72kIMbClHam^=Zaig7cEh?kG><dI17
__`A2>cFlBW1L_loQhfD:HJ`RUc<NBWj=[mkVDDeIf<Ae^iZPDLpK6B:V[QE::2B
G`djbnE>AW7jR7i_:aDBTJR`AHZ=;lD8`THG_cVJMlRj8@L<3WUmoB`A]g]6WP2>
H^ND9Ahh[F4OROjFjE0MOARI;O`^=4KSHeZXNB7=R6@^b?k6RV?dK:=CI03M2G_6
HLPGNkn8EjO\`<9CJAPmO6EDqWi5FcZ4Hl;W1>2I>I<R6YiiD\OSGJb\U:9K<<IX
CVggTWR:;gV4lBmj[_^kZS32kdf4J<M0hjco3d]JFR0^oCT^G>Ni:AFgNJI@kH1n
6lLIEIBaibBW=On[_:a;2;HeOWk4<P9`U2kZXd\kc0\@<PUTJ5=EQdeUUJZW4qfS
]Xj3oF`CNhHNkCEiJC^B;K0W^6@h[nXWT5]I:0nbH:UK;4[XgZiNEF[;7>F4MbT^
09T3EBO<RjCAOSEFbQ[8IlREkNVlZZD7TA;ldB>9BA4D5jlKKH;l^^f0M_\f^=fo
dA6mHC57iCCDoY[Tg:34W`U7elKSl^D9e9pKL11EAAj70[l2RcnhfL?gH^0;^b]h
\UIBMKUV8YdCcKG9C77^@jd98fZOTGlUjIQV8O6mZnBOH^?eg2>mY0oE`903fQ__
AMVkC3DN_:nGT]2bfmn7P<YL^NZ6OMeY1S9K\LQPPI2^LT@e2HM[b=N6;AN\\obY
fEfkjI<pc>L3ji7LQK:]mke:N[4LTHNJ059P`7HN`h8cGl?d<JLmEH\:LL9]1bdF
]Z`I_4=iBCe4F5I[8e4=`W6GnQcfJmNk;BE7XY<9B?QCMgB=<ZN^e4k]fNQcD32G
enFgT4gRceD8kHNLiY\o`GimgNU`BN^89PmoT?PiBZWOpF=\WHdUe7IZjRQa?\aB
A9WcTTm?mFB?0R94Mm@2YSdgmn`WoZBH8g;jPVSVB?]PVTcM8mj5a9?XhL6`Um`A
V7>ZmY1oAgcYfVWT:7M\:ebLJ_Tm`eg^YUVd:O1NaZ7^BF2oR_=EdnDUlL4MS]V4
=_D1K=[>ASik7VRkIqKbOj_AU;n7oJOS_@h1`k2;mLoU=gH4nl\AOITfYq8M;Tdc
Jkmn<BOWHXhniHbUTD4d:QVo<APh][j=YBPOCNak@^E9ef;E45h3DbhD3aagdZj7
QVP1Z6\RZ;^b06U7C_@G4>``PoMh]2okFFVh`SnXWjmLMa`T2]DUJ7bYH78[66j?
FiYiSK\LX2nkX:Pal1dbE93hm;M<Dkph2ReR^i2E_2CO6OWR<llXhch8_@:D3Q5b
^5j:l98L>22B?_Z>^na>ID0IMJDl:YMWPJ]laI>XD=Qc[^7Kgm7@<9`_l9^PO>b;
45Z2TX<c6Pa3\9bkb?8I@FNb3ldoc?_h456bHTa:XY^c?ZNo<ge^H59bE>FgH1R;
?O3pZ0]M^X>QmbeH72FOJ[HA2QT5ifMo[SSnk3CZ>0S]7Uo:F=Ul7HEZJnGjN9RO
WI;_nVQU7<ha\7MeB<YX8m@8CUI:a_?eh>YPD`CDM=mMoQ?HehNX\\@L1cAGQ<`n
5aPHZnFCO8T^WkV9BJ`A[BB<S3KkZ8Qf^b83DT6lqdKQd9jaM9nIAd8BORQa<SLc
C2BM0SC@m<bd@oDG;Mi1;\WFdCNRB5^bRl@BbL_>a;7SKFE_[?bPPmN\_@l0O?8f
AT91CP0M\hi14k6;F_QK]EPdA8D3^DZK^aF`KMRXFdJ@><J<BZRSGm\FKO2\1hE3
8jY>:l8SAh27kp1Dek1X[QT3\R6WJAN85]e^EFY6H?P9AR\IKgIfSZ4;oQCi><<D
b69bVSC7ghSLAK2WiQCFI>a[[L;[dSebV^4R?DKX[nYT32I1KNFhFT[dej1VGUiB
lQ]=Mk8j73UgWC19Ti`kRgAhf1;dTMXlNJmQ2QAeU;L\hSIoU3qXO?aLj<Ie0]Ae
D:cU[[`XElE17AoF?Ohh`cJGn3^jfi6;T\^E<AoSoKSc;3N>WCP9CF_aBP?d\2lk
ck^EDdC5n0L[O5Nlc[Z]BcP;b6XM_?1:05DZEI=nalScX6dY6cFX[XB`4SkUgKNk
5eiN=9\ZTPS8PXSYAJb]M0?qJ237TH2e6lRnANVo8ch6bKOb8ABl^0OOV^5Wc[7Z
a:2P^CSAgfK=J]0@KacQ?knhe52E>Wm^`i1YPob2RDNBO3:d5oE3?mBECCEEb3M8
DoF==gB`V[H]V2jO@Jm[LRU^Jc=8i?U_LLU^Pf]VnB`RC>VC]?Rb?_=AC[O6p^DJ
ODIf^Ieo_?1>L9gJ`mDZkAC1bUCo_460HY0:eRj7c]2OGf;L3I`H4NoR^NC\2S^A
=_1d:fi^D58]B<1ceHjNUR29G7lFcE=8oknKC52g;BfI0F4CM34G:9LoDkSOI^9f
Ol>m7EEV>5aGI6_6mMNd^acGl@XTZEACLql[`dRSo093Cc5@cL@8615VdEYPBRg>
4V;PqS9^50XjPIjY2QIn`@EYji`J>f1cNn=?5T4gFlYmbWZR^DVHMB_il=KZ9ZlI
7;^P2T1CB^Qoe1h4?VP4_fLJ;8i;gB1qG^<=AokQeS`YMS4U;L3GoK5PNGLldD=a
QC81PO33@=kc\B>aZh[a7nB`2fMDi7hZ1DmP?:b`N=:8bG5=DQJBYNMC6>6RUSZf
6Z82ln99\ZSeLZ4emcE^H8BC1:kHchBMNAPI\`_]q@G<JSEROM=QA@>:XFEFGXh]
VgBPdUAQlEU9<RIHfPjd\M0[H;c3a4NQI2Hlj8kW`lkC2Qek6E6>6;fZ7>ZK2bB@
In=D]9A8@T79;BNAHk[mGd9Z3Yme]_ZQSDP3NZFa:PPdN?gmJqTfK6\b>?Ma^2C7
<3kObAZ[1In=lYXG^BZ6B40WQgpT6dgH7lbbbQ\546AAb\UY?K8i9HId67Ug9Zob
Yj_;NL62G>L@LUhK;_NO:S_[TS8eQB_`RQI:Sd:N<6@O\X2n]LX7fSS1G9H9lZI]
0gbFPecQKS502`9kCPoBdn\99Nl>01?^HfbqHbXe2mFoLO0B@TLRQPU@\iViWMim
X<A_h38_:g2Ge9TJ69aMTh4RedDfk:S5YM\[ffMR3C=O0f7;`>?M6>D`MjhBB;;X
366Gb`8OcH=;<>Le8Y^\CNgL3?DJfE]bA@H?@;b[g^]XqI5ECYI8nj8VMZkPUWPa
7D@TEOESn43RbJQoeVM31Y\XZhQGFFC;Q<Cn=e]bePnT1XJJK6SGZ1NXJ[083N;0
15l[k`flWYbD?>RoSGHcNGoc^?H9N^PAl=2eLl5h2`=A`af`IE82:poWS1N9`hUc
3]10R0I8N66[IChh[oV[OX37AVJg]_Uo_:9dP[G`87Ql5QgC8ml;500PDJe8C;mY
gL[fMI\P3M[FEV>Zhl0jPC2eA`XNL9YociL]7QX7P\mn5a4BL]m>h?YVIl:_O8pL
fkB9@A8`Q3iY;ZDTWk5icZ48U[W3LbI;YnML6V>m2\O;<GEEYhbRG:1k46fh3D?c
?NH\6NG\4f:4U9><AACUY@iKMYJ5Rf4TWnh2EIAkohmLaFIP9FUQhf;@50j_SK^e
HFGZ:m7p:]OL6ZA`YSdK5_ToaM?=d5EXD[??`0WZSn:C;VJNT5PC<0EVWnOanNXA
PIJeU1N?4kW?bjGd\f<X4SKOCQW3g?5LZ0STm]T\ET:]4_OE8BXY5nW\<eEPHfiC
:3^WQ:HR<l2^Q1==qHD_?i7fZ8abSJ;TGS;3c`G59OGNNn\F^YL7=8k277OF[JaL
7JNWP@Gleej6<f50ZcEY]_;<[V?4]K]Bbk?NOEc:T]1?FpJh<ga4>Ih5Tii@0PUP
G9lPdn_TR7=:7I>Pj@^S9A0`SHcc_PKDBBKIe:6ZhRUlFd\4CSC0QkH7l\o>>cfT
]1DJ1@WG[X]E;[o2j0K`oP8HhS<6WQe7>3CPe_eL\ChQ4Bk=L3k_Z7q1Fn1Fi5jB
_KJB37>9jlQ?EVB]F8>OFkO_]DbM3k9n0A3`hDdL^2Xd@3Oc6O@Q??lU9lHW;fCA
SodYYFcoHNSc\?9kbV9HiGbf;D:DL7lK_e4c^mANg<6UH29iiPaITS\Wog8>7A\p
jSjJW^A:S;jelDALkH62\cQfp[Scbm1]WSXigDD<;Im@Y\2RQYa2USNP6d;1;4^=
fS>6kl0DCm]^c_PQeD7[ON>VhD9EBRa22@GH;m8_>G0>\H^^WEfS=4;49US1XmPM
]6jlX:DSMgG5L^nQHK=]<[O`<ZkbdGMT;pFJ=dH>eIYmjjGY]8DW\eAcF[:6a8oa
SV<BbeD6S0;`So<[EARbgFL8@PVYdiE>\\X2<_bRFiAK1@TX]Y;<QC9OeZL=YU3A
QOjPb2mLNP\MFY\VM_`LSn:o2i^d`<>6]ng@h1eXoOqO;bYA:X:Oo[R\LNIT8=6k
i7C6BF=Udi0R3f9iN]`oZ:_P4o30A;W<RO22Pli=VCR<A?K6J6FcE2;?<OcSK@D6
Z2BY>S]W;9;nCf@=\baE3d=<KXg^[YK[?C2`PZ;jVM`DR?mJj;YqcFV=jTfeF>4i
\c4=o33eHNF1EU8;;\RcP9gf]jEEcg6OR;8gD\6Oef?ORIRPggaDRjc=eCbnW8M]
J4BS9UGH?`P<b_ealMECDGg4Nj^0gW]A0IU;o=:4LH?W:<7Y41EoMI63ZIh1qR1J
7af\7ROD:B=AZ6W;6k_G[6:Y>>Y^cnJAFWA;`4E[6meOgE?TbcdAhif42U=55GXU
D4iJ<`FL9kMLSd6nPF;HT?l=V6Bfd@^AS1;EgE[=YAKmYl>M4\ZA<Oa9:6<3`26m
721cEp7;nLnTeN4JZZkP2C5Z7eN3TY2l8PQ7>7]nb]n5Mb<H=b448oOG;Mi[9>KO
HO6OPcO=R3@@ZEKeRUHPN`o\9i6>LM7=g0DMJEUmb?^iPJ::c9OEbXl7DkZ949n`
\NX7Fl<Hcf]H1KpEb?E8U`SIi\<Y5gi6jXk3eS`J<jQjSZNTh?D;]DRXHGi[O3Yb
[]Z]7BT=^]KX1R3\6]dA]MSDKjOKkf@^d1Soin[`_BPpUPPbSl6QRO^EhdJeJ[f0
B9NCKbfo8Bq9dL4Y4jEZV6023gedEQEKl];2IRkOPZmaBXR=0j=`LdY@=DUkKfM<
6[1F_ee=8WO?MNRfl<cAG]ba95]UCNm<[:T2H[El?4aYieKNZF6YXM43=9Ocm`D5
b3NI35KOJ9T9Ch0q<d5nQ9R6L98O>?bGm5<95NN;TJ;9MVUc8_jI>4N8TNf4T<:>
cEGhTWD@R6k8ZHT<aE\`QPQGkaLd4<<^851oKNg;O57GL0h6UgR@RnFa`FbV9`Q\
gf=oQG1K<4W2@<O^<giKqWIYAjhY4O[bDe^C8:e@f]dYBLn@\k[i<m>S2d2\2;^[
CeC\fO>[IoLh8lWU77d6V1lULc0EIE[o3iU<:WA1<MdL@;li4h6iGfM;:]YjGVkE
m9WiQ99EdKc`NOk7WE89;W2aeqO^ZFFS8j854T615Z[1D>0[<CHU:mTW9c?\F_SR
akl`\k>H<Ho^8C68H>NYQnSCgfblf5jC@7koifH5lVi\SC@nL6Y\aR<^EA44g@IY
N_H08JeYa5JKB31PP2IG8;1Aj?OXF^p4OG_d[:eW<6c[_;3UCXgm3h`WU;maYbja
ID>gg`G6aRm7\hTcWg1CNi:7=l\:078;D<ENQ3DgIhi4I:7VDdIN3mUe7V7GSOe?
VF^;0<K0e661n>IX@mh3UD]:[^LIU`748cMqD>Ng[5g=RFHD;>_JV^e1R0Em]2SK
?0Bdc>^JCJU8k]l=c<2[INIMbZnm;I?QhVT=LZU81JF1_jKVnio>Mj[:E9;nWi4g
d_oPBmEP^JG=FC`KRO=3ZaLC?3\MO4dbC<SdDFaRp4`8gW[<j1S:?aEd8`RbFAUT
<<Ko<@bT<9`j<GYk8cjaCbbMSWo1@[AIU@A2Fa]KKTo_[]Z@\`]HeT3k<JVKAjUK
bN[0T\k2B8MD95_f1[B8P[l<CYb>G0M=MSY0hfHZl4HZZqR;JgEdL=G<lO_Ua3nk
M894hUJ:^E:iZRnTXm@2oiKo3TeRo9cE`TZ6k^WabdCoUBm:^LNU<821]mRZP7Hf
8oUkU0?m7TOOAL:k^9]gRU14I_Q]<B89C5JlL@?]gU?D]^R1mopfVF;VZITK78cV
GfYccT=a90COfVOobmj6g@eNno=BC^1_RG@TfaP1>djaj\j1iA7pk:AnLXWmmh\2
R5lh_oE4fNLBUfY;DeohTOil0\>]:oJaZjJ=TBM<MSa><^5IhW?@VB?QbmJXK`[>
:H0Jno8?E]FFp?cPXL0qS1N8c6<$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX4P(O, S0, S1, A, B, C, D);
   reg flag; // Notifier flag
   output O;
   input S0, S1, A, B, C, D;

//Function Block
`protected
o7;`ASQV5DT^<8YH3Li1APl]j3>^nVP@T6ooh6W4:nlO\K8bo;][76pfY2JoBD24
gDA8dW6X29pB73dijJ2@41TibUfgL9X@mbaY[TZfNG<J^R`b];FObhb<<AIM?@jK
Ac:Q`YcJ4Jkd<p;^8L:?qc0>G2B3Tb?^FdH`WJjk1cF<1B^EFIKb3CD@JnE6:SXe
f?FkOjB>R8A5O6[m_a;HkpPhK4JZ>qKB5NZQqh=9c4k8]81j=>R@ag<nKZiI[C1e
fNdgVVTaOpKXnLU[a8[Z5UoEUYHl\67@i:S?iY<PS<dSkY1=3F=C?`7Aj];JEodH
E=9ai]WV5K?W9=QfegT?diD2N00hmmO5AilemmX?AYg:kUPIgc6m=GV]o7>fF2@1
Fb1Sf<W[X>99EIdL1`pbm82FeLQlF1`^a]YWUSR:;@o3oHaHlcAXdhG0d]PcIlbL
LNDDjhS>P>Ma\GF@o_11[WDXojkH>11m9daoMbYA[1M6jKeXeWdX7h\NoH\Kk\oe
g;cfedo<0>bA0kYblo`nShP5JKNpkGY_`R5HK47OPWLXgKAYXjBIm30N^4Wd[Die
VI]\_ORR6P2jP5eoeVM=oMl_j?[6A^O<A90;TOni[QaRCSNBO0MVSTQ[XFh96BiJ
7_kkk<IjBfK`ZQS\I0REHnJ?Ci7med4J7ig5qRTSfkGMOdOSBP:LEf\VM<XijaNV
o_6KB7;oIoinUSF1]clhNKGVNTnl[b0BKa>MKB1Bd6]PGPS3OJS;=Y`1R`0a?U1S
>gTiK3OoQ7b4Cj0lFZj<oRDK\7IMN3noIQ:=i[l5;GWOFp]220i_eLKhMEj<F>6]
3^G7c>B>?6VTJZ[N^oRX\GZcc\kPhfdYkjWF6C[_;38SXZJ3h`b?31UMF>1VU_OO
okee5md=;0XicfWL^0jFX5>egVjD5^0n1I5i6IN?SHJ]Xa[Z_7ef1@q7`;6DZVDj
?Ngl7V;oiYYlK<o@\`d:Z79]<1k=JQD9@0;G?EZPa?@jYW08=\;QaR;B_LmVk1>@
^2Y=M<M>CR?M\3VeoKL@bb3SF1XdQZjO2WW1XJf96mD]@WYXA>^1h9:b?PUa6]_p
WDDSF9UiQP[eUMXThaWaQ?`ZoEnE<[]@dNjG[;eMQ_ZkjbZ?WZefZdB7gLcj36?n
UXj5I]<G[JNolTN2MiWUi2?_6bVf\nW4^jjG<K[eiaT[SG6IPTP_Y[I6e5c7ga[f
Ug^okD3ipX__3>GNN]NlIeihbHd\1\RHNTP[o_VgWEkf_cMd>KHiS>DB:8Jq^3Za
MMZD@EW9G0]U1eK@TYL]DjGkQ2eLG0F]i11c=oLJJ7F?C;gZYU8S_PFWAaZ0aa`T
0gZ\n<9LX1L0=mV^?`]d`:nC99honCF;ZO7Q?R^^LSol`bn9m=8W1cj<1DHVe0jc
NV32qR;n]6cnNHF8aF5SoDg_>UKhjJ^dhcceJMU6jIeD5FhTTQ=nEEj2Z@P4dXY7
2gF9F@YVWC7mGb;Jj0dGj`?ZW0Jao=RhKp6?g[O22d65CD^X=<HS:e@la@@:NGRU
VD<\L;iSeG@[BN2Gj7i[?_HF:g_f_eDUifh4J:Dk:3GER3bcBT^52fb5P2l1V6ZN
;XF[=San^8QSPO]\BKh[`28fIIH1KRLnoI6QS>91NGV;[bbLHR8;i<^_Z34V0:PY
KVFkm^qfLmn3fUkRA1M<=^2QOVXiZ;H6`Jj<lTkefXM<\FK:M>8i>@<F6ac<2PM?
[DXSgeY]jF1I^bGJc34iAV06P84`?U8:bk3KdSa^;Xhck_4fHWdR:=k^[ADHYQS4
I5:lTE0faGfA;dj@K]Qi>mhLO[9=W6J[mf`9229^@liqXM8GgI<U=j6cmQ@VbQWR
k;`2SBcL=0^RZ8a9CobZFU71`8R=8V7`T`W465]S>LUh@WQOP2bKP6gnLOD=oAkD
CWol`=[G7m@OmDFhhAnn:@X0o_0aiHWB`C2][MjIn=9NXncS`i:ildLNLn_B3OJe
X:14k5P]D4Lnm@=6p2EJaAh;DeNf6XRT47g[E][i5dP^l9fD<b4icm8<f3D6;Z;@
ANe<JUfa`i<RG6Zg?jNjdd<JeLV1Ikk3:8;SHCYP_VBoZ7B96WIM[C0`P1IHRI0J
6TbWBb?6<OCkLkbnE2A3?`\fCKSkjkOX?@QOl\co6MDM0H]QBWHcopMBaaKZTX[T
5jE5gTeR2QlYTZU?fOTgXFE:8IfSYJ;JjBaL\3e?8mCZLnD@n15K7bGO:Q`UFCZl
Wf?l=\S9fn1_1C:>=RLokMHd8CN=d17X\o]b6WGM>Ic@YoD68=gIOlMb4]UVkJEN
ZJ?m[Z:RlQ8<7QI6\L[e\aHAD<qG2MUGId^<KYam0YZ^9\7`82e07^QJE2mhm?V6
:Mi<]j7lY\;20BTC>S;L\fCQ53]B^U=IkhA9[WNEP>oaXo8gR9l3WkVb24A1g[SA
X=Qf7Ki]A8iNkAf:Hf?GlHUlK\QGn2N<l9JdA;=EMP<XE9@1KkM2XNZcF4Y1daOp
JTQ3nZOK;RVAI0W>AGcQR1f8nSfFoXC6e4LT5ICN1X=V=>4KCC:jeM:gHjWa1iE<
W1929FibiX^a8L[C4ofKK>k5>bNE6=j7>4LkmOjj7KH=NGAFUXJHRoH[RTHcnI2K
JE<o\7J`Z3WK8bcF0R[ImFIQ1nGHkU@f>KFeq?PZS8`DBK:L=Beffef1ULG0Cp]D
O`QjH?25n?QUK1g6REPloMo4o@ciOM>i^N84lOje4jfEPfCCHga@eRgRSKoKS>n1
SA7]M1E4^fB0?WLYTnI94ng::XM>A\f?^8KU@4FGKn::SnlP=<g=^mJm?egc:j]k
W2j?hHJnP`BA=aMCgMVR6M7g4X4cVSfVZRq]HdD8:R`]EU1A@k?QZdk2c=h^4`o:
?BdTSYNClVde2[F:LW2>>o3]eI3ceAUTV6NaQZFI[<E:nFKCAV_jDlGGK6X9ZH7g
do<CgYXcj:IKaY[i[hmlLTWX>6IISkDXf8O]TlF57I?D?DcCa5iNZ597oCg879nW
QLnC50opi?OFLZ<dJJ]SAiOYNHLgW7CGYQ`am3AA_n@^PQWH8>fR>E^b:4:Lk=7G
o9Z;i993W@@X4:f_fRZHU]lUSe;WTPLfUBWj]MWNJ1@7D[2c4OQ`?Fe0_?7l`M[>
=ng5J:cMinNUe1l:F=koUe62>HSCbI[0ni^d0D6LJ60kqgY]m92JfN@;egkY;_i`
V@<8Y`>i7b>d8Hh>^V8PWbeUgKoZIbU:__3fAA`RkQaZHC4NZ>CagA`9Fd3nSRJI
Fo`Z:ADS?XZmJAdSolS7k66@a;UElmOQ95WXNjVd1M^jDgold6oUn<GcmdA@Lm\j
dMQXMWS\oGb1;AjAiqmBb^hKh<M=k:G0[dkUKc[50i5fI]Bo6<2VHL8Fn5X^hZ]0
6b^eIPSCg74Y]4k`\Q6\1Z\PlE>_FA_\DX_9^?o6@Z76;2NbM9QTHUckFoQ1g_LL
LP5STj:<d9H?HO3kcbm>Sg8R_OKnVU_JX]ZhR3O31QYc8=43:aQOG<q[9L84Cg8:
[4YYA4L6ha@41\`6L9e5SA<kYWn>INgGRH;6C<E4ahJLBB3]FccO6_CAR]jN7`q3
V<N5fn]e2;9\Z?B6d5@\o7d<\U8QBLmP4[3KaIkHVlFXHi6JV9:PGU6o[6lia?9m
3K6m1CfmY<6^\2;DYl=CURb?mCH6`kDHgTAX6S6<AkI6El2BD7@[W6gf\iPVOgS3
9KbEA21IP1=^70;nSYEOUd1i=8Ln3hJHOd\pA\^Y?0D6neFBShQG9Jb6SCGQ^?C@
AcACIhEeB;H<Oi40QfR5_gi::geYWXFFA;FSJ6;omAcg;CBlbf:=AAaGIV>?D70k
MeFh?:ENOChb^DWIXK_TKG_F]7kD<E=kaojfA`C<blOPh_;bb;i=HG_B8N`L2;nV
dGMW?LfVqa?lkd3]V3h8KX>Lig?aJVKdaPa\?o;M;okX7hCc\o66S1d@lGkR3o:]
NB\fEEOIK15;bPf8f=;RM9=o`2WE8X`Dm5078M:4nZPXS>_i=^JEQ>2Si^7oXo:d
:4EGIeleDa^;cPG8GGG169g_d:>6dL150^Y<kPSGQZTUBp3\7:G6:h13iT[RBU0l
004kQf5g7AaYC=CL:8WnAbgeSg1je7FYRAVQG:qiQnHfBcIoP[2^fR\JXbn1Z<`g
_OZ?llm4`E]UbBkgQM33GfTnbHYC2=N]NZ5b[YNLj?\Q]mYMc\IQYX_bgafGUPiI
EW3k2@Id41@oP2FJgGSjGMR\3GPnm:PU`<n`:9DiIc70H?h;S21Q1me?j9j?W9nQ
MiXi>ildl??p>:=CiL`4hSAG1I2DSP7hkY;P1b\<a`bYEb7\Ze@b`0PfAQ1^E1n0
<=KVN8DjL^I7V?D;SeeZn0HnlZJID9MGTec9i?pWXM?2128S5H@N@TWJ^2P5>i9]
?dFfikNd9n2N3d2625=\LlbSBWhHKCM\L44Mb^PRiA5HU`d8_nNW1@\;hKJi1R;W
?23MLH<6VHeJ`?AYhOmA4P<EFDo^Lkbl_lnod=]1<F1kB0IN0f7a0bb;J^^e3eWe
k^[n]hm\T1EJH<aqQOWhc2?lC6`ScVD<T8P7E6GSbOK]6j63Li]fUfJd;^_8<H3f
nc3OjE=Sc3fiA\`02WiVOlRY<DlfjeG?ZRRcRl\f9OWJ6_BXkNm60ifTNH5cPUD?
4V22LF_<0mS7>5j1U;O@MmBOY`3g9NBlZP;:E6<H`\EgLl<kS\<S06^8pd3[4FmT
>^iR<_6g_m<Rhifa`R@JgYK:M26jC?O2d4S3HglT:>V>qjQ^9@6L1;LYhcS8UR8?
K>c^M<QEl^8m6kI_gLbES=a9j3a08aABN3oO=EPG4Hj:iT\KO>MS1[3_AoBL;1]L
1i9GKFQjeO6N>`00PHSgA5@oZCJQ\HLm8POP?XemMAgR=`XaYA5UAYbli[[0W1n0
1>cdRa:0M;LQ>OSM:HMB]pYTlgL9nX=_;:<6:]06Lh>U3\\5Q[EOAGlcPJ=HS0CT
VGiZi\O20eQ66ElR<X<IJ\cBFYjcboX`;h[7=0kOg9T;ZE<5R@>;e66dbC5A23aS
YN5Yg7IgcA5M]L]caDCiaLE0PlaHXTVHT2>adHkIEjLU05VmXPf:j\3ENK5ST4pk
Ak:No0Qc_oki1Dk<SafEAhA=nH3HFMnM7aI6W\eAg]g0FBHG@kh=MJAFaJR7jSbV
Ih`\b]_0VLKa3R7j<QfU@<EonH31f0lB7mHDn2?EoiiLjcQ?\FhSDL:Mg`0m8169
J5UH5W`OdoBNS<TjARJVA3\gCkdUohcRUV9D^CdqKZ?e2SI_E@kQV7NX>i6k]S[W
m=cVKdSLWe<TcX6_g^5gIGPa?SM[gnmlYY;ShlWhO4K>`B@kfJ;=AQoLHPH_QkVQ
6=Jon6=Re^l@WVV\flW7ZcKB;M^i_@Yg`XTUngOZSffeU[EFN?C6Q@PUHVa_7RZL
0g5n69`VBG2BW]_?q[R8AWWSd9YdG>`>aQSR<d\o\aODm;l^8p3a8dC5=hP8hI0O
:Tm:[X=Ue7Af=oe4_dZjZH9?m^jAgH6PSCH7SiZ@nFli]g>LC:JZ93h_CQ0TBVP4
O0Y]W8bR:M1fa@6`iL1JGhBb4II\VCaHl47\4^\o]O_:G51@_9F9L]imIcFk3Yc8
nUY7087UGeDOkU2Wg:f1IlB:QfpUj<=S9K;>6dAT=Enb8`L`NQb?:nLV?TVABEF8
`Sf4Ql\e;K57ja6CEcZU[O[\:GUfk3]GWAJBR?GelcmaTC[A62LP:fUBoN5B9f9L
h5DJbgBM=M[ECXZmUfNEWEUN>cmW7Rj=_1IbEAKVi_<aHV[dNU0Gn^J:]8NiTiZL
7;kqG@:PBKHK@bJK?j8RBDoTm@j09[]h<AZFS2@nKeKM9;dKjK@m=i2UcUdJ[jA_
dRKjF3TnM6jl66JRkNfCeGci]NCMm[\UT<bl@YQakGX@6ZW\>IMNOmJU;SBgh^fY
;k@^`a^760?71>M[87POeIE9S>g=i;7FZEZ6gWT4kVNOqU`Mo:lekKS87^0nggn:
U`g_ZDokS2Z\RWi0:9ZOZ<fFGlZX4T]Z2>AUo=;[NEG[i3P=6UlU>M5XINO`N3Of
=coJo_on^KS@17IPemUQ@MZRakH3S=c8IXbTjnJWYA`S=n\bnin8dom36U_Wo3MK
UMThbFDkG2UJ6DGTVmX?hqOg@@?2M8CVg8^6d5_E9:;PgQOaG8e_2La3dQQ<>S?d
?BeV7_I4lkK5O1CbnFkg=3EhdBWhX0If12LO;aTObBP]4`JaEGU4a`XJ3^ViHNaH
LFThFJ3aRmQ:<\o`CIGV[9cKdnXgIdM1^nPlgOT`@6\P2ic06VM^6]V]bOVc?;qN
f8Hf9SFKk1WNU:UV9cUdWY=Z;FHc>>aeNUfE2LLjZ\fmLFC29nk?hUiW0Oe02AHF
Y<h5lN<aJCnYHSCL<1\Gd_YM;X>6HQ`6Gl?==3mLA^A`0cG]D90WSMN:j=HE0hd7
][GnGZ@^68OYSbULNo\m4CCWkc@h`VFGPnO=8SZq8AN0L6i?kN<OUQY9kHUbKQDa
X9CM7CDK`8hKm<mZJg[a@BKD1iQ6ZdoegZNM>AX\d3oBLV6J^?;\\7XO6k?W4iHF
h9CnilnIDhglG5eW[j`K=^[6TKBUM1DkO@BXiH9lcoKV9oTM_NM_Sin=6Qkk8QH5
PB8M7RZJ`5PhG:4?qWIYAjLOKOmbDe^C8Ho@BUdYdLnM\R[PSm>S2d2B25^SCL4`
jOTFEa0\S<0N[fF[^JWZN\Zc7cJ9>kkObjoX1jnFH_n?>lAB]:bi;oOj]2?gVZf7
R6cE<6cb[cf:kT8lQNlKTc5ORN[E:iL<mj\GhM6LF;li4kL;biMGboQANq2UJdeb
EdOeGbm@3C9e3oe^=NC^4gMdH`WeL0[C[XaeAGA;GEBYTWY4IJD@?HETXU_T>F?X
DYb@?f=WCajbHW@m40J^K?FKQ1TP=bjK2hQUmXcWh4JFT6K80MOf0?31kMhoR86A
nIAj9l1ATfjJdWbFPElZkQk6=@o6c5j3TCp0bNd7G=[ciQ06AKaVZdJS2ZLiZ[P<
f?iMM_m_bHWI3HaSF:i=0UKL5J0p^ZQ\eAe:D7Yd;CHE>=mP]nX7UHSk;fFUnc33
nHXUTSJV]Mkj=h2BOYiOC0iO\k>>]JMlk3=c5B9hX?P@=3Y_H7;:AHScP8=gegn8
hXgmmM54OmMSX1eW@99N5YGAUmFV8=iTFWn8VDQGgjX0=9=ionEXdU9GV@7ABe>4
hU=cpGkXCCIEMn:UATjT?]M8:fLMXi6OlWj;1_Q7RNcGcO3g=nf1CS<[;5ogNhIO
oS<EI`=Yh\_52GC2`?1MYM`8[4=U]=c69Z2plHbl3_ShnMMSk0k;Y\T]GSV@C7NI
E`OA6Q\=1O7UfKbZ:ChimS=5I:4nRXWa_B122;^4OU?oTTNG08o?hkn<3lF2nAHL
Z`=RCR\>X\lZ\REcVJb@g\JLZn43Z_3_f[Vo7bZi4dTIq6nUQHSXYd[hoiC?7bS\
LXY[LPcbE^jPQD45<TIFb`AgPkk38ao]jZAce\K4PIKmhGE^ee0OE5Xc[7SB]KoP
Mi^bd><LDF1T2]25=7M5=U>Io\d<VlUD@E\cFhP5WU6:;KdVk[nAYp9e7P:OLA;h
N5fd\eRI]XCF@Mc=@dI]7:_TDKK[FH_?:oWjcjcmN>JjY_G3@2VihZ@C<EgI[g^D
@6kI_VDd2><b35>h6BJSdP3iD>L0[Q99BR6L\0X1>_=@R]e`E9gRFS960jXV5Fq1
kM>LiLWUNTjVmEg1bD757RMk_6ZX@9JTD=RYL9oTAECDQ@aS`fX\DZXM7HXkN^<M
g7mGO:Q`UFCZlWf?fEEBM3A2b_Z:DdIiU=39?lQkO02fGliPW9l1XZoUgWY_fO?T
IJ[MHY;qC>N_S_7`=YidYomUU4\]k3E^@_>_9oj6_\mCO_Ha46ZZA:MkC;K<ZI50
Q3ljF<SN3];Lg6@=dJeDXB<k[3FY>IIOA3]Cn=\AmhmAn9QE<`c]mH[4O2l]Cb=1
85hoYFEc?=K<3h7Mq2gkNG7DY2=h?[>BfDZ;kgOOF15NH4`?UIg:1b]U0i]^GEFL
m6k4k\aZgB_BQFZ;@J4_LEf4cM46d@XPf6DPIHO7OAe0PSkQ5\=:85m=m?UjC\lj
K7bkSRAZ51N[W]a\CTDOHd=Vkpkc>J@?ViT2H7ln:MWhi2?5D4VW7kUBKM1WJT9l
A2A[B[V>fNLj:Ooi3>NLcBlN[G^k3Kni69\==Z=B1F7F9DFdE1CB`P1IHRh0J>Tb
WBb?6<OCkLkbnE2AFY`\fCKSkj3\V?<fM7q;^`eJ:nV68QNb@9?i>1F2ik0T_d:7
J=nn5o[ed2LeP?JeK:L69CKg7nOdlj>IQ@q:@5M5;_lDSBBccDKe9dgXnKRkXI<R
T5^mBHH=;2R\J3K[1m7Wn:805A09VefoEc\ZB^jAXCP?3PIP15e9c;kmnY1a7o8:
7VFLfHIih6Wh10m@A@[AI\=j:BcXAmcN=Db7j]=W@Voqec<CgM8;dbFYL@73c>1>
IKej\S6W8@K7n9l;F656;DF^o`F5o4T1_REN9@^b?1V=Ki`XA`BnGJ\J3lX8Bkdg
KK9McQUWqR4ANOKfPKU`CN>:9Tb[eJ3;T[[>]Vj;oe7J]FjRA;n@>NFdSSP8?eH7
S_A2<0LKNFb]g0nADb]2Peg0bQKPEbXOQ=`Y4l;nJI`JK20E=YM6nUXkP\E6@\47
MM=;GV972@`0@n5BkpV4c^UbR5Si_9Z_o12mM8i6SkY1BM9_oLV4DXO=f4bC^EVV
;9\g[IT?@:]U04Gl[^fkZc]hCcM5=NKLJ[0U7fon`k_?9a3LhBM7Dh?iR4bV9cHF
@mDAf2g\=DFL0OiQB=_H;VM`?ApIa5Tn63C>Tm<A<07HdKZ1fo2gWQ6?HlI0jXe2
F:T102IIca:=fAmIa:YU_M^C9jAgYb=U0d:G0k?bEW]NJ1Za^n=_<OdgALZaEX2c
l<]:N_MRQ;>k1adi2:cdSVkUWM<0Vcc@IcOq0QUiTN<XMPhkkkh^]oPBL?9S<BSX
Bc@>k2G4WU[]17[I4@7i>>=l4?<SS;81bJgC;k>BLd@PJ9J>I<@HhbFCg=MCBX:f
d@jlKlGHnR`1oMaK@jh`U_ll5kfoFTZ<E9@CS@bKa7k0q13C\B]aFCT8Ul[>bP:>
7>RnJQD8cU4JDBPMeW<LhGBbmjg6dHJ^V:B5ZP;5OjG0CjoSZkVoH8`jIB6X:FQE
^ihm<NiWS2>`CVOM5f=8heM8bSi0SiGlKSW;Qn2B\0\bK_bem8EaGq>VDYm34R=N
<0XMPZkDakKb]d=bR7?0lo=YK_nWQnFmoTVZ9dYfCo`X`6>C8B:5SPFdAEEack44
:j2AG0[R^m18\edIfj;mgIFTK_HGk3FdL015RM`c>:<j`]0Dd]R;b`on>EVb1dqY
Y1c_BETRaCBS[WV>`EDIhl8k<8l55nbhCX<fBoZc7ceckKMnN3SD4cOqoeF]K34R
6IoJmd1CFh<Ch>BX]FAk5m<Zo0ViY;H[hAY?RgCEDjAoX^A`M6gf=7\AG[20fQZF
;e\_200BL<W[U1=5?HS:e4XD:eVGBJ>Gh4FZl1_QL`WZAVA:lVXTJcHd=<d:79;3
pR=WO19JldVf^@o]QC3L28HagT5a:Z^Z;\N]_K@chR<`PH^^>aZf3W6XCW7PYJhJ
Z[1H6Nee9=UdWjo`TQnM>1Y:D687c=ONR93]gmb[URh@iYA6n2J3hl:3lG3hiYdd
[nWkgcS@Ap?ZPWQ8=m0NX_D<Ohm[Q5Lk]HMJehFO5SB[fWK]QC_H>0>9agJ<?L5]
lDUW4kSblO>gAfgOX;[i:DQCSKSa4IOH4eid3cpF<mMeQTXg>K0[4`O;2^S`F132
3R<@hUJOHfC4@PS84MB68=g_32nmNJClFUmP9D>jBei3km8JYMU1g8PgXdYl>Lm3
g83>AYCeRfj4S[6Z=YF3753m@mBUYJKK<Pn4InWXI7VMCM5paL]UB35mM1:FCC8f
iGN?IgbDFN0f@4MK8UcFX6DjCh1M`]UgK?kCN`>C3[Zk>6i6EO_UgNh8d=ZHNTW^
lj^d80f]j0`_GK_Q@2c`1PcG:W?\g573JNc;ncL3PKLVBFeX;J?3cmWaqTaR91Af
d:<KPh?M:1T1dM8:R1^<WZF4OiY_ee;NBLNOCYNDU?YTnNAlWdYL?0>bMIhF4L5U
R<5Aj`Oncod6bC742P1\N0CD_iX_h=YXQjMMhZVaoiL^\]YlJZN@5C^f;3V1d3`S
YqcV>OLd;9UNYCCk?CUT@X:QJQEHH[C1:MWd>0N4MbLj1`15V3FnH>ki59P:VOe\
PDi5:Y]BPnbcFIY_0CdjjG=Hf<nG;JlW2g8S>bM6I3JKjI6XhFF3e`j5K[o2dRbj
14a]<o_G6@qbV`]DX0g441hS=hcT__^d\Id@WGm4PVORO;G@Ygk[TUTLOGlHeI87
]QXCdb5]P7`lCOnVCRm9\_G?[G35VKbn;`hHbAj0SGhjP;m25iOhFIA\;oYAc2]@
K2n>MhgPK?Qbf>;Uf_lqg?T8kWmU>Z8YVaZ_<opRAcSeDiH\Ko\nl_Y:hG[5@V<K
CoiHHj8n5h=UjjPADfM@P[9990THKZ79nRae9<7SVDm[ARDm4^bb?^F=YIi?hoO:
Kh>FeI[gShk7`gRXl6<3Md_^oS\G6Z7k2HRJdZGFTgN<b;6p`\YXaZ38]f^9iFi4
AQ?XeNFW[cJPWY6;WO4oDF4KiZF`:nnP5m91DSBBccDK?WdoXnKR:;kh:@J6W]?b
jUf59b<WFJi9h25@<24UYAefZ2LJjjkXPX79?8Bhk1PI9G;cmn5aQ]59qIF6AVkf
PjV9Xol1cBYf[EK\==A?:ZFi<7KfMLcA\6[_mfc@7h3bU=K80OF:N@8L]jUOSDBm
20>JQhQf@E67cjS0FQNBLC6WeW]fFeBDVCVcm?oaFff>BhZOMQcSj6G9[AWK4`MS
Jqi0;WVCb8baFU0l:MMDFX>oC3ifTE^ZBlI=HU>;:T@H_Q35433PhD:o:Z4]KWF^
[Yf4I4`cobZnMd?FmojRY42\J29`oOqO54V4MpDT073UhoG2Kh>RqT4XfQd3$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX4S(O, S0, S1, A, B, C, D);
   reg flag; // Notifier flag
   output O;
   input S0, S1, A, B, C, D;

//Function Block
`protected
[Y]0RSQV5DT^<=I:<F<JdL`P@iG[iBPCi9CEZa>N>o@;1^lhfc:O^of>7aO<JKWG
_P1pS9N^E<PYA9a\Mkpf7\7\4anEJU9j=YS@RJ:K[4HJYn9pNA7>7?qS4FTN]?Pg
gk3XaH?HZbSFCHK3HS98n\3Kd8d;B@\^DBk5VgL0eJ_S4bLIk\gRV<7qIY?Pe@Kp
Ia@A?>qLZj<0d;[M<k`H8Sh[[J1]RB2>=c5RPUn7`bG_^2SG4iM3Y4>:_=\GacZX
]l32_4Q[CC^M:iQa:`MN78OZ\UbZQd0]868XRBZ<8bO5Z`4GX^]3gTKDeSLJoV:3
dVJP]?MadYb\g;kqaDRE;fR[\<_8SJc6dX1b0kU]`\A>bmeQbBeX=<6KX6RQDUcV
R?jSL1VG1;7XaOXF=fHW2HcCLG6>GHj=W^?AdHVjFfm^=G3amNeXXH<@N79[AS=J
\:VKn1VnO]H^nfee46AVYl\Mp@;9ORl>[;>oc;a4NoeE[j6Kl;?P_\=Q[P>K9HRn
k;<oK:\Z=7TLl3GS163XgoMRFg_>DAC9=OK4RbB1R4AP;ZSkYIWFjac89@4K@CNU
`PQ[f1YoN6a2:>D0Jcg8j@?Ba2D1JdKdfq\la;aC_BQjcXTE=3l[?g_lTS7\X9C]
783QLXgV2XJHi6]OU6T^;[`>g>@0YF\>mFTVFWGTh2=WlNo765DWCfa0@ZeKgM2T
W@2VLF5:5@A;VaMg[JdG<CjBo12e2<92XOWGBUmX<Op`3M1:lj\>8NkPD7JnRBeO
GP698Nj<\_U;WQ6]bmi`V>gAD\nNB[mof>ck=fm>9nL1GZN56L9l^VA<[`<O9Df=
K^5>0[U@02f5JQWU0<T`fcPhYU9H3I^Q\>O_6dnamYZHcXL\T3VqL1CDc>UCPA6G
GD\L845XE<o\KbPX@@1Bl=N61;^_:G1d81qEJi<h>F3DA;;]Na0BYm\6cae4PVA3
abeo<_EElHB53\2mkG\NcYHmEbIamdW=5k`PjoU99H279Y[BkLW@`CoCM8:D@bL>
0c>Tm_ToW:c5S1^<Q`@>ggR3EbO:6di]kC?JA__1bX\qoT1=iBW^AD]0SjV4NIn8
gaa^SfPWlgeL:o8INoaN<W6B@fSkLaL\H2Q8?2Nc<fYMdQUHWEKCMHUiV6=mS`m^
7XPfhAm2202Mo>8GC5Ld<WHJXkE;g=@55IeW[2;V;<GIW_7lTL@5q45?lVR17h?R
CG7dHmn5JTGTfLbOPRIcRPBJIjN`;dEP?H_fdCk`?Si6\OCD9MddmDUiDM`gM0F4
_OT:U=NB@ZKJcoU`:BA1`j2JaR73IN]T2l?n@801L356C7Ui<AHE]gO3E^5gLpd`
MEGYWb?V>BIZ`j55d6UmNcQ8n^:FD8=ERabhTAk[HHQRF_KJ:Xbl5NoNJ^2\6D2h
3AeXo2kOBO@QchU_^Dd;O2FemGqX^3Bj=QeZ>DlBjF>]h6aRHEL@]lTWm=RCMW3n
_7`IlH;Te5eM>0_[2IO>gAA53RIXRBU^5oHEi]mgUGC@T\75:oAdWCZ3K=mH1`bm
On5mLIIMNmLhX^@0SBVnofjEDkcelDM=fQlESi\7B5i\@Hb`IE]lJaN3M^Ap3GI_
m\AZ9DB^8TVJS\Fb1_]dS[@F?d;2_aD\BVY6`^WYBAgWkYT1:WgS=^C8hdGA3bDO
NFda@neJTPc^LiRD2oYI9hj4LL;2?flFn6:9bho<@@2a_RZ2ZIVEL=6Z_8;7<>Tn
iONk@icn=CN\A?i6[^`Eg_8lLe=OpQCgb^mSlJH;\PioCP7G`^?I4JD3c6I<::]X
=OQL0RK_S94;W<eXd6bnFFASEQcU9Q<S^3;cXF_n5K6bnDeYm2mC_>HSC1Q<OMnU
2n5\d0geS\iI;h^GB2`Yl9mnM0a[8YBR^`AbLFW`C8hUESa9o8gV:Y[P>1`olq`Y
[>E=kGJ^^GV5K2OnaWGTgMl84VUML;[R?X2WmVPeX4Xc5L=Y3fg?LNF_m7>k7C`W
=WAFKWZUMm6`8m7Nj><IGadi_CGSLOk\f\Vl[mA]ZJN?ILIjFkbCb`g:@XXNfT1O
me8kUJZ[X^CISGc<<AbT?COS7cGAT[qmnA61f@jZ\WSYGc3gTC7g`\Zn5o_d<NM=
jmQn8L4?\<oJoeDY8D>BknT4;dX[QW>L_DqGCJb<YO6O3g_H]WShTRTS8n[R8nVE
DZK@mAZ9O:b0j1`AB7V\9c;Y;a1WXZD:n_KGe^Ti?7JQ[oGl8Ke_nS]@N03ENPCC
dZCFKYiQF\24EU__[V<E0nEbTIO12>Fd8P5`jONg3bOQhWGnG]li8>9RO62hg[SC
nQSpKPH1U:Wn9>HgXTIRfng<VV@mO`4@6XH@@>TDh;oo:C51Cffn32JGKdA3[>c]
9_FHKeiR2mOo53NEMJ;ajnLof5YlaZiC=OHc<O:6lm<_R9=WWYajID4MI6g1^ee;
5WcUlMH9N>f[5QM6kFLI1d27^HM8[l[j=1GFpL2kXME2VDDJ@JXA@Nl\UO5X9j0K
`E;EaUc32ESYFNbl]FV3RYVV2KnTQa\eP:<S7LP0Z\54cGgeNQ4Wc1j5?OC8CefF
7DIE8UGYGK\ll>>VBEg@NK8[olOkgjTY:aHm[^09bbT2OGfFo@bCWES^Eh8O1Q^m
7DBcUp?jO2J\BCS2S5XmZQ9CRI;K>WAXCXAZ5\h14HK;RaR[D<JNNQO3aGbA3M:=
TEkLCE?`VmioH[d3Q>KOY94\ZMQ?1MhRoc7V5<]]44n<OIXLR5gmVablH@3FcXEJ
?@dmI\liEBLgBodngnWaSLOKC=kMiY2ST47MlOqiT0K3E@d;_CdUkSfKSgif]BQ_
]e7h2J0cJRnTeBa_TYWV7^PR]RTBVKmkBiIl1;0i1E:^SY9U;EAY7m0kkZ<\1_UK
Wd\NKJ\FfX]>QDj5`LVJ5@WLo^N0[T5dQa>:JA2OGaEl<jRUlQQ]f0c@J]8^cK\R
ENGN_k;qLGHk=M<8F`]>A?c0N2Yf^E=e4:UWfhLSR[BJ<3IMgQK\Hl<_b85<TeaV
U24F\l[DLW2VX2LQ@a`DQZk]aB[6=1Il[Rkf_gL=SEVQflcZ\Z;^@\fTPY5mnj>o
8=K8GMCYQT^hl;co@a5iOa6bPR8=XEAUcWP]_fj^qgGnW@ci=TN3FIY6^JgiZ_Dm
2@0n[0JSe`5bNhMbj2dZm\WjL2K4n`c]XKDXlCY8h5?Ep_V=]M[VhFOZGODPYA;_
YPC0B8c\6M3@S>n^C5NSo[=WADZg6Qbm[Df1o`Ia43gH\_a8<lY\];m94of;oj_L
`_ABA:ch;Sh@UC`f4e<gl8A7aHf_V9ZQmChhHL1e\jWJd5G2]0<]^;eXL2eZCWXg
jFfP^?7dhSVTip0>l^L3Xm`<5fhcc0=XoTNl77L@AaAgeIQRU3nT<8?ZhJdR@R`U
4MfVIgE:@n;;ZA0ch`o1DN4f`LMkDa0?KF\Sd0Qfl>aHeY?3Z^XA1`6eL<=JVI4W
K]H9nRO[HAL:gd7dW0OVB:4aM<n00F<DO\;;V[MZ1LaZ^cq>YPNXjn_4<A11a[W^
oKCm6oER3R4YRlJnjL9m6dPR;ndCH3]W@EVoJSd7VDZZ2Z_>CHJH7bI;VJYon^M=
WRLm]>ggN>8V>lmFPTa@Ei_=5AVAL?h4gaGjAl8\`75nkjX1LjeSM3X;5>DK;X1K
gBniNC8o9DMV68TpUe]m`4PkN8IK\A?m_JohIh:aL3eUKaE95oeQ?W1AhGN\9RGg
\<e9cnLb5>lo^MliUUSIAF0>>BJ@1mdfeoj<=k95V;icJSEJPDba]en`?cn8;<7@
ZRI:oPG2@KSh]JokN@0Y^XV6>?bSSbm3202`oCWf]U45J:ZFqPLkAL<XG7]D4T`o
aO2^TmZ@51\YQj;?eKbf@3MTo?N]X:O?:jTBin;hJ:mW>[CaVPZUPTPCZdh>5P0n
>SSHFG;3TLTKS8C?eFRiUE7073b1=U@hYh>3c1DidKefH0RQN^m59na3Bd4X2F4;
6Oj\B3C203RLK8HdepKQ:1dd8Q:5o1doelCK6Q9ZD:3d6Z5F1NR`CC5^`GI2XKUD
QC]df4lYF123UoW6@KK\ObikIW?2QHIRF`M4=d6KC83JG2^`1<13`EZkNWanUJZ`
BkhSKm6A0=c7Wn]BD47gWfgi@=?iSJdHbNROZ^>@KC5=mH^jcTp4OB;YRY`m]gFb
MSl[59;3e71b4GI9BBkhLYnq7QZ;68@ilDDlNN2\5oERC4TQlY]e\RcES:HVJ>>n
Wc<ERPX7eJVkMca_9WcEISAO79dWEnaAVAb9>D3I@QaEmMpAJ_CD?bMjAHK@::32
SUo72R8LGC3g2P1;[XXb?dY5j<hd15\RN`cQZPj?N\DBn\`1?YAONG9WR3Mki0Qj
1XP[84iFd:PgmDE1nX48@?M0FOG62>_^S1ZfJXid9iC^CR7Ao4[k8lE5R1nk@NQg
CV1G@DBE;A7HM6C1^QMqbfNWnFa1egUjicm2d80eX[^n\9``Y`:X;ZE>d^_QF\Q[
i8A_jh[jiD>2MQT[AeLam`FdO]AMehc:kjl9Z<X`WU<eU0]MEV6_nM2_XO[Jjn?U
gj?ED<0Ro4Y@`ekAEcMlb7E[OlGB0]2ekUTLUnTCIBUO\E8SolF2n_M[qOGh8DF9
mm=7VV94Dj<YT4fD^E9Z=11fZHU?^f8FoLj<2SOhNP72F1d6E8J<Kfk@T?1OF=b9
N_Ze1lJ@F^IP@R=g>OnH0?n^Jk^?k4haM4I0dV_cl8<=YjTW94@@cg7XFOI2MZ8:
\G]JWl97UgBNncmTgMiP1dHTMk\E@pU=[R4Y>4Td?Q3ekGh2>021D]4?PW25am<<
l7:3e:]DHPALl=m8:1PHD]iI?01=ZfBoTPmb3dB@JBjILoon_h>bW2NJKcWOe_42
Ne5KJ[n6cePR?AUD_hgZY2<F\599\mUF\ZZTnlEco4j2>[gHf63_EO9lYTJ>G74m
TAqhJA0U1\Y:nL^abQZJ6ajB?@Ap\1XO^LhXGS]`cNn[dK=WgF1fbmQf`4b[[NGX
U94_UZLZB4aKoa4JHm87VC9FiCZEJ<KIEF23OPg:G6Q596U_>Mm8G0oH1]Keb]GV
4k<>`c>VAjP3jGkfTMUXDi>^QFAb\Q6^@132FHn^GS@9NTT<IAb3O?mLfELdb2Jb
p2[V]RRfg`jVTWY4Y2cj@oIW7Kl1H77TIZ1WPHd>?1B<RBgamkC9OInFMjL@g<\b
IM1DlUhAQVlhfmKaULa4TKiX:d5LJ4XHQnEhRii1U5iNm_:XEQ2GGkCDgTZP>NU7
^2H4@VW3N[aPAm8f@c3j]5`]LK[`ID6ihnVW4qE>OAlRKneX1]l3kU?DRIkVe1CF
Zk272]`<^>5Aa<3>g24`n8:6BJnSa5^8=KRbNkTQHYWcP\6VV20`U@neaiRdFfh4
m_6DmPnoL;J3`i6F?X@5k<EN9o9?2hlX]4LYA7EEGVXFd6bi930LmQ:Ym@fX0TE=
ClYbW;nJmTqVAZ>R0;ESYeI3]IANJ61ckladHgRMfUBY36]993VX=dVfg0Xo=J=m
h78R_\X11kX;WblN`;I:eX6RO]]TYAdOo9AD70]aSMZYMQHCK9IVbXb<[i4f6Zj<
8AjAL3_YjoBV6eZKF\oE;65RfCM32gn\8gbRmFM5eb\YT]@pHTgCFCXoF9g4[W0g
qUE\`cLAS[[2Gc@Vm^eg?18@aF:GU`L;gUO;`FCAMg4E?2Z^@=k^6Z\4@AE?eFk7
O>f4VBmbiHcbooVb;<bPf3o>jBM`fhbOLW:;Z:I6oI09_f>22:GQ0KDb]U];QmWE
ZUeeP2hM8UE1QoYC__j=>kH?kD^Jg745>WZOopn>cB;M3ckUWeU1CNdK3IT^6KEa
2A=8H5`BiS86KPM^\TG4ihIY@U`VQ?i2eclTkHn>7SZi;oBhMn@DljbReHjcLo<S
F\@HHCH<H^7COi<0in77Q;ljHEZ7[I0PTSnOBjSLfgHgEgB_b\8^4C97LY[dI;]W
nE@_S^p<4eHYaC_`T`B>C8BU5SZHdATLj[o`dmfHRZ:SOQ>CDgW0[2BUf^]CYCEa
iW>Da[S>5;L>eLNXePPUPL0A6dl1\@_iaHg4jlQnmZM8@6WnSm?Q1C<dWLj=5K>2
GOi@=lb<31H2c30<CQEU<gQCQnI>2UG2FNom2iDnj96q<5^2S\n`]`VQHSL1?<bd
1ma;HIZYYlh78fXQDiHoHf0[:4diqnhLDU1N4D<TdW0Rjn[a3ZN0AUl8Q]a[gB;j
;BZ5mGZU@@hAn4JSh7GK2VkITEmfSV=`@EQ?CUWD[F4Rgij\NdGNb0J>IR@05>Rm
UDOdTH?f\EWRESJcKQE6;Q`[afS5VnOi:O49>gWUMFOMgXOY;M6\2RdYB@h5a>`j
:p8Ujcai[2`V6]?EVF9iF?eOlXVh<KO6=MZ@=WY7PF^3Vd?JHS=AI\Pi8_;T=N8e
E[8nj]a\Y0]<b[PKG[Lf?<;DMQg9b_=Y=oMCVfd59>=G:KaeURkUgO2Vh3Hjm6Lo
nJL9m]>B7=]fTWL;iWFn7Ne\=Ji?Qe=HDRqPo>S]nln4\InE<NX:JIUOKS<?Q2JR
ZXWWee_VNnbPodkDPbZS1;O`QTf=OK<9S7CEJG>^B_h^R1d@JTJ1n<fnhAYl[OB3
cYYS6e;YLZ[5@e^if;?CN;eiV[ZaZigjV:gP7D[2R=1[TWl@UeJ_U3`]ch\eS68k
6ZgSRd6qgn`iKA;5<8XZC6[b3e\dmNaH<n[bA_F13Q3IcYIdEo?O<c_aEMg\8mbS
dIk0LfeX^IDP`JBA:OF57R3lH;mWRc6:7K\B63C[VTQY@W3f1m7fHfc]1TMY5K9a
9LC0PmIFgN6BLdRB1\A07S^3VKh5==3Y<P@<HM8_VfhZqmVQC9;k`a5iSYWM<:1Z
@n<oQ][D:cm>O3IQ5RC`l5le[OJ6OioCNC:Y6A4Pc`98VI^lIMPKWUVl1:>cV1Oi
TU\5k3T@Y=47^:QWjOWA2mUXZhPSnVVON=UU=md7^mS9lm0FCa^QVjfN5:26cnQG
TccUY]V0HTNbF:[4`qbUO[6`>a=;:_:EDhX7jiCm?mUn3:5DNAlaIg`aINPOSimn
3CZR08J?jmP^XeQjkAaL=RB]1:\jaP`kV\1nKHcBH;PSq1n4N7;UAlk6:]7N_Xo]
I:2==:mHK3_Whk0j=8c0^MQMN9iN]U9KTJDE0<k72DN[21mBT^5W;_n;d7E526I<
UEcm`no;Phla4lS28U]eIj>V>58UObL:SicZeC]JD^KdeqToToj5?lVkHbLmnJN\
57HQ36neU[`DIQ;BL?kIlFqc?m3cY=6jnoSZ;D]g@3>lTULC0E2DSBYRA8Fb^6C[
FQ9RcV2UjgJCf6_^I2oBmY0ca6WXLYA4h\7RkR[_Q=Ena?G_n9<@k[=`Q<F?[L1e
EdGjg7n6EZ5cfL:AOOA5LUHqjM\6m1[2^5@k4@HE]A6[JhM`^JU8CmACbSmOJhOi
\Wc^9Ybn8iVd@mLR4[3NhooIj1@[<b]b1UA0bk>aaL=`ATKPHabZPG^^^o\kgf^M
dRm\:DIi^8Na?VL^;Dogk\?5q2<SM8YAWb1;0DLU@P7fb555^?;Ud>6EnG=;nCIJ
Vlc0g`XCIR4oYb:0NZGdXjW`42TE4fCcbV77X`SBi1]41`QogVX^R7?f4Rdh_<BM
=9aaaSgG]YP_7MlA^CXNAL1T;pAfinMh;UOU5CjFgP]k3oJaV7NdYSX<]k]L6<lU
9M<W3L]IkmJ8@40RNH=oe8_1CAADE>^2`m?nhi[Th2]Na?M]2DAR<SdcaN>KBSbb
4HF1oBQZaI2WLOX4cb1lUf>KZSqVWITQ>`mmm3;]7oML_<g\eej3mDf>SRdnI9nY
oTp40?Rg9Sej[on<68XaG>J61V;Fh@9ngh_EXRmf78CW>c64SFli=NTV4Th<8R6n
hC04LaVjng80:R>SAF2ZdbHl;Lall5M]70e>o\O6SDHnlQn:MgjSU[kLnn7^KI[L
bNopV9?\AWGBi5oYTKg:2D3S^l^kT3XJL]\eYn2@WN`X78\iJ3hH>:@BKJ^HDncj
JL7GVR[gfSLG?IPQWhLhShLI__?`kJ5][?lIQakBDKehAB^c]g9m^=W:Wi7Zlg`4
0<?mq[]mdGH7QR:TacCDQA<Xig:>Mc[:l[2<NkHf<;Ghc5c\?9dd\4lh`1g_5[e9
VEhCe[k\ChlQZO>i9aHS7=iEkAl@@L`<OI@geeh_liMMe[=3785?QR3PPh8A:lKh
DZe>2p`BOJFdi1^W[106\MeI?1CgG6_]h9H\JKO3Sk2B^[b_a<6^^;^QdR6lOcg[
7Wc[`N`0b3g04XjAA<8LSkSI6BpocU47GC[k?DH`T<Ghm347SZP]55jR>3bEoVGf
WXCdX]X\2\nDh15Dfi4W0LNVDEF5cSmdH^h`BGk\RM7Qeh@=ekd<?14B]J62:<XW
9CVecdI]XLYEDe5S;IW:dd8QIk?o=04q5ZUGEe=<=S`NegQ_U=jV2S0l2eUB]0>F
<1Q@0S^Mn\RM_ANQjh5TO=H@TlMHl0EY31H\c`bEMd;<T:9]<l=m8S`MnOOHAJB^
S<S=7QjP[U=jS=aei1On`USePZ:R=A_j50_hpA_R0Ihf52\mG8HIHdW8TQUdVVFJ
]ZB<Ql[HmPH><1hV8JkF:gEF5T=T?kO]L`<CloaXDdOZWgc@>]D266Cn?TUmY0m6
@[EdPd81XLF?5MXiimOMXoAniYXlf:n42aoHeAdVQp^:kXEB3JF0gYD5faa8^ed_
RC:>DF[gHa6dda:L36i`B?Chc7SmXj<NlC8LWcOYgRG5[<W@OmK=VnPD42M3F]Ia
5X?U[LbB;n@0TYFn1_74<EWV?fXXk2:JP9dVSjhaUY^hgEqHf[EKi=2WZBJi0Z\1
ZF7aTL9fIIU6JOdb0]iBEW[DMS`IRkh0]n92QXTAkgf3ccdRB[><nXZFCk=8m5hC
a60DTh9ah8;<o[FJ=\]]U6;oDD[0[358KPXFej==l9:Cl4MHE85qg=9kA><nLMCT
j5KDKYkV:i2H3lbVlNA^a?_W`2:e3KbIKjk^nD9?Y^knhRoBpmY5Z`e[TH^RHNId
ZkRQ3NnkK?=7MOlFEc@]BUTA^mAWWS77P1\87XUSYB<GXAjnT:TN?8hRlX0f^1k7
Qm@VWAB0`j9G\lTl`Jdo9FP3nZkiCCn8m6XeHY22UF3`BXha_mIWYp3PnOHggQ78
dnQH[k3?L3465<^T1`WJNba[Ci;cjWX5\?03HS_l:>Xhn_562h;9BOaBFYWK\fj<
A1mZLFQ6QbS6BTIMnLk743CcZIk>HjMiiRd`jH82\FKBfmbJd[mX:R3?V:qF]d_J
?R4[ZROCYd[L0ZlL=5i:WoUl`ck5I<FP_nB[T?IT?U`NaUcHdO\SoPKEK^jV3QoV
cZbJGXfFZK:GOnLXo_OTCc3Fa]4G4I<9Al<g4Rnb7V55Tbe8>W\8MDA_LlWFTRWp
iTnY]MBBWlNGmY^NoXmlKIEeH8^D\njZ05L0DMf]Tn:5:kTgV2Se<^Qe]j17fA^9
nW<YKkbITYG=o?<b?V7ZnN;Lq?FdCV0eZBNjNQ9I91>?n3VN2m:=M?]>C:67AJ6Y
_Ym9ffDZU2l@KBQkk`CZ^@Zb2?Vb;llQ=V6a\YfNX03EQ^b`OIEn\^C<ENH:T9]@
_hoQ[``<lQBK5aTebjlb?5AF_pQ9Og[KMXFiZY9DG=iD9Ei2l1`jbVaQEckHPgH_
=<dgm?5U^>Ch4WZj9J;aJC>EEfQZJlcLma]]Q6jIb;lUcjaHP3ok?3AV`MiWkMCb
5j8HSGHnL8NVJlYVgWTGb@GTHmqb[<=DXTTnDSV`VbX1PB<WdmeIS\NWO_jU2BG9
NO@<HTdK5Co\1K^@E3BH4C[dlXKb=_OdADI6K^ldnWhag8N2<WG<=Oj_LDW`Q21O
2;3?McR7mf7FA<N9g4LIl]Q8Nf?pXPRXIbXWB9CkgJ[Im@RYGBngOiF[FQ1G>:fo
8Iho6^9U>3PfV=C;BEDfCNG4M\QfXRRHIWFXi^YL4Q[a261R3Qh7JFlQZ>Gf<NnP
<98]l?:0a8GE_V3QGm[DT^T>>CE4p?RDYLhR9NXa\9KdmS]2e]VETiY1q_8TY9lD
CJ2ddPl7FT2TK6<BYddEE79k<@;I@9Z=72]4k]V4PZ;KH]8fP<d[LMZRO_=VCon:
\]?P8h<nYnCL2=P6Al]gcMgJJ0kUcmF1SORF[>kZk>38>cPiF8c=nCEOeq_a^^Nn
9M4FOXoP2Ji8QRZ`X^n_7iPORSDlLX[F3RDfHN=YdUUPNke4@>1DfEona>_`8=<H
D3k^DdgFhD3BeEWTQ]LhTd8]X2FB_4m6WZNAB:O`X>GdIRbEl57Fca[=M8qC@LEP
ci3oiJITSMk53KTXkZhLDZGF=@abYFa4AJ]jk_DiIW[]mG]j]jclnbe\J>dCA9N3
D0IT<Go:k000WN]O39_TV2m`BZEWlPGjTUlZ[?<aXOPhG=Dg>4Gj\ZB^BFEqe]9P
PfdDU]6EGJ2MgeC4N8G4LP]:LA5B4ak9FiBgU0BGA;CRZb1V0OG9Ld[l9m^MehHd
`d7P4P0]@NAIM3SDC3N?13GFhHRGI4?S_DE1Z[eF]cL8RXlXCEW_fjKD=lmMqC_5
3EPj=RTlXJnPiN?]SWZkAP]Zn;f6B<XLjT4EVHj:UoQkAM4M`i@`^h8N?L]XdC^6
hP9<UQBV[j5YY_FjfpP2I6b9qa2lHXP0854A3?;lB<[gB`o9e1C6ei<\GP4pC3F2
kIB$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUX4T(O, S0, S1, A, B, C, D);
   reg flag; // Notifier flag
   output O;
   input S0, S1, A, B, C, D;

//Function Block
`protected
E[FO>SQ:5DT^<h=`7m?6inpJ5Od;X_]\2M7M;W9R2JNA@G4`X>Qb52>F^ocnjhPW
V5PF^bRe__hHonXI[27RCbkdMQVp7KVDKLKegd>;AL@Q4BV=?1_TfS5kP]eWJ8C4
`IgRYgNm11qRe\ad6qm5JUfJafEi[@f@N<CP`3SoO<N<54Y:^?hN[7]R<V3cH:T8
7P2V[bQ>1IY<j\PbF5q6EF[]OQpUlKOnlqh@nUUmVZINUE[kn<_LoARCJdije6X<
T:@ESDmGA8g1j4I\NhCc^H4<W>_@D;alF274Yca40c2;M>7L256k_l5hXPI>XO0O
NZ6dS8ZmJ4Ooh_bfM9_Io_1:Tnco5TlLX6Tf[9gjj3p>8KC`YNabKemQMeX?ghmM
H=42=hAnZJo[YiWS:aFNd^8Z[OOfVS^XI?njAA7fHP7BJPGn1n;mBJ=NGmnQ3gKS
DDZZgTa`lhU^@iFC?g^cVET1:0e0moo0H?C?9AEEDD5GlW>J8FgpcDi`hA4[BSNI
38V[TBZ_0EcZIm2ZlIBePaYbneb9TCA7Z\EObBl:WFe3h_HRh\HUecjJ[CeQmRFo
\2@ZoMbVl_aB[L02XSB<l@YNNBF<VMP1SISW?QFTn>bo=?]@fenBc[N=e7a4p1gF
S1f7TQZQ\9`DgkSWoEmB9A0>JnYBc]GAq[d:f_iOdVGJgma28NEGF2LQSRI7oHo@
kAic>DMjj;M;d9hgcb^7jdk5kZPfHi]1l?dMYcMmD<_2LgOQenP<I^\7cFQU[\m:
K;@cK=l9fPe3@Q2XnH`[E8?oQe0Q5K9AKcWP]_nCjp;>KbSeOL]G0Rd=mKg^5dI@
EJDh]2RO`VMK`LThLc=mJ<eZ`_CI3I`1LF\^lAYQF\]amQ5OTHeHaY`bMUoc06K[
o^]F0PgCHBN^`76fP0O3kkKWHljhIDC6Lf4@j94J<jDA?<HC?4q<>dLIhGaB^D82
l8_@6Jbobfenc\MKIlO@G^gIk;1h4nAQ1Z\mGKhPC@UFj2D?giJEIH;aWQ@g_<kR
1SA:8M8bbNo1iTH^4@8Uf^9gn?B^@ZTM5jQl5IMlC@N_5GIoY:4cn44cjN8q5F_W
TRQ@=oC]MhYWmVGj;b>PcJ3c:kL^;<Bc4m?R>Da:flZh[2@LaVR`[C1hRW\jlBPj
Sfg1`]]CGE;noWkR14G^lC<K69i]1bBN>MH1GiG3_O`\S[U?`\j=WGZ2l;f;i@FH
Kan<qP2g5k402:GeAdV^eoMdL<kJDC>FT8=R[h@4AahiGHJ9^bZSePHa@oe__FP<
RHT><SS?YB2C;EL2g@m8j4kk_@5R[cH0FMSZK@V48k4[7e34S:n69boOnGh_5`N8
27mbSG=M1=9;hq\MkAiid0B=Cg2=a<n1_jj^TEWQV<`G1_g268V;470CH3oUKL;E
DgeN15Bmm[3odiJKj=cTF:FR3PBCPkVQ\o=3?jUR6<qT_dc[=RnTNUboZMX1?>6a
F^NZ`Rk5l:J[HnJGgjj^8KgFYWAYG`@?4o``UL]7F?jUoe7K>8hSOG`=<NW^gO:2
T1\O`g4>okADkQbgWO8d_2TTo8OV5>[7n@aHj^a:Oe1NXSNKj2CQ9FTBH63^4dHe
P7Y`EeM5Z]8\P9mg1_CqBkbYM9_7<QTQILLjZdkZX7YKQ@daV<`PH^4]@U=jZ0X=
jUX00]8Ef19KKcAAIIoXlRR9nDN?OPi0Jbd0=8JlZ7]5>@do`CBjFC_EZgE4E:6`
2DTIEV5cmW=Vcg>bc3P?johnQb6>hYYL3i23=FNR\6HX<S<KR2ii@AK:ZM99q@oV
3Li;Xc@@AhN]YGKKlO_;kFJ::\Qp]KUdBV2W3SbT[Kd:G03bY>G0GggR`ImRnQhR
JWm7H?[o72M`5BkJhHLn;lUKfTQ<`JI4lGaML7Z<eJb1JmRhWk9cAgA9XmAT<nnl
]SMJDRM52<l3>E^AL31ScjUZ;Nib0CZR0=EI\;G?4XAYJ0G^]4Bm=GBd`ZoI6=Da
]PIkqn3L44GL9^aFg2;48AQfM@MO;[8n^?QMl`B@`10YbO`VlU@nT<Yg<:]mQn@1
Z;HFnZn@MNX\N]oSLK`hYL0I=OSCXT8fl]9iCieKo0PnDZa`BBFEWHnZoZ`E6lJ^
0fA1QgXn7X5J33eO;E^_3LenaiMUbl8YG?b;K1MT?0_KMpXj2<2c7;iaTaTDOmm@
[@^de;^BNd?_TfTJ?Y53Yk@7H_h8JC@26W`WiemHEh@0S2GhN[Y<YGBfOPiiDm<C
HMoDV>MBNdVoUh_g]P0TJWSM6k4f79Ui3f5MA:;_JY`1S=aecYM20Rg@Z[H6Ro<O
Q9l\QlEj3:8a`5B^]O0nljqa8N5\lb[_gG:U;`]?0SaAEPgFVNI:cgG]42hkFHL9
UeJgKm3dG=Q]9lR0039BM1KF\UlMC92g=:YOkj^f\WSO>8gDV;eZ2W`07^\EoWFb
>7^@>F4YP]R:?Z?kESh6dIS0>ChX6booQbXRDc?f5MCEERXOB11:USG`C8bEA1Wq
?nD:F:mGQAg@d=[o:>[oIZ?>:b?S06<^kiLb?3a:P_`IMIJD]HIkZc6Zfko7:mZ9
Kj1CD081No?PVDKe2AIgN0EQEbBOg;jON1=B?>n5cX6OP][o4R6V6=>4TMRbkO@j
k@=P_J36KLN_01TV29FfDZadf2i@mI<\UIAa?kc?q]56`>S:NV=@]j>]4N4odGAd
YlNTl9dg_g3oGY1X7]75TTCQN2bmGQmOfJ?<R_5`@U6R5X7O;;9=KbIPC=?IFWIM
k>N;DW=^mMCfLLH@b584`d712FmQZ4JU\OV2A>`RiSil71AD6d=c9iKS9=UmSeAO
Ah2o\P5B9;iaILEedpM:3g_`UZ_OkT^C>fNO=Xeh@O`[7_dOKKa8nfjPV^ho?3iF
PmId[LNVSZoWGZj7Y@VQNN:4CTYL4;M]3HW8jn_IPg?[7_0dK2=I@8DRon1]lJ6Y
N\WeN<SPVjaf2ZYEfM^CNJRY>g3[h7MPoeWKPcBNlZj>4lmm<8GKdbD6K`pm=4f:
kc0J3S_kX8YQQ<B:dVFSBN53G1WF9EK?0:KOXP1JXN90=P9XFI8KA7hQd1c9FfP[
ieLdXF[R;YIlKQAg8n6<B=XMj0eaV<eh8QX3Bhl9AYU>CI\MhV<BjmZlBHi9AnWY
2HL`1nKG;``loDREXe\?P_NUUYjHg6;hJ`Bq>Vi:`ZfPl;R@f0bcd`feBO9A>@g3
Za]N0Kkj<N]FhBH4mJXfQ3W<H7oBOUhSl<]8A4LVl1<<2@hcaXLHbXM9=8SnO@e`
[Alalk1iI@nEJEg9jh2K8IOG;iF\A6TjS8d9S6MIb8i`Bog;6cUXbES@Qd0?jNd3
ZmX9gQe`IdHBpMTREREAkA6hlT]cD]=^]BnUh1A`3Q??P8TNn;GTPhXpRO9b<\1n
WFON4Vcb:YR2VeL7WO0i6Fo2I4icWZ<M\m_XMPal?_46IFA=SZ;Pl9k]Em]M;98@
;K>Vo9cT4HBQLl`R1Ofia]d@Z4a\LEh>PUdPJRX8D]?A\SY>=hQcFfC4?h@kca`I
m_?6^U6F4HB3JejE<1d>HcJZ:@8:Lfa]qCVQJe[9BL79B1LHQW^@lan?F:XLTK[A
LS^>f?<68NFUWeKE^H5D<;i]^DDGR84=I^>@nS1V7>GbV3`?mj3=j_9LcWXnVF8B
>HRljaWenc7MgN;TB_YGFS`2Kh<MhTEGUA_b62L4DaM\lRYjajbl4EHATogMeKbc
1G:[jaBoJph_X:1WmKBamJANAF]ML67dJYb@8hm]FJo7a>Hb0lGHhLh^Ca]7BC\H
?FT\C<88@m`XdJlka]Cn9OXZM=Jie6k<L`^@QD>UEQaReeK@YL2A2mEPPJ5UWC:X
0;b_V:]k=4kim1R[[iRPmX5X_XJj4S0dMEeiCX_C6eVad<Kj0=p\45YBNB6T6_`o
ZJM`KpFNAZ]MT6;?BHa305_m<iVR=>4@JId6:TgTW6ek8o=\;m<NaKm@[JV1PjXM
F]HS0df3_Q>Ik@Dm4?j>0>>lDn0`KGa@KYKn>NU?iS]\78=5a<;]F3b0Z=ZjDZ<]
\MXi]Ga8\2XAcR]6^>S3gb>bE;GRUD[O58d]c\nWP_]0dIpcln=Gih>S=?aj@7X2
2UkKEK=d@;GPW_feo;ZAE?WPOMmecN?7T`:>oFT8NPP_@CGE]HCUdmMZQkXPcOD@
Lm\;J]cE@@m\aXWePm9C]FJb\O[Pe;9W7T?@k>?Tag@8FEAi;=2=FhRF>G;;cXU@
d0Y2E8QJ7N?POV>:Yg<C2Z?p4AjA@5XA`?iJmHEhRcSG6hNg\2Q]c^e?ieIEKD=K
V>EI:2ZKJgm9S7Uh1oToSneS:DW<:O8Q]GKVgiY<LN>Ea:^OP<Qokaq6QVS_@=IZ
DCL95NF3SkYGN``^T?9fRX>XAYE2^3R80NdF66<lZ5X152GWJ`_;bWDCB9C`AdfU
\Lhj\9@idETM804mTb2JLCH`9b\g[Y7[i>h13;3=P^]Ri<^nG3Y3K;Z_MiUVkSfg
12i1hUlioc^9TaR639=n]dL8m;AgC99qc;SoBOkVGok]G<jLeTEbL5>3eD]kL4N1
18_fj7`Ui2HiBM5cT?V=XWQjBnd`If;GJmdnaHTNT\11EF32fX9>eD;D3DUjZOjk
`G\62Mn]YT1]l]S^OF;5D9K>nDKYP;CVKdM:Y`78=c5MW1RifUgLX5WocjhWnj51
[^l22T7HqlNmdGQ6=\@>=D=2PZHPGC4LZZZi3EY[6@4Mg8JoOB;W^oVX>6LnA6XR
:22;SSH=9V36R`gE`^S_8M2gaCeX?P>kFcZLicoV`HU]`;P=LiFPQb=LAngab\Hl
nSSh\AoN=eTKTi:NP:ek8<k_1C7g?M4EhbEcXT;099jc[;[k@qeNOMMg219:fJK_
VSTFKV4jA<S[>4;@cij7bO>e9hG[k3T8i0agB1;?gOgc1\5M;]hBWm_8mYY;;0]G
1O<dD5kb@7Z[mk2Sh]ZohRAeWgHbFCeahSoHWfjSFQAIoif7HVVocUki]<GTFJ8E
j]<?:3^ci_MUT\2A79jXFgAiSlp?]9[hCLb10<UW4?LROUTNT<9l3j3mnHMfWZR]
i?26Bh>@IEkk;mdUX7aAWoU2lH_Q3HI8UImT?AAiJb;VUH;mA=NS3E6emKP4eAb2
4Lhij?7L=JooZ>Mk:9hZTHG9IkJZn5d8EiaS9G\hGoWVX4IPT?Md5<1JHi9\kYd2
FFdpld1cfF_Bm=\`?kgNgElOi3V4LAEYX3`8\CPbN[O;QmkfoOSBO9P8TlQ8T[Qb
m>X1RBKB7>4fDdCnFVJ:H9Q1CO>@]AiEH=]Eg?AXHYQRH;8ThNElLmnVnf^0dZ3m
3dGW`fkmLMMoO\7P3<HLH8@ae8[TOB^^5C0hDmNLH>Tgq[AHQ<e0AnQgWOW[ki^^
bTJlPJ6kcW1_\3BqDHDBTngK?\_B9N:X@`0IEob0]O<OT?f4n;7bPSY>0_l:1:_`
bbJH8>WY:g_oGfMM_V?lN:<l\;_9Ul@D50kQf[DIkOkeZM5TKk=meDAKMTjmdlRa
1>2?<@iV0S?>E3<ZO69JRB>CVSg^5>bY5?OchoQ3cEB]h>OZH9^Ae]`XqK2WiHW;
Kl=OC=<ANdWaRSnjEG;3_elRN\:;Eh9U@C29P^\U^oJC<jBIOP>[ShY:ER=NKIGL
GPVM@GUU[:fC\Ya]Po;:K:>ZHJ8:JNhV3HLZ^JaTZkAQD[`6_[cQ=:KW@HS<klP0
n5jc0cUD_:`K_En\lEGmna]7DV_\DNh=dqj25Mc`fZk1o4VPg9LK0@;lATliL>QT
2Mc`gic>c`a:03ld2]?o?8`o]k:RjXE0VQGLdj3ed;go>COIZRP>0C6K7MgiP\hg
PV2HHH?5ojZgbUk5TGflD8@d]RkKH6e5Y`F<QEEFn3YNLHJZ<;P_X2E9\Vi@]dYB
M`X;dP?F`4p2hRh:hEohU\>7flk4WUiJ^Cfg_\Sl`QQfX30QKmXNX=8Q_f\M;ATb
ee_k7TmmTg`SKQ49ga^jd@^2]B\IARYaOJh?_J@8RBA0FOWISQ>JNS<H_YaV?3ZA
1^WNiFY`k5]SETC4G:^ce8d=Vl1I66aElTCCnh2kWkZ5fCFID1<q<;clj=nUeNB4
03eR4mcfW@jO`4a>TCjU6cI7Q?PfUJ@F:TDIW39aJXXLX6>NcncN4;EPg`5nk7m]
lCC_a;KC[>i\34a>W4nVliZa97h0i9eU79cN7P7FioCg_Dk`05EOYiT2akQ^5\\n
P`f:aEUPd@27^E7l;XOe>;CF9JZ;pJ5bRedSH\6[\8Tl\RT`Y6J6WZ7P^\Y;f_\G
U05`CgS50=@?<m1^<SZ:GaK;a`hEYbF3jg]`Z_OVTF_X4l^180HQ4b7Z<aIY@Yeb
@9l<X;?a0ZbD7IAYEkKT@E4<Ei6EOYdi63YBolLGJTS8=lGZoW7a0Jo_IA2;DOm>
699N3p`]1A1j]Xm:RlX>^MQ20oj[_ShF3FgmI0RnJU\j67\^MB9JGL3]ODcG5g`k
CoaT516jS\\1JJ10k[OFoNSA22VXDi8FLlFKGVbeBiSa`a8D7IkbGMc4E<ilJZQ>
DRRHn[7WS[5O9m2Adi_2S\Sh8a5[A5JLG6h]WOGS0@S]R@pmjkE2fRd2\cAZh93X
5h;ki`:i=J0lNXFF>JPSj_\N?d6lajMR8jSUkMMPj<E7[eEKBe:neaQ_2;ePTfZY
1>B5n8E2=SfCgDQk0Q5[6[J8b`mM43GEH1<dnELQBW[XKP`_KPnoCR=JGGABPI3Y
EI8fhoRg<UW:do]I]I7[2Lhq\eUakXWYcBW:k0UUJVnnJT\<0SSS]^K]V7L6qH\a
H8lAT7OU7jX[AcMI\1hZPXTPZ@B<V93Mlb4;RMVDQ6J5;2bb3COcD8XYF\hGo^S3
UV=XOlc@<:2QE@E8WaG`?IT25nin;iNE7QeZfg1bgeigfoU@:BSK@b][Tf_MZSVP
AoAMe?iSGK@jH@2_3Qf:RnWdXO2dS92]RQh;3qYd:njCm`80X9>Tg=o`]:ScKTd\
SVV0PNVeaTLV`PbX<=SBd=j6oBlR]n<>a`Y\X0I:NaIH<ePQ[@l:>GJJA:Bn`8A\
]?KkM;Dc_YfSf9>?U06Z4Ma:I4Q7TgeZVJa2C`=H0K?PTNhk:_R?YRJd:OncM>jW
_lf1fNKOKVf>GIq=Q2\iFQ8_GG;R0PeBDjOBI8Da]61V>aj9[aYTXYFKGjA@3gI`
BVPlS@bGVISd[BDe?H:TWUQ9?hYmV<a3i2C10EFXO4^RmpE26V=2f4EBRQN@3=6^
n6gm:;5cMm6co9R77Q=?iQa@[EQJBQH^^51GlDdAY8ecg=9Jc^]1N>3W<_C9P?2`
REmadbaeD@BeETbY7NoE=0a016L;_BcCko0elID>_^6cNFAjE4XWlJpQ[4Zf?SWS
f7a:dV[1HT2ibB3S=NgO?Z=Voc4[b6__S4;>8N<B>^YOg^A<HXcaETd0=o[ZZOi;
WBK^@LFZf7TEJ1aZBFJ[@YI8lcSAlcS_Gf;0Y=G\FPID5^li0S0LJI:7=:D\I>Wp
bo54CX\b2Wk1IG23_a^Ynk@2^5EDcGVPcCW:VCgked6ZfJgf_oEniaFQLLRgoo;k
FKERR3f9fhocDZi30lek<ThSQ?=]oKSM?7W;>o:0e:k98EE]gBjo>\jDhhZLD^G^
8nFNYa:4qk\Fae5m?`P\<KE`c5H`Q`AdSYok?<hRei8?U\UT?k7:8ih5n9G^:BDL
1CXaFb0_>=E\lc0c6aUc7;dNGJ2T`i^AVQllk6=nX:c?W_ng7\1Pd`]8P?LElC0L
L`d5AWF[BHU5d8Tc\poLcCaE6d0cS_E=A5Ed=[IV=FUecX6_@HLc[LfS0<GgWGT?
RgQkHPmcc\E5TQT?=WoSHJdARafRkao9gXKNQ\jlMSlLDME0hh?k[7@OWBGPWX>[
<LVQHV9<@Z`RRnVIcC7^RYF7MTpQZhg5ma7_9fFl3=J?>W9QVD?]Z0M>fOZ@on0=
[SN1JY5j1?[@K=N_`:FFBHq`6fOUY1:\AGG9[kQRZ`lQOUGR5K4I]K_55hY8RWZS
a9?jcT2JfUl;iD:5L3DVhS1L3lBCk0a2]:7GgBXjSNea]kJblDH=hJPX4hPRRW?f
b30Kk[=e[naH<DlDiobE2MKdm]_Sl12p6D>FM];W7h<@@7:ZYZTc`S1J@DR3\PfT
4`Ee;?aYm[hCXVJ:Co40]1jg\hVcf^\8[NfNMjCBXB6iBo]AHN9aHHg1^Y9;]_HE
S<E;K4\Fm6`?R>iiT;2ZgPa:42e7Y6o5mRHQElm]qYGL=cJ;\nA]\fbFKG3G1bj?
Tclh;PMEUg=?Ehe<JKRQNZJK;QHAiA08\oUkX?lkfSVUbXm37:e<jlD=\7\Y^DX0
H^bA]\>Yhd`?Nn:jGmV1>M>0I4`j5f2FjM>]KZkB8<OO6J_IKq]lGd\dfSN:EXmA
[mb9caig@>;`QHf__l6M=XM81eDg7\e=R5_DDkKQG1YUNnfnG[Vg0icU?<LmZ1^A
7?IES:38cCf2nMpU^J>:e<FQ]QR3lV6EmdEY2`j@F`S8[>[nO<YOCDh2ehYbo?0g
>9>J9LMRA=C`=U:P@@8=12\J7k`g7QOKXmCPLQ[1?hB7GM5;l<65ImB2DZk=Uh\A
m7Q6<LRM4:VhN?Z99YinnJEq9SN1mkaO\KgZ3`hIQW=W9FlD83NIhVJ5@\lbTB:o
HbGkAQBFma>m]0meelFJQ7Z2^GX`H@RXK5@>`WS>`E5ITd5PHR_jgl2OQ^lXG0J_
_[P0HX>_Chm\mFg;X0fIJX0V>Fd883QZpg<WmYJ8lCM`g5hIK8bMDjhaAkhK?cPm
o?9246G=[2c20j1:9UX6F7PYk@7aUgG`I@<KP`OdHDSLDFoY?d`k<2a@mGY<7J6g
5GH2;Z>P12K[OLGak@RN[JbYPY?g8_YjkIFZATS>gq_>]:DOV9Wo6DKAeAb6];=4
IEW=VMB]0T51:5n2[;VRFnLCp2`U=k]\\8dMEOL@^VdVk:?MbW^8\VO@LEK9HCMO
AoCVB;lG;hkD=E4cYPYmOZeU5\YNUZ5WlBNQ7ILJHDe9RhO8cjW=oN^89<^90B:C
go3j46SDNJl5ikb73WBK[3PmMcDXo=RYNqc77NAe?_3Y2kS9H9T[N1l[KY;]`YNA
9FmAALbIEa6JVJb0H]3j<9[N8IIRkh1Mn\X@WNC^[BA7lKCB==<\JAjCCkPj\n77
SMJEA>jmR76_[Jf=HFKmoU]RWdB[758;ZXZeRX=`[7plk6PkJcZD>O4[RZ;d8Z[S
jnkX9\24XYjH<]maA3kjiGaXRXM1^P^Xm_8TLjleZ1A=bkBUgOh^MD5AT5N[FOWm
PLjlm7Gb_UbJN]bf2kUATmT=jO2mK8LGj_8OF4?T<l>FO80K@kPpEk70[Qh;d`e:
T>0iL?oFKMN@;kfSF6MHm]5K1Sn^^JY_Sf]`0Da<D9o`C>C2U^^I=O`nPZL_T5R1
4<FT9GU32eWn1eDWbbT93456]h<JV1TjYTUh2=@3T?oXOl6?nD_Q_@GojRCTqm[<
5nkZiZ7j@jFfQ@kSU\AR]dYc;AhmY2OTGa@c:60;dJCn4=k0;dk_6lM12;o7p=8_
OCA03hC]4]UjfT]UP@QW0Xfa?G7EfEg>;KWZ7b=ZiIS=R0_emFLfIK@\oYYJYNgo
bUCGO8T@;k3\41KUNfPfWNPf6oi`oi2>i0M?;5R5dRLV^Ocd2KcEgAJ@=Z^Na53L
h<lSep?PEXNK_NSE>_?KKa8S]<kTk0P_o979Bk\53Uki6n<`IEmkb>K\Tf]]O5AI
=h=bK3FJEP[jTFWBIoPN[32aVmCQP8LH4ZpbVOQDREnDihI7iaHC@[<5;:9@Hfb4
nI6WHb?_hA<YgMeJ34X6QNc<T;J48JW_K>7<G7d@D?L0eb@nPdi[[nA9EE^H;V2b
`nlQ<boW1`cfokP=h@YMAGnE;;=1TNZLD`5cG:iIY]DpTIRfE>B^>ZRIMc3_9?E;
@ZX=B]LEdRWVVGbHhgmO]HZ:>6@Q3^<:YRlnj;6A<g`D8E4a:ZigSeP=gWoWGDA>
0SlXC2fFj3_Zj]b?[D`;Il>PSo>g\\GQmbCPU@OF7EMjK2l\A2kmpdVJ`:4H_4MX
<=]\=WmS:4S^V13HQ?4m;APX0fW9Ul4KK7_6X7f7SDkA]kgLI[EGPHbLZCKf0CHm
VAUVEVjII<P7RaQGh^ikN[BXi2<6cN\34B]ASZ^W71TADSWUZc`?V\?<0GmaHq?B
hc;]W\c9N?e\f45L:eL@fPRnEm5HFXDOD`3D=@;Z2k0?pdkfh^ICdd=NTh0hkbPY
5hJi?@lFf8dUn2dJJ<<I1n@g0A3HRLW^nW=b1gfZMBM?;FnO@HLGQ@FNlc7e>RCg
2cPF=RDW4_dJLHkJ^[a3Dge3MmZE^g<Xgf4Eeik2:S3@lCPG1OQ;ep]j@__>oB>0
kA>n=2030gINn8LA@RSN[P=]MiJIZ5^50;bIFb]LoM@cNkk>OL6o;RQkE>>NTX3c
4[;EZKAV;75;=jHXfR0o1SC=MY:RoaWHE:E1Z>[om]H0<2QH_1<_G3]YdSBZ2Wq:
6@0nn9DlImZjg>aIP8[FRQhc>AW7aCP<WmYN4mJ?I]A_ToISIoXMEQG@>:Xm5Fnk
h]V[hJh9;\:?TldoOHnSL?\V6@SGTNIMCmf^Pl_HBCUGP1Wfe7@E2QYaf3V>dK2b
Bg[CfPEqIbX:7Gi^aj7a80EXC=@F_nZ3TJ4;RiRV?]Vnf;N;`OBoJfjh@am>IbeO
UB>hLM[>GQYgNLBiOC2Xjh=l2[EAR`W?Gg2A4=\RiKVnh8=;mX7_EO<nlhbln8ed
R_>nlUCIB^?KiOeIpW9i^`M6V8cijoMRf2a@Hm@2<WkV2CJKAYDL=K4QI3m6CqFS
F6ZEYEf3_P3M>JFL9=ig\4cViV_C9CnYWYLUF:\I<XZ@0FTX_i@Q_a2<JajmHaRh
c;ISAO79dWEnaAV_8c5[MPTCN1G:6lT6W9K`Ki1X6NRlQQMmC7UARW`cKQGgAF]@
TE>@8aq[cPPGXdR9c17f53>n8OQ_8ka5MYD:EgoIU:Im0oaPKGCfo:UWd\UH8P>j
31lKk24S`M^=WBY1k1Ye=g6SW;OPQJ@V7N;qSdCgcTqUPcDl_B$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUXB2(O, S, A, B, EB);
   reg flag; // Notifier flag
   input A, B, S, EB;
   output O;

//Function Block
`protected
:UI^XSQH5DT^<TFH;]g4c`e7k[gCAh0^U7`qIL36d2O]?5WZ_cfk6bC3U`9ahMj\
XhL^BR`aY>71H=iN@alUAGA8j@`SMF>XVOQ\EhZ[0ApTjBYf=iCnKnG[XM=cW0gk
[mWq]bLOD=qZA3_<nC@=n=U3N3c^loYnR_nigIH6bhMAH^2hfCl^lma`e:qidMhd
M@T8dRV4[>Sma<d5_NDTRZZqanT^?VcBEAR\ol9Qnhh27]YqLTTXBG`5DZj`Tfme
=S]A23VNEU^W:TmF;`q4H7S[JnpEa9jk3p^RcB:HbSB363I92B0Vol[aM48XK=:F
6FG3hRNdL6=Va21RTE>SIp6AI\oBn>jS4N4Idl:JNbf1:>j=[S<FTc?KiMTFNjin
[E[EM?6LJo=F6Z6I]Ga<Li6`458^72f_gGi]<h^3@G0P0o=SADg1T_OhWph8SG:_
DQcAE7Dh4BROI33<Ub@_;iKOkkaQ?Gl3gFX:D1V_U`<JWSO5VCneCf;UdmhHDU8j
ULTF^5=_`=Ac`OUP`^TiIP]dk[jcCpa80lYMLS`5anY4M]a8UeaIc<GOVakeeocj
fH^\YT`9h5GS8EEJh[?PRH[DFYF3MMa]G9ndUmX4Kl3bom>JZmpPQ:3DfRl4AcNX
`[]IohF6fKM6TTe\04]XKTLOUahjXC;46okS6nFFd7EbYFm<g<fP?IBoh7cOakWV
_o<7HVjhbLSUH7>F;Z;2NAjSKSYWO]>Wg_556q?59^`\Q_G4mH;ABOMVG7MGKVGn
MAjOO5nkTV>o=e7`i?_DN:J1hFfWF0]]HEmT0;?\B[UgH>h>2jJTOP@n^9:Hn]6n
lUK^0kIdXJLK^61C95=B88haq>2AH9KgA=ihUWOSE5A8H\cf27Vbh73EUiKn_HiJ
=WYC>7<R]eWo1;I_I4XHWYHMC>?Ka7=Ac17EZjX:cn@[`pj3^>V]HR;kXQP]HORZ
>\eGAOU]FVAZSNQK[;f]]D[lgWALJlMR0XUBM?nMX7m:DbjhRAfj_H7TNIAA4ll\
>Nm>KE8RW[Z]SZ=d2MNXcVO\UH>Lji5cK6TLcQlXUcP:30S1po<]H`cXTI8Fok52
??A?N\kJd`B5DDSZ<TcGEfOWjca;hUYVefBgW>ASKgWJhZ>b\o3Z88Abb7J5T7lc
J3^?2RN9ZR@>nXiZF8o124<7Sg7;c76`QaOOE\X7Pec:NY>Oo`kq:[`>m[2V6J:;
>1MJ[0EebE^HLi3He3PH>nqMeHDk@F[n?kbXjl]gKZ?cWFod5[S=3AHdG=1Oi;g`
^gfbOioBMPMOA\l0ETafXJYM3n\iT?12H\9gc8]YmZ?oTh4kba6E?A4NcITUkI8U
fS8h<hU>J^XZATnD_\2jXKmSKqD4R_542[dFCCGCFO9EN:ilB6I63QUng5FM_5Pg
PZ6[lW8NS:jH_FZoA>P6k857j0Dc7WVHUK>=HR7fSPWAjZVX8enFf67og\dVTkUd
EUgRNf9l9SQKOb;lBYVW9c:7`A4Aq`4[6<0f:bDa2HW;?[fK9N9L5_oB0>idook5
5Nc3O8W9IQA7]2\MSXF2MIo1OcDf@`VJcDDUMI_W5KTK`Q_HmNEq:Qd^gVQ6m5TO
Fg5D;2K`[OZD9YA]9h`[TAS3HPUKb0P:YH9@P:SFfah2e^1C8HV0:e8R@h\M\BPD
A1`5eYFh:lo7Jj`Fa^`UDYGqX8>I<jhoWCRDloS3fod_`g>02cI>4MCeSGnoRg=X
JNJP6P?S]:<\7DkR^[E26NeZX9N6@GV68h5Pn@G<o\<3W4oI^l7<h=Ce\=7plHnA
kVQ7269:]okfML6Ad6:<mHP?g;`aeXFSO:Eh6G`H^30qMZ@kEkIPeSQYgUI\TIT0
eLFUa00hm1QWY=Rl[IAn3Ue1Y@0ggg56_fUoTgYFiKmOMcONJbY3Ia?]6g7_cFf8
pN>Wc:DqPUWEfg`$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUXB2P(O, S, A, B, EB);
   reg flag; // Notifier flag
   input A, B, S, EB;
   output O;

//Function Block
`protected
[;R@9SQH5DT^<FXYcLNbSQUGMh=PeG=:C>cfNd<]X\i??d5Ip=42VTM1a^TO?GMp
;@^\JFXU1cUg0:ZI[e[b<lFlpCdjaKQp4hOCM?:95k\ioHgA6\8kVR?iD^_E=Dc@
@_>1o9DNPblLgfPqnnbja]@T`jM:f75bPl4WoK>B@93Yqg0l\W>ZlH5M:nhI[E>]
5eUZe;b\dJkYQ3=qdnim:cEpF=XUa1p?YZLMeGNd4mc;UmWEPDC;A\D`Bn4\6?fX
EHOKf\K6FIZKiXcX5lE5kBT;9T6ACF7\hcJP\H^Y:DaLLEKQb`RFl^J50?_[dQKL
BHMX3;pcV?8c22]d3_NDY8Sh8f7^F1lf1<egaQQjWkETYe8ch55LVT]XZ5o9V_AH
RJQ0jB1IR^nlKm;GMN3OddJ?:l`\F\HDE>[O4Z\1`k:;^;qEegHVJ`QYenQ\S2[C
Sbc0W70Qk[iJ`jg6dMh5G875ILlcEGG_3SW[G2@0D7HplEE1n2K0>_dQJV=ZBafZ
hnI:DS<edQZoOIcQZUl3g1OM>E4]OG60K?6;UFiEI:nQJnk_m84OPF@>cZ:HoJHc
@IQTq3@H<C=LLOZf@XHHWLK]Z>LPio@dG>lA]bNYLRgH[NARcJ7O<4_Y\TLoQ@j?
U<GK9?:iT@J`5WG28]\OEdI:G;L<mALXTACQI;?YlVF7N1hAf:olE2\G6K@D9C@q
L82eU>hP`;n=N?LkGIR11giVE;RQkfVWLDThVg\7W?82jdlLQ?Ak]gEUhAPod@BS
\<SA_9h;h7RNFVVeM;<ONgMVUAlCS<_^4L:8Qlc9\e^V<L:935j7;gpKCU`k3:hk
kffCT>W4R=nbWHUe<0nH6NODUT_c3S1j>7B1;7Xa_XI<54J;jF:\jn7QHe;Wf;9e
Hla6il?Fn@nOc2@q\2@eVFJb8\FhR9@Td=DhUQ^iL\cEK;lDA1JEMCm_\m<EDlh1
?G1=niR4:9<aeKKn\U`VHU0o6Afi>JaGBkDRWjDG3CnRmAlZn029O5WJ`[l=Bc8?
b6?`_?5B0_lL\KGd:Bqod@WbLf\:TVH=UhUJlKbCkDkhBT?>;>DP5nJJjbaROn7D
n72=bLd8]J4k18C5Ti\o<Z8JB<m<oBnac>h[FKHg4Li3;b[UK>jY?]AAfPVL[2O7
eYmS?1QMO]UVLC2\TU3e]pWW24>7BHGhAcoO;636b1k^XhIHSkL@C@7?::7lS<1Z
\eaYSFf1<`gbB]QKAogm^QWi8jf>_]1Ah5G^1g=@b9Hbi^G__2>jCgkJF6@YY_HE
CO08G5\;dNlK\0nT[=Tm7R3jp0N?Q3i5V`HbKhNSi;Ep_i=[:1i_QkFGhE0XQSg9
C_Tfa5DNUZGNCIY9[7SUf2iRQjeWaBASTKm6\VG>6jb;_<g1S;kKF<Uc2iM=:Wj:
0>S9^IAXIeGBa1ISdlgg^e85<WWTCmZlBc^nLEklSj\;O>q7dgXO;O^@9e^GU1=A
6CiCY2f@6`:o=@0j4DMbk?h1LmTcBNMbEoCgWL@nF5TOe=>7l?jElPRDGBgS7TB`
S:TF>pcC@oZWMg1:;@BiO@`fdC:TKH7WnjRT8;LZdR38F`>FC<\`^9SkW@f@<3Xi
j4Yg=aHK4?d;JXGM?PoJ:Tkm:Mf95CgBZFiUdC;kdHNc8pAoJS>ek44^c0jIeZa]
PB5lX1ni<<F^Kqn6NFMOiX7I57>E4]<16RYE<EaKj_RIWDU1X:7<BOCXc=JV=ZTX
fcKcb^XfAe[TZU8QQj09chH34QQ2acd6Cj`E6E`JKh=mC0lNX[<RUqZZDU=E[=[g
4b?WlNV>X6^A@U^cJY@Ghm?D:::]`hlCER6<A6g<g=oO]Lm>Hmn0bnhOfoh`dKNh
T;XMK@<P5dABRfpFTPL2WpVoahU5QMAHCHZX;f5b7?oM1q>?AdfmX$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUXB2S(O, S, A, B, EB);
   reg flag; // Notifier flag
   input A, B, S, EB;
   output O;

//Function Block
`protected
7]UoHSQ:5DT^<7_:[iKF131OCIG_1c>>:XKc[]@fdRZ4054aS^1]Zjo4GBJY9opN
7ISTgCWN0E5Zf<^hIG;YX\PXi9nlYR?SC4QOO23a1lqOY;0Yn=H6H1nOcR<=h2YT
nWOVWTdP>b^9EZYEGME`ZJPO:`K;XpfJeG?>p6BN<>G]hhL;n6klc@7:DSW[MHA9
bc_k:NcnFkQEjha3M:M0qOCOgRF\Hg@VAeV>gk12\\;iD=@?mq<QiEY^7?Q:nCcG
LAeN2LceAf8H_8iikKocSlXgUJ[BA3H>]6;eTf2N<opGF=5]V;5aB^91R9XBA73A
T>kNHC11YgkN=pL;[SibgplXg`2dpAW\hR]XIPQcAJCl_cJSJ2EEgj53Q9fZQQNA
;NH`03^4Ii;bbgbXW7gDZQZlnJCS^Ak1_o^f`lh@V>gRENiRYbNX35kL\inZNC<C
p1m_]W?Y7R8M_NOH^Rh7aMjWFRelkHC^Kh^IF<@o:DDU?086dJhcUZX18JI[n6ZL
31gXN]j\5n_K:Fj202UaIWd4XfVC=hL^NI`0qM_AF@85=lRT=D=9BjBRX\c4>g11
65j=EXhAJEaV\4J\E_N3hpLfShLQ_gZ8i>E^GdbY@7h:L7P;k9>acengW9H_URI\
50g5CnLUoJL@2jaAomLnA:L7Q@3XLE>@n^=>VomdATqFG=caRN7_fDZUMQ[mKUak
TQk19e1_7Rc;<dKQaIMfMWj@EkW<8Uh7m:j`69dG@9NFKEd?6Q14OZm3dEF<KJ^S
EjJjC<a]Rj>5fj<OCoC2kQA]XWUm2qRED\kn:U=20W4WC08nT\M4_nV\EGQ>aQ?5
61kH@EW5J:n>B3<@G>d:8Q:5o1?hhWRUM8LKMh3hG2QH<]1D`EZkNWGnUJZ`BkhS
Kk6APDcmHIh6<oW8pLnQ78?66Q`V>k>K:iagaGNl@NnWm\l3KVm3V7fCEFClgjW5
KeVNYFFICFIEQ_DU7LDI_jeAe^6[J>TVdCf8?q1UfgJ5LGU<5Ue6[cHSY6UY6=NO
YTkfPHiia^>VD\1;15Fg4`SnFLf93?=QJ_4BgX19bPLZ\BN3CX\AgUD[iD\@4`1S
XdJmPf:OSV]CJ=bEEeo<Ie>F=>;?TMQ2=;MBMK7kpcR^j19@GjKULX7`lfjK6IV<
mZ\EZg9\A<42E?MXNBQ<dDUHgHAW\i`bg[hJZ9938cn=M26[24YgBSbh2^6H5@m4
eJ37HDM\`AP=7BmNe[=^VKLmN?iQCY<o2SI;Y@9[Lk_pC7Q6dL0<9XMI?X89Ojl;
>60]WRKOYm5ZFg_GN?T22:O=SR3h6QDS]gJIBHEI^2hRCC^hCkK6`GCD<12;KAcI
:OOC9i1O1m5_HVgm`kR>Eik@DmK[0g3H@JUOR8Z0P2LhJWqJng\XBZNFMaHOFJ8d
<MVY9Hha[X6<5TC17JYYUM0gUYfmg9?fXLCi`b[Hd2ib`VJJG7XNWIoH=C0jl;8A
eAP2n8CJ:GXLcTHOF0<?O<J6;MTZ>k>jH@`J0Mob[HHb`jQG<qaiL6HSdnj[D]9?
9b8hH;>i@n6J582\DpGoiG?`F6[o=O=I[l6V18olOb3=nonV]^E=;bM;AEBiO@?\
dS\0=S6FoBiWm]8O>`GHmLo2hlKIS5BB9]G]V1P6qP2T_Q_Uji^iPM4e?OUCV?C8
>4SQ6lkBCGSNMAij4bcTH`W?A8Tib2eR5`ZO1oA1VP5<^4f;lQ@mU;IC2;W3>\V3
QAgBQ2SB@G2`pnDGIR5X`<aTVQYfSaOKXdHe\kRg;Y:]g3VE5eFCC=]G7nUd3i5h
\Cm`J\^gGd>EKn2:aM^\=Oeoo@55Tj2Pk9FDiH6EJc3]Z\fWq4fASa[M`omDO6og
6MR0;RFhN^l9KS=FegnlaH3A4@E?lg`ciVDFfk_fJM?W>\G@A4m5?X^YXcZ47N2B
n9HdGp^>T6D=pUDgGm9Q$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUXB2T(O, S, A, B, EB);
   reg flag; // Notifier flag
   input A, B, S, EB;
   output O;

//Function Block
`protected
c]NP_SQV5DT^<k]R=WVmWhkR@0_nmh`F4\^_kB0aJ[^6jSLRe9caB0WmR3iYUGQ_
NhhPiD0E_87ap5\48:]IobNCUabAh962Z`EH;A819\hGYe@H=6o[Xk24<UVh5=aF
[0A^SO2KnWiB8`]dSnYp\BG9<Mjeh7ICMc<qlV[?B`p3:@fV4\hjfSGIIN2<[Ec9
lV9WZSmbQj4o<9[j5SDUEWfQoYqV9?\UgZ4?CLPPD]F^J=_ZJh;Dl_`qGmDW<>Rb
`hIYiD\0[Z=]NPkWA\?_b46D8jqe`CFVFIpR>gHeBp1D;9Hl1F08mELW<eZ<hc6X
C4Q8<5eOb1fn:DlnC73Tfi3JUH;?BkJYTfdJMIR7D0D9Z^=ZI@N2_XN9TTnF0W6@
EDWL_?J0P[N5<n]9JUC?=p`^cWbUN246@:4FBXXD8g=QBPO>QkPk<GFR^BBElWCl
d<bNoRMoM1_P9R;j[C7[`:iZ5heGSYogWU0[KJlX?WU@GHI;ljef9K9LZ\:jScR\
QpHJdeWNT7Ih6GKA0aiZeH@^<A\9jKn?0Dj9TiCaQRP:6HDfR9nF3c?UG`HQ>Iqc
Hfi]F=Y_ZDHB08HnSTTVI=65\DYTed@9oe81^1hZ^?cWm^WDKcJH:;7\PkREc@:[
2iUJC;FibJ7@?VaMEnX`=fQD@hOqh[US4VUYRZdHb]ec5kLjhUoZV1YT`?I^17eS
e82Q0IAXMeDleP:3;b0ajEZbKI4<OMkCAl^>SWF8dAI@j^F05kK;9@baUObRDjeS
TAD^0o]QGV?190Q3>TIlT2pAjVG:eLYg4OaoOLhICb5]3fhI[1RT0RX>D?2BiY8_
hSmS1IR\0PJXkY]8`TXba`aKA[V\MVRKa;c6`V86_4<:3j;NIQZij9:G>J02Ve\D
?MM7jSHRJgP9QpKG<cPg11oS_4FP<RZ5>>1S?YWGGleY:2QNUUE=_d@h>GDLBdo@
DoI@J9[Ri1Og2WhnFV@D2c2T<2<Ll3YNl]PUN^qbb=R]JP813>6f6eTlTZ>bY[j<
mbo35\@eDCb><h\gTmO[_ma^4H7l>kb9VLMDlNdbk@?lg4G]>HlDjd^CMZ]bfb1D
ID9VY\0ebg\>^^jmJilaDSd@OD3;J@8EG?4>l@Tbcp42l9I8g6@94Eln=CWMiY0Y
GakgXEOTC=_D]JChR0;WnTkjZ4SBOk5@0l\1SnaLWh>8IKdCp`mUgKP``h5k0hZb
em8U4h7ZB=i=5JENHm9`4>9F<6QB=?O]CZYH`Im7]mKAfjVOa`]VFFN>`WSX08:<
eL7U:^ejk\3<FDAN^:`EJXo^CHc<>G^WZ;8AgM<O0[DGMeVIT71p=R0dW`3dT8ME
UXTg<j2n@^WHAVBgPWEX;SC6@Z6bBDNKVL`QjNGQ=;BZV9D3SN>O=\^A4Zdm5?WZ
bLbMH\2b]\DY?PY=J5EJ^I?F1CYL9oYD[]4<l`M:S33Q6JoXON]jOlqfaZ6l;_JF
C`PTA_H@0_WPZV7:=;FejA0h8P=Ko`aVGA\:f==mCIn`GccORe0k05afeI5e:0MB
1;dd=32A^Liof0S3N_9PTATNE@cL?L2:5iP<VD7?Ch>SMhmZAL=<0XoMkp=49fWQ
SJ?egaF>JNeZ\@PULIHf3g:oW_O\@h;Qc6hn^Jm0U`V1N@m:lL4CBAdLFm=j6]IM
W^]laHZXUHW^V_]1q6@iG8f8hg38m>]^L`gK:CBmkXLYHV69[KQCG>dnm5eVXaUS
6B<3fAM6WdD6R?b`IUhJHZ]ckoJCVGe51j]iA8Sb>@e]FAl3mY1b2KZTQkk_pPV=
bF:bb;VMdW<4gU2DBUi:2Ub?h:3Y:Ln0gn:bQLbn7b]MEaQa]^;\J>bd_Ob\DXXe
;1d6QXocn2B\]b^4GXH<]LQJj8Sl@F0V]J[IgVUOqmi8BQ]9JZ\cXecGTNnOV1[i
iPbgG1;N3CnU_Dj>hmcO;2H3L:80J28L[JL6nEN[>^og3SWlj6C>jEeA04aB7deN
g`@M[pPC?j64p<8BTc5S$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUXB4(O, S0, S1, A, B, C, D, EB);
   reg flag; // Notifier flag
   output O;
   input S0, S1, A, B, C, D, EB;

//Function Block
`protected
B7i@HSQ:5DT^<9FRATjd17dIB581[=p1FaVOb]\?55]j[E@bdoW;;hBR3]5E]=GZ
IGd27hJi4Woem@kJIao0RpQTa8AECD`OS_n]OBW]eOmW=e5JDnSKg0l]Vc?2d6B?
moUn79pZhA6XjpA7468P<Ej[@=b0dQ6Phk3dVTR@fP^T8dgeL3@TJaa4T5]5SU;i
EckB37OQbQ8?QGfOpf^;[UDdGeH>b^IM:VcGm7A5LRmq5X?Y3E0]Y<gUjTacWbO=
6MA@bIJTB\bqYjhn``OpB<A[`Wq4=cOT2OcP[S_:3WeJ:k>U_X;`Wn[>=6PS?eA2
h46;Ud=of^3Ni5h2Wk=]aoNJ4[WSBKH@Y9iGC[2Za>\_cZEIEKN]7\9cAe<`eejC
i`O2Ne2M8N?B:<9miTAP2?650Nd;aH>MQ3EpcGnmoO5M^jKYG]<Q5SKIXmbGR3Ok
Zjca^DGIFA>Oq9V`lCa50WCW[ljOHG1K5i\fRg[ha5XOZiS_bXQah2h`LU9^`RVe
[XWbXeDUMd]kNYhMAVBi8jT>3\Ib?1@<5l4f;m5@4`n\l1E_HRFcMMFYB:Xh39@?
:9eb;=W2E8oV[L9CinLb9q3>`Jeo\Zd6_:bXcR;D[[SST`nnZ6m3^A90LAFdkKT0
9RWo?X@9;c^:F\02JS:i4Dn8B?eYUfZP\DoIh]FXA94O=VNE2=kAc>ScLFI`;edT
l:3gdg:6RZ5LomN1cF0^D3fR<8loaapZ6QmbLO`mP]8_6QPT6?mK^cRQ68S;Z1mf
Tf]X6HbF;@k?FTf5P[E<]X4WECVGb]N^L\ii]Mk[RB@ih9XH<>hJUb]?I4=?n^Zf
Hf2FlR><_j0HTI8O3[]\Tb2\=DGWM3cQ?0;NCn]q311O8Zh]NMj^CMZI;jRhbaEA
[4hlhhR\dHAjaIbO>SclM]2o6cHfNaFWd\3KVoEVqI]bc3X6InA<mW3]^TgWQUNB
_Pk?7>Za2;8S_WoTDfHV63HPCEi9n]<^hnkNNUUWYTa`nL<7lm3MW`ZfI7PLoUgQ
>YN;D@nMgFiS<7H=6lnf@lRRK>cWL9L^@j^2Sj4NVA=oXLPI;q75:WLEbf\eDW4T
OjIdJPXY4\0\a`Qe?Fl<VJS8Jo97D^CjX^@GM:K5h?GXTCM@BLo93jHQ2<DiOige
5]3SU_GZ]l:X]g^f_cCSV\QoA`9?i:@KUCT@27@Qh:KnW;D>cETi_=Ba36pCZ=Mi
fJ2iDFEkjLamb_KZ4Z3iGd>K4:6Zm79Q7gGfEX]61\\Ye\@\7<OnUG0Go`JX<o4[
0b>ShN^\][EPO20aZFe[65\N<C]=o7aC;Ag@IjmhP14llS2Wa:eRQ9_=A1=_Y;Lo
?69pPk<^EFEAlIlGP^aNodHPE;9fFifN1m^W4l4HNjEPWAK\RL7XGdQ?il=ZiGlL
Xb\?dD_fRb:[XElhOkoj;ZY^>VI7GQ^S2o4Y4[4Lico@J^Y>1:DhaMWnaJ=>7XFG
CeTNEGIc??TRq4Xhik[h8kL6B35\AQa1J=aMGS>9EP]?Y`;PA>g_S15=efD@\hH;
\HX?3dcSCCo:QDoJL6FJcD:fZjEdD@\nEiD9>M5A[pnDGIR8j4<9TLQYA7?Oh<dH
e\Khg41:]?3Vc56F4Q=]G7OPd?o5h0CX5;\2gZd>EKn2:aM^\=OmFh97DP\L_<^=
hQ<ER:cI]Zi[?QT;e\D]d`SnTQ;nj=<L;6Q8hgcaNVG]iTl^1]OU3iO6Q\>J?AUi
8kWjVjcXhMpD:@nDOb4GlRTYQch?E@GUI70RWSH?L\2LRQZETlZoIElp1JLfEAfS
fA?lK8fAAn\]L<?jZN>jlAI<M>ZH7;JjW8GZNmb=UOP1HO[14`PBVHE31Rh=JZ8S
2kkP2NUM^2k8^AY<kF5<XGIiaXk5Y?7J]`a;K[GC_:KGMNJ=]FF8M04BOBEcC2dG
2GU=i]gZ<]nAJ0[>YXOXXI;Eqn[O>B8]d^I=Db@QGc4oRS_FbN8iMC82oaKIHWAC
QT9N:9W6mF`Z?=]2N8A]M1=T;n@I1E6YMgfe42U1eAHmE=i0cVjQV4b2SS7dhmom
_SDIFc`XRE3O34728`cP8mn2U]?HCLV8Lg[AFnAFSih\jTlfF1l1j4G=2qi]7mW=
i3X9=G<Ef0fI7>o6]S0C:`SmUE98go5n\]L<?j6;>alAVEaOSQ[^]E<7JJi^eP=c
EO:OfM]N0Ne04]OBEcC[d:2GU=iogh<]nAG_n3OXk0aRIFo`IZYk^GXVQP[[\U7l
=V:;d74R74M]YkF?ZQRZa[2[K=p5TE\dFnH:?c`H8161QSVklp3O3_H[GbW;6MMA
=d@gmdHE<WN\mKAS[IKDkcKI]BUc>f3_[nQ<BkeFBc63bIlJ[V3L==6g_cmQY5dk
ISe^=Bo`O9:4ERJC[81KUUX?G6NB@mYd>X5aGG;2lCJ:`2dXiRUOl6glQdmRne6M
PFbV>Ghb_f\SWVJI9?p2OF1Ek5LOHSImUDU_Ph]na][=D>0o9?BEa4H9RmVnYNA2
P9[V[22>LGc>:Tmg=Kg2fh329Kl8EKD59VObZjF@GWFjQO@eU?^0B1h\6SIR?0Z`
GM@Z3RRnnU:e0;gD\FF^;M0]glD8]VjZB>?dig3bKZ6DM4@e:LNp[88_`7?D[o@e
f?m\4^2XCJHB=M?^4Io5;_Lc7CiYN\Njc0kaIMZ0<hV?WlB8TegZ[TaPaPJhcl<Q
ohDKX4jiV[M9S8g\Cgogg8J:oea6l66D^co_hkR?n7]WnYToLn_SY:[JN=\Fci_Q
SX@TRAM_XC_CGjEWCGLlpnRIVIHYj_;9JG2]7@4FllMm?M8H\]JE_3cS\K<:WFd:
^JH>2T<9L:kiMkEnX`949nPDWD0;<hf?Nb;Q9U[KhI5^0iLXEJREok08ajP1MNiQ
Ne]G3IOakRhHQc7gTfB\Q[ZNRY7;Bh;g37nXQZAmAfSR4NkP]JIBepIMf8\_=L0:
MAUTcF:XdJ4<Mk2^b<LjdQ@BIO@G2iD]kK0N3W;[hcV9CMWAF3?`imIYmi]1f_HB
^biGg2^ag>[FS^U6WK<ddE=^KS@IcHSEFPAfobC[PIFc0Hg[PU2bcdW2WFL:h7HE
IbETiNRV9B`3`?FDSE<<Riq]QaBd6I@c>D3i4RaiE\^K@\oYXJ4?0Co6o0ZfegC]
Ujf7gUa`_mUNV`^nK_mmGXP]g13FBfA?iFoO:`8;cf<AJ@=ZIN6=eCeCKfY8lHnQ
ULVGblSgE`>4e^ajfDK82[gSMmd_BEn?YK\0P<nKlWj_3BR0O;:=NVBqjg40FQOK
;=99K3AXG>UipRmL_aTm:Z?SFWEHmE^0o4SE?U\`dKTa=\dV7aLd=O=mf]:289la
fM]SCgG[DVB4hR;@7RlTRkmIdf81E:fI_MC`Q`@;]0KalhTN7c0LaY:KkQ_kL5TV
a8l<?:Z``[mbi75VRlaf@kTE^EOJ65in:0^7RnB:<0ViMplBeg[[<FZkd^lL[<V]
l6b;=YhSJ5PZ0S34hSRB0QIkHOcidkG64dSc9_bLjZ4OHIl=@gnTZ_o00:J`m10S
K7Qj2SUOg3=a0<19LcUS>LN:L;YY>c7E2JNeTd:Z45>QLEg7ASinL3o3D3bZkc<4
0_f1bYAXO?=gVNp?kJe73;]USka8EL9[J^5jV5PIWn@7GIj59<lZ0<M^bRnk9W3I
PeXmFc^EYYF4POe?akFXXHP0cm>FSFZ7CU^<h^D;?TPFJIR=WHe;N75TZ\CZVILi
EDObMdi7I5bGg:VW3NfJdBI0^O2cC^XN08o6ZJIDc66F<YKp?\fL_^\d[m=o7mRh
mLoMH^h8:NQ`eEi_52@5Dm[XiREAa[j3m3``HfNj]>O]G6ib?_@[L4jBY1k@nNOk
98YkKD=[G^]J`Mi_?Qga_e``8I96\5o:@FS>5YMc:O2Mc7SCX0oMQWFEY0\67`JD
A6[AnmENJWmc`fM?pD0TKSdUG0@LCAd]K\ig?hBlKOj^AXlA2S@L2mk>B<6GI7cl
E7MAL95>APf9ROk7PDnnIKO@lL=]d?IS<8YIPhXaFTPKiR7ANS270jLO7jgf7=NP
S\Njjj@UO[2NMD19TO9Q\VbPgLQ1X8o3AA?ogEoTDQoYiRcfapiF;D7VVjZ69?J[
aefFb]T`f?U]a4o8kfJeiJdeSgZaGTGPeCEBXHfl[aegn\oP?gi2aHU3eiC9V\XV
K7X\QYb>oRn`55UhkBeaeB<UUTHk1d9=_EO6cZ4hQE<f_M6FZBkTVIi53hCQ`nP:
^5HeDeMbBoiZB_Ua\mqAMB]^?aNnPDU]iKI0PH4Y57X=e:E5mJYIaQZBDIK@51CD
[;CVdV3iCXG=K7?kjO9AUJ`<6@nRkLV_cDmW`GBlWp6fE]jf[PlE]><>a`hVXSI:
N3dPm^FEJDNb33;ZT3hJmF_Q0E]V6T>eL;bW0CXf@DF3akf3OBV7\cJn@_2R[`UV
17DH]SP510R]35DbDl6@`E2D_lLk8YV>aUf]WK<Lb^6Mi]kknXb]aHJ3VSFgK;Y0
RBRdoClkV=RdHBpnoZ4>a8KgY^hZPgQmF7EY]o0Gi\OKSahNZYERN=L8amLDS;I8
oIai^40ca;hF0VBf[X4kXK_^Jl5Y>eHom\a8i;boiQPN2dIV\ZS_Ch\9:n`XeZH3
lGCJfl;AT;c76[N[90<@JJYk_J=c?2Io`HG`]RO7G[ZK`K3fi=__So0q59od2mNY
SFAeTZgLH^[UN3\2CV`l4Ca7<kGGn5Pe`>bkhDp\m]Wm>5cEFjGS]YRP>4]Lj1T6
ZL;R3FW]Bn[Oh8>C1UF_@09MKn4^kfmKUb4Mm_UP4i6\Hn]1IcBZ1hDlQ@L??;1O
h[GnXjUb^nI71Vkj>9]`iJYgV\NfQI0Ed1n2W7I\IiDG23?N\<4Z:n_L^70W7:II
NmM5l0<bhk0qTHXD2e1PLge\_^\N<LL0I8Mi`E;R^GeRU?gk`EZiWkLj`:BJPHVX
8YQXiT>VlXNY5`ok<j4Dco`CbgQ58`>P:W04gE95@i@5UoOEKh;IZL_QT>>GZ;G`
^;TjNHd^C?2MQOUMCDL<AEA^2f;U8cI4SCJ8CcZ9O<7oD2XWKNdBq@m`0fc5<MF^
Bm@CG1DReTNcD9@gZK0Z]n1mV2W;W_\ZQneSi[O75OlJL^oWP90CR76L^5GDZB17
_0l@o_4gT8YA]OZ`^;3FjF=mP]ViCi]Y7^kclYm2V0Tj<VB=_Dg^g@fIoLN;3[jL
;0cAYG8E?lc<hHO=KJINmF4LLp54gPl>IUIaOlJ4PV=@KjUFo;HLVmQkH`hY95PZ
m`:WDCaT:Zf_jfmXSI>OF0Oh@1SS@OcB^MJC6J0h92gAgB^aR`fLVk[:WWDJo6Gc
391Q=><ifCdA`o8f8F9?JlJRm[<EffJ;@lg77IQJA5gfa:4I_mFaDWo4a;[g9RG4
k=qOK:OFfJPU0NO`JGO]<`FiWK_fFBgDkI29M1`8da`6^ll8U4Of0U3EMIeN5@\2
X@AZoWii4Q`VXmQU9AdJ1;SGk^V^F:oU<G9XNoe=aL>SSTn3NKMdCZgS[E9[b0a[
dP@o1I84[9A3b6h<NVUJA@OJW6DaFeL4Gbnc^l5=[cUp18_5ge969=Ob>@OWWlK]
[?0SW]X5>2QJncPak>^]8RU:eA`k7@SSG__CD6go`02kIMdGD>64NY@SVhD3:dPM
XURI3]Xj3naMRUm]cO>PP;5??5WCckgCkMdJKWKD87B>K?fkVX7]Q5<CK6\V:?20
J?PV1ToK2C0l127fcN[NqC9<5>GGD85=gae=HIcE4D@9^]oKdBJOnNCKA5RI8ABM
lTCDM?3CBRJ=:]UK?Y>]]aBM3H7gf4k13NWlE716^=o@Z:<T[CH=IHHKYl_]MTH?
^O[>NS^@C1e31:H>bQQR?C=PN`NbLh1>DNgLL]5ijnAHK4fkSI]V9Hn\\pJb;HI8
_]ZdQm;f362WOR>Q@DBm9_fc`j2TPa?F]ZFl^:jAe\dnAl75D5_RICSZb^6n57^D
W0NL9b^CbfbDig0P2BeHCS:e9[RaPAPIdO1YJIk21RknCAI30RHjZJi8\_J9^Bom
n@^g_g^=3FAWV[fS0;6PPbZHJgRmbXqkiIWQkYho[?]G[J1Bn:66;8_fWU]GLQe?
44APGZ=DORXc_n7>U>?J?22RWM5X:B44O`RANb_6kaM4Qb883BfHU6Z?iZgN@aXh
U4hfH?3_Z1k@:_]o^JCj;l6HM]ZKfSFk6mTHU]1L9VN4BmVgYYlcfFT[F`gmI^Jh
D2Nqm32k7JRW\;?o\\?Ii>[1hA]5QJj>p^W9_G^H;3ZMb`DG6MKYCb`fj2KiO<f7
>W@RfK1lS6jbYmJ6T3aBP_>Idg\bO8LVj8^LLY5no?J\T3CXN^iR`ALogKKiOFXC
\KhS6H2Jnd8Fo]c:gQZX@H:P^5g5MY\N7g?oPdEYo:ZQLaV3k^41nmhZ\G0;W[O\
<dMPlHoM4q2MmL6SC2YhGCOEh`=V6WX@PKk\XOADXZQd52hU`nGDDdG;j4[S5Bi4
fNk^eK00XOLnjS_40^^nlHXI9EjDCe7J8KVe4i?2:=lm5:D=Ca2DDY]EA?E<bUVC
?]J`dhQMX`2LOHQQN<\<Q\X:=Ce^ek>PAl3^eE:0lYld6Kpb^7`7TV[an29`e1;V
nKke7F@WcPe4UcI;9TbJQbajeT5o2_YA66K1X=alkcBTW1F`>Obd^E^XDO3RDiEY
R3boCWDf3Lfm`?g9^TA862eeBi?9\5BBNCUnENVh:Y3G?J[b7V`\91db:X@RZnA]
]eX>j`mS]5=h0Mi9lPWq5fC;YheBd=736icCjQ9Om\MZVB<i2>im`6hLeYoODmV[
HXHiJf?>gghilk\o1:j^9UH7\7Z9l]@XLho7el<_^PC^BBLZ<E29_Gnl\045f_4h
5>:7;LXBI2DNKOja6SK5KS_6;g:e0ZS;`IXieEWOCW7JY]mCi]Qa^ecl\h@NqONc
]VGVJXmHVBdS:N2WQa]8^>aKHNXFP:NZ6S[OK0=iOVJU9Zj4oJ?oDRmg\RPlDi`O
iMf4?LaW>m4]8kFlcmOVcGaD5][[GH<fbH\Y]5X36:3b@f5610`8m<ZXMZToJ5aA
B]Q_MA57I3Gkkk]]WP]HjJPZjb5][9R73HUF:q4gZCd^JBe;NQamKCGSW3^m:O9^
0J@KVBRk;TL83PCTY6G:PbPkmmX7dOaMKEeI82@JHK;mP`K;E9lX0BOBmVG\0@eY
lh92pmZe2UTBgc\\^JCdE5<EfJPg`d4:AJ\6HRiaEB]f`<aA]cScg05Y<XMHn^Oa
;FO>om^L28S=mg;fX>H0WhOODR>n?kZ<MW]6Ob7bHVbA9NH9KX2PA4>7LgN_fKbV
]]F^F14>>i0G_gRjCdNc2k]FRW=8lkAYBL1m7_2YMbn\<h`:ZCMo\pgBVdCJ2<ZZ
SeTeamfORmKf=Z\UU0qWRO[1ZKHfOlXQk?PW=@^Z6P04eVB1T\AN7R]hegfLT61L
3MMWE;fEWLc0k@k;W9[WBG[>2XoG@][gJcF0@f2IDGdf;]Mh]\k_2U6UYTjQXGUL
?8Hdaj@N=_=R;6^U0;QV9GVmdYlG_kRDkEI]mWE_DD7fDM9DL7;cLXfVbfKbPMRN
>?PqmUX^X=?26I0@9mehKKYL;R3lfh_WccK`W^LG3Qh8PUA_1TXYUDD@3g5[?O3M
Y9YVm?;hII61>jHL:W]VFnbQI8RKFoOCEDKBbAA9j2ZAB[=Ci5Cf_O8oZGCKLKGR
`kg_9>4o3kjT>b8N:_SEIA_LHafPF=CmS\7Z1F:\eoTCk5Kjo?`ipYWi`Li]TD@D
JX^\_<k3<aL20285iOmJ5L6ME20;VX;HaeGMBRHJ9EH7]1CDME?nbYUZM?`:G=GN
oMAeY@[YnKnjcfR<d>FJLL4BG2R>c@iS2Aocla6IIQmFaHS=kc7gg_jK6o>FI=aN
hk:[a_Xa3cjeafohD5lHJQXHS97iK=U9?;bkQq]_ZimECgheiPTU^P`?ULcXm_o3
A5gKT_9]17>[RlE`9HJgJVPXPZ1fRP146gSZMI]:TS5XedNIjD=PGg;JnS83B0_T
UE22TH<b1MoD_6k[AfGB9jGeiL58dY\\^dn;gR<L[`eDh<NCZWTTf[EO>g9Z_R__
c1DE_@6CC?fJ`=BPkA97?GqOiUoUm6^1=0Z:`VbN;;n=:BF0DkYX9RUgW[MIR:e<
NO89ehE1Mj;fcdU=8CV`FcmO>Jmj^3?SUBjJX3QnZJlfdS5el640@RTGWC9LI<<B
\j5_3dmYWJ:S]6G1hK`I<cTZE[HIPZ8S;CF2k?X<ZgCe3j;eJZIR67Ag\jOZKR3M
OT1KjgkqKcX1E<fQCM]Qb4a?kZ6G\Dn:`GA=XiYTMOLlY5`SEM0U>Q`T^X;i6ldC
e?35m378KGj28FfFA?i1K6l8RbBM>cPoToYH2QYT[jHRmX:@g6B?nl_lKIR:N^5^
ZmWiDaIC92KBM\T6AAWR3IX;\1fLf5`GTUZe]PcZL^JZkG5@GY1DdJY\p2W[44JT
XVha]=D4W3Ze=4Y^[PjHb?[JBnkaRJKiYjNTX218b94km_gg9hfSeW3HF2AMF9Zm
o\fAZZ`Ge=:O@DYHN;P4[_2JMUn<h=R3A_Qa0JIHJEOYW:`\^Fdedi5?nZMlB@LD
Z\HKDO8oTVdm_QiUE;DUi7H6SVXdUJkndALA_2O<cp]<iIU<7SkYhUVAKmi[ZNoB
WI0>d\]\2CkR>5Q_f^VDKI7^qn]k1kN@DknWjU[O6U4N2Jl1H;M7_7g8XdZP[PU_
ndHo6S\iQWUQ3C`AT@`eAQP:9nD0?6DLW>[HoGfjDYc4DKfZV[]hWGb8]m>[Mi_o
[IQVa2^XId779c6G]S>9A@fMV<SY]IHk`>JTLjaJMGl49m=KG[M1UTO@8@iH4iG2
ad9jPH4F7pnCHeE97Lm>3fA?bO6BC>9A5:GISD?Fc^=mQ27SIK4k=CkWb6kHaTF6
FifX8<aT_8n]5O]8Yj0MD8@6Ihh]3Ub9c`;bZ5mPc>[PCI9YKB6^_9fmfPL[dPZ3
[mS_2`]P6m>lMB>llI0Re0<AeQG1mlSS9D;L@Xc@VMd43eB]^]Z_a7;d8@pmPBI3
DIN1\od6a^EH;A^iVoZWhOL9kW2i=h7]n5SbA2_KSd^IB@[_T1=IBI;91MOmHGo1
f]eUWLYCi=K8=PKD3C63UlbU_Wkn`l3\fKk]4oIW91U]SVnPCi;?njD4iI^V?ACA
3lPUUIASRUDHAd_bJh03^F@>42UWU84`6L93LSISYCSq=H2f5jDXQbcfdS<8?_g_
D1YDQ:GK[P[R76f9U\XgR79gfN<J@GFo93Z^e2IoG[MV=X^BIkEY3nQTQ^:C8<mE
Ib:WN?7Ylh[YFNVdHf2\[e6@j@LgJmemG<o`R_2MMJoJhgSHV[=o37`\XMhmKo[5
5OgYNFPn^dOi6Di>lQ]D0f:OGKNLqP0BVR;cbaELRYY>;m92aXl0=R?_Aa09ONO<
`hGQGSnkeUFaRMji22d3OiVmcn8ldPD2]f^AeG33^D;GPf`<[\\9@0G=\>S9cPSf
8KW]1YY[[^R_Un\7SGA<YTOZdS@AW7iG40;;iGZd^C7eT9[[6D2LE0j@\:32WiCC
QmifdGX75cKoapVJGWe>8h32E[Ieej?^PF9^gK_[A27m?_URASPFd8cf\i3N>1OK
Z[T75X=`]:j?eYVEakjXi_>c_ZKQi]ObO:4<IOJ`o4D8?:AnK6bQ4BO2bh6^P_Vd
d7Lm6Kkf\aD7D`EnC1B4GV>_^jEUQm;>Qh@a>aJM;L\3gUcmG[WV>Kbg:G]eO2p`
Rlim]S5Sj>2Uj0M3cM`geTAbZ><KT6n3NXAEIf=_Pi7ZLbQNiWF]gB0CJAVde01`
kBjaN9KTd`L1eaVD`F@`9@3Rg3KR=6Oj9ZKkaDfPb26GWnE\iM`Ue<\o`iZ]<KmE
;@hN8@STMU?dHcoVfgH28e5RCU[XI]P\aQBUQOT4haC[1UBpg3gOXYW<]mi:nZ;F
D69gJJ7c_LM5Rk1<3a1ROLbY\m9:8Wi75IXOq?09RmTMHnXb2jRIPXRBfiQ=5j9N
Z3lBF;@RU`j=?RcDUD]H9d5BQAWE4PhV8G``??jK[iI3=:E^:5E7mZng<6hnYXXK
[\VBFBAXHgU:`4h\YXQP^3QRf>WQHXMNJ7K_g6Y<P9_m3:33c6_hkhWTK8\LbX5_
]>Ng8A65f]SRO4i5XSJ\Qp]B7dnY[ATF6a6W]nN89eIZDWkT;i8nbBn5:^WH\Md<
FiQSPMYcT2g`fP0O6g<Hfm]ECnMF]8gjhcPJLE@IghDj1]DHAamdb?j;O_\9cdm9
PQW7ck=>BmN`Kn_6GB7ahUm@RCK7?bgek=Gh57IM;]JH;^DVJE]G:TH6i]:QC9@E
S3^k5Ap=XIGN>5k]B<8Ui2DQOnnnV^If`<2j]iC[B=M@H10b1U5V5NlkWQ;3eibe
:AXYoQK=h>cN7Q;g:049fibME8o^RJn9U4`1`i0=2igI0Ke8\6h:nKng?XZf^2`C
c<C:oFDQP_N7AW:gU2C_b82dZN5d\=<91o8]AH7U1f42Q7hga@>\H[QqPFC=92:T
MQ:aUb[\d3=Bg@@Rgk2eehROoIQdK:aoJ_]NI0Xjj3O><KY_T2gdn65@P>FCA0>9
TYIhOV@MGAc^Fjh:Jo^T[hRTXL43^A]d@PI9aAdDY7VKbJC3Jd`MXdM8JBl@b24j
Td14LHJN8Sl@LXE^J>Ig\m\EB2Po?<3IJhZR4bChqf?P9h?a67D8cOae5F;YHdBf
ClK@Fe2o9hMdHn9jZUZnLX0QSBH09W7WKLei63Z5^fC4nODR2l>fQ_lKGO9iFb:3
48oG?hGoA@VE?_;Thh]G10<9[;j;k8MZ1iT]PFlEiXAjNb@6UlMjLPCoQIgS_PhT
d807?QN:NOa8kUH3kf8`@8A@SpL2a@KAWNDLNgH]L^J2I1SMVQXP11=[V?JeFYfh
WPROKYKbU3fD04E>WfPHBljeSIL^P9N]\]8VhBUI1RmDRB9AdXbLlf80VNSnn_<E
QoN?j_l8:2aBCSGfJBmUh@KZSaLaP6hNYK89jUmRU^6h`J0e]^bDVTL[WnRE<VED
C4;;X;:GNjqEYIfTMHU6RKYBXpgT159K=_22bD9jGm[?W6[g0_O4l=C\CghdPb;`
>jMT[aDo8:ObZBW>IIZ59NM54`glK[\gOOkB]R>\[QJJif^V2R\;9hXoC[0AGZd<
jhgP23JeA<jc>QgTQ^>ML=jRmJ5eeOWNo<k0Ji^[9;[VV4l=WM\N1C6bVf\nW4mE
Ge`K43o<=EqU7^TYDZhBEMI;TdL93RhnCNPmO:\UJYC78;=gMODX^ZBPU=j[emS5
3NEhB5iCTjmU_\dcoUaeEUV[mTR154iF?KHYLNjoFYoJm2SNme_o=aBhn2Acgho4
kd52l:^2FYm5U8P;?HdeOIAEl<>SgK7GV]YYef^LFlT=QNh<I1IMPM2JkSRqYa[H
>8:WhCXS[cbH2fb4?b6iU8dZ@Z[]Mm2GkGJkQ>NS\_WDl6\YPB`iK`O;Z5N]YclH
@5DQPBGiJRYbCljbU6[3;h;bY:[SIkm1h@P>K43_28cN5k4^5Go>6XI6a]5XiZlI
gZ>WP[KaEZL`BB7lH@]=;1NO4gb8bKHdEY@eEe@P4QBOqeej\U9?_g:383C2g]HX
f\B^L336NlMMRY76]`2O8I_0XB7=H`W_PXiDIi=W6WUU[eid\MH=YUIc352WFa1I
XKADA9<lZ5;M^1e9C3FXf44\NkIYb=`m6X[=?Ynf_0ZM@[Q@?JV5GUZg0MMC5VVk
_S>>K9X[lJF^1@`\<iRnd9YS`UI2BqI8`30]2a><@;_Hc;cH4G:fiKN1CcmO:JnV
inYZ8F111f]De5K<CU7l\V9dF4EPUlIN=\oP=oL<]L>LQA\GRdZFZ=CC]cS::F9k
\Wi1ZWCjFKQOLkgf=O8YmHfT4F]M?\6KXjQ17PLhaL:gDHS1A5c=h[C4DehN8g2g
;0mda^_25_`=1Xq=<Q9OnfL6V0QUaVm2j]J0g8SKYlm=9Z@L_8]T0@2PSiAS[@3I
LZW3AL9<4][f:l==4=>oFRXPGBDmc@g40Z<4?;jBBKmh\ZV]lbP=@^hZV[DmXDgm
C@P_eDnK`[6LXCUbHcClaKjPDVYN0\N0_nL]]]fBKEE<F3Z4C_GOf;ggAA`nGk\p
QGOo8IeY]j\JJ7fL=CO=ikF7fZ9SkZE<>YLX=KX:ml?TcYkB?:@h0k0[cmcBe7Ng
Q7a04;bbY[1[m;PLh7kMJmMRdHYkZKE\G5:RPDJhWmNZeGH1OIJ@LNWOIP[Tf`?D
Z\:Z]RHSYRl3>35jLbcLfl?fdF88URLa_\=:_^^GA7T8;aRFqLQ2R?NEQ?EKiS>6
1?e98U\H\Vc`bW;fS70@l`86BRS@lB63f=WK>P3RMWi6\jna8L_h7>[XO6CdGiYX
a3o\_VmEI@;1C0RfHQgc[Dd?_Cb^7FEfl=[=fk_4i@LOXNYmkWeL::cjW6clmDSG
l7K=D2PDn@=IaJe<cLN=eNWJgoF8VQLZ\pK:oWGEQOSUNCB6Eo?_D=k:U8lRkB@4
M?<TN3P;1E1oE;7[leVL=WC_`XN<XXdZUZp4?YLaDdneDk[2XeO\g5TS5l[XI`RW
eZZ2KecZa2Z>@bC`I7jeZ:jM^>aA\B7JG;o4BXQ]N=I;OEL]4YjPhQ2@CKZTcBf_
@Z`h`AQKmWZGbOUgO<K75DoB<K0d3]@92=e^^>34N`a;]U;jiO:4lgC3VZDTkHFT
O81T7Yc_Jo0jmL8MakBq9j@7DbdBFcMoLbVc2k4=;NN03aBAIZ8I]QY6>H0`<=^2
:lVL:D@=TRgd>iDYc6Q`9TY7[1TiN\8X\bAJWKK`lI>8?3[<f>8O3MFG@8ij62mX
RR`Lih6g0b6@S2mO^eNSWbLdfb>LNW=Ymnn8DHQam5CD?[6S:`YgImF47d]j2cA5
bl\epDdBP?HI?jmkm_i;6U@TJTgE0g8V@nOP3GQ9h4NWe[HiA;IBlE_S<WV5cB@B
X98c0D<hMJ7:4CDeg<jTm<NE2Cdi[fkj@1aPZ8aAef^PYgVK[fA;9j\>6QofCNiJ
OEQ`kJW>@IAP_Ch3:d5BmJVDV;V[mfA5:3MSkJhkBORP]S0_e@MWapE;;94jS005
SD\b<@T>CjajFlk2?NGm8HkWEPB1V:5dEbl:3?GG4SG<KaCoE?77qN2<9I1hf>5W
C:io>PV<i5_ToaQ?;kVkh<[SoD04_^F6>@L8Hd5dVZ3@3Aj08;6b[N43Sk`5k::S
7IagSMA@:19ql\\fGVaC:H8UZUa?BmCXN7OPPBT;@n`d1ecReU8fG25:dbQR<ZH4
QG<@iUaI]ZdS5M1_VEeTjMCM]U[oEgM;9L<W]J58A10_8fcD1QGMD;ZFY;BBOVBP
H^<<mPE3ShU:X[oJ?2`[q^DAHm@NamcT]iIH]1J[8GGXD<1[Tn1QG@XZGP[F:eYB
EZLL2[nJ6b6R3lZ64]7M1AJKAU6AcQ1[X>m[B;G`n^beJ1g4i4=\cG?Z_^]6P?SX
[4NIN7i5:\jR?=kDJNR7[N2gZi2J`pKUYOSd`>fd1Z>0l;CM`ZZl79?]Plj;63SL
Q:WU7VVbniK=T?ko=l`dFTKK7FoNCkYlo51P<9O?HZ8>]d0J^hlKEI9n>Voe?4N\
QkAOFL=mUCLX\f=3`Gf>fT\aJldoY`fcN@]QDVq>ZkCRY<k?G8>m0jMK?;3I@;?a
O:\@QJAg^0<o5Qh8GO0cC^:b=9CaGEZjWM@2?Ufd=UK8hgED86@MnZNY^F47`d1c
j:_0S35C[0`9j1^:5S7a5WZ>o=Qj=ER[Eai??2XijC_9X[7qH8E7bY?\3=X2n6gJ
c7FKQ6P>@b3J:Qcom4Hh=d^lf\QCXe2<ha=LkMXNH0=YVbJKicgWV@bJPK_V00RV
S;HN1RmJIaVLZWEebLHA`@CC_4MM=IFA<CFK6IU^`^[;0ieR31l214@EqWjDmaUD
`]\^BCj:p2J7edKT8F2<]oVLMRQ0R8I>o0;2ndNkaYNORPBTPgMlCk]iZX>7\oh^
1QVCP;R_80[\1e9[0\o_[jZS^0dW7XoJBl`SY]kM:T;OiDLgh1o]NfNH9Le5UTm^
g@529<=P;>ONQo5?Nq0D:E_j^^I1g;[WGNdA<[?_Yld:Ulc=^hkRdO6o=Q8OGhok
0jn@h?S_O\bA2_KGd`]1djgC>F4leg21lMmQE>Ff478]WYj:=L00dNZ3o_79FlI@
8CB5R0\Gmj3LQOSCDQVL6a;kRWp1F4`8@Z`1;OAd15\34`fjIgVODjk2HE`AnlIY
6\@_\HF6B_^g3<DP24[4PI\dgT`;7G_o6Q60Fa^e<fa]0lEg;5\?b^AT<cXHAloM
8\HR<jUR;L]j]ghG8m]Fd:PgCD9@6VWn?[1pOQGB]oWLHe<19aY3JlV<Ol_]W4B2
7l0WgAPo:?I;[AT`lj=nQ?YEf2;O9_RE=R]jNnRjG=6nY6<:IP<dP^O:7RYLP;B9
qjGoj@VYoImbUfjfA>^kC]SQ2lU8:mHm<:fO^1VnkEIe@6N9Lcb4EQ>ZD:Uk9U_c
;2;D6n[amRe6\YOS^T]8@[FHMnjfWAVDSM_O3>;Wad=_S^\I84PP^k5ZE>?T6W;Q
P>[KW<kElpoM8b14g^OGR]g^mB^_<AM^b?eEkM@C94\8JOiVcVR:\YcgEUhBPgd0
mf7\aP5YfLJ;GbIa8QjC`UVf[cUAaB<2h<]20e@fcB^KJQfWlP3gWa?iE=hEMIX7
VGd<Cg_ZadD7bnFTfQqWQb>aRCf>mc[ODOa@Q6T[4Tl=SkoRQGjnFQX^4H6icB`<
GZ]7Lf1R2a0ed42CYk^AWKW3iUg:?heUT<]0a_Uh<oODZ7JFjNgRcQ_QPc8laQlj
PLml>5eodaeHMHN8@38e2lY72dOp4k>6n=S8RUe6_gPQR=hP2F68[?G[@N]9hjCM
2?B6iReJ\?:[kHdD3_\=1bj\l=S@gX38TlpX@B=9Y;Ni3AVWi8aTMYJEVk@MZ:eW
dZN@DV;SL9REooP>`QJ14a683HCNmWFKah^OWkCcgiR9gGE9jZOc_g7G1nOV?4Co
=d5]RV_5OF2doek]8F4L>JSnGKaf^8=OBYha5gJ>^gcqBTbd]\oTGA_GaUN3Y6gP
C0BK[5blg447M6aMhhWZKnAhhljB:7<Yf_1eDCiWo222=<Ddi`5lK2JE<bkKA5Y9
8[Q0A15dgHP<@3aGm4dkh1^MeAjo:\:7GNCbU3:8T?kHdDcZ[U08pjA^Uo:TkFK0
\F@WBZ:CQnWOUknBCUSc[4HJ2l\5Ad]F<3QmlEB>JfBTNAIn6UPQYP_Ta>e8F9jI
jVGD@mHO@KGk\fifBDMX59bJ;Y=V^CVWd59RTG:e1eUTRUgAEVGZgDM4@e2fNpUS
739YHaO^a=0:i2fH8V0VVj=PPgZ^`akZIKS_JEJIfIPUc_N\\?<bhkMJbS7hlkik
<2C<<04UdB297C5C4Z3;INckbY2aS:VVILMke;C7eLSJnVn?k959hk?W9@F44KNn
6_GZ4PqAcP]_5d6>b0QU@[N5N1JEP:O=Y\6;Q;Z3Zdj0\9k93jJSnFiWlkkmRYNa
b6De_V@^b=k:::D81I_JfJW^Z``6dGJY?[0hRo<ZLdoj@R;V2ibCCamD]hiXk^IB
XH:WNEXQml]O7>?p;MbE77fOfE9M_=JJTE9o6fTMK_d;Z]Xf72U7nl\O_P>kBhQl
l3lR9AU`1_BV><]MhC:5SFA56KgOK^gN?e^HSMQ8\?hJq:EX2E<C<cC6CcAN44_Y
5<LRAoX?WCLZ>9KoJdj20i\H>d8:E_KS8coQ:RBBfCK^UZbAo1VZqNTEl^KiEBh7
RF1aNkh7jn\90eddOfel>8>U1^7mci:Lh0XXE<mJb4baTCh4E[gd]Xj;0Ae>O]Gd
KAa2a?^mQZ^@_o;A09AWmXGUYB:XLiRU4N4oj`Nh7f2aam4E:S<BX`]nRkd@5plm
4`m6oM8ZZ0S^XPJXon02kkmoD5LLPA0E8k7cfWlj82f0F:a7@^Gc>FaS6@OdT`kd
ija?LmcE>fj]DddNfPOHP;o2G4M6a5]380N>@5eD^bfEUXn?VinP25WNRHneKL@l
Gmcb=jqJX4lJSDHWBB[Ol;6b4ClNgDR5fWWV^RQ_RZai4\78ggD_76XL90V`f9AF
mEUM=P6]:PaMZh=a@Feb<=ZXNoegeogSSTn3NKMdCZgS[E98b0D[dP@o1I84[9A3
b6h<NVUES0]Q2^^qa[V8EJTL3V\9ZEd0KL^^d5fN7;=[LkCkb\=@X;dcNc8eW6D^
LYBTQ[8[X3IUAFAU3K7EMN6XSi5BnO>DjTGf;e^1XcUgP`XFYK=DYPS\N:3;m42=
2?S>gY[56Z[@`Wom_5HRObT5pV^NhZTb;S]3:58m43]^R\69VNPRQ@^WQeD\fak]
2:m\R??;n<bVCP?`S0;BA[;9FfCeU0e>@A;WPo;EXZ7_jCdYTCQ1\\SJSOd\J0?O
Z:^;IggEm2YJYE3m@YN;03]5PWaB6HL6\qJ2baIi4i[6ljUCT5`Y>LPN=k><ElJE
3]0ji;EGO>:`TFWK2?FDn:kIndMcZ=^[flSJ3PdKCX9>6oclnW;=OO`WHL\DoO44
U?`6iJ0OT81fU_G^oRTeih<;nXE1DKe42W_dQQBBBMq?X;cAl?4bASdADP3TI]Sl
fgagFTm_XM0JSEX;hRgWF=VC5G\j7[G6h<n_eXGGnE?Mf=j;`ClN`05<9ceCXSH_
76UURa:j?CTeGEOQ;Lfl^dGLdFCFcgl58<n64]ad4I=>KlXj799qjZjZik_P9Hai
?ZoM]:_CVC9GSTN_3_AgLIZ;KHKEa<4AT@j:a2_@YZCJ@`mYQS`gaRRjXnn=f]1d
Xm2o_f?9?2[1M22VTWVln;Z3kMC>1P`=E7G[nQEkB:emiSCoDc:<7\[`5PFIq`PZ
JH[n_26\5`U_:OcLO:`<dh:CCQV\hb]27o?VX^gk2PcPkXN14E[W7n47]b<gBPf[
K3olM5^kBKj6YL]Q6SUT?RPnZq?T>45TNl9cFM@KHZ>L<h9hbmgDU38<JApW=7CC
Cp]PSI4mN$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUXB4P(O, S0, S1, A, B, C, D, EB);
   reg flag; // Notifier flag
   output O;
   input S0, S1, A, B, C, D, EB;

//Function Block
`protected
j[;5GSQV5DT^<HTh68Ydi:FK?iE6^k]3nQJDIdP5;NJpj:;mH`YWofMlkLIn=@AB
ibRkl7UR4RB^9iS2H5DRl0IhdNH4^HabXBEcPVV3?]9ClTgOX9GqFBa2dQEMf7`;
\?8HWH>hBLigK]@9Co1XXJQeEQl;Z548:m;ZdB`g;:Q;=\CB7GXTkh2941p?l<gD
HqcR0`FeD9l:=7G>3D5Ua?>NNIV=iGTH2@h[gH1NL@dm]F3S8hPg]mZW[4]fK<c8
Vkl>q\dS2RQ5ULjUW]``22M>6`nd=D3pf9W`iPZYH2oLjh@RGJ8lgm_n[fXD`[SY
R2COc3@V@9ZFgMDo3@dDY_Nn9Bp6^J]]XHJLcDGU3VN>55[DY1=`>^VU5fqoWUML
Jiq1bSKgdpfY963_HM^7bU6^UBBV7AFhRbZV?GG@LMO6;\mhl1X7SoIm98b7[8c0
1jQN\6DPqEl4gg2XcZIFN1=44\H69IZ\0deee^QaG]IV>05DOn8Ph=2[2BCLf>5_
2NjOT6EZRX;2APSjjm<mQ8^YDjfN5Z6dRnQGTccUYh[VISN4\NgWjVN=]Hi=oC@D
:gV^HA5lo5dN^91=fq:f7[;<iE1mLb:=U@ASN<_0QgF]>ONBeFao25P\4J8LZF4<
EVn7B^eIV=@JRnI7h`3Tm:dViV3TRSV8QdLlRFh=6U^Xo6;J7T\n2\8CR_97k4T`
Y=J]\?IoV7c50I\TNOL1Ri4@@Vqoa\^n[fgMV=FhLn_8A]]8E_2^6KjiMdUlLB\W
?iAo]A08;eUa\_<_\hYifY\IXn=W18`8Q?8JW2:m:=6Te0REOI;YCBa6dfPEoBnZ
c>G?GkC3N=^@6FVP4h5m7_k35U9i8><dGTNp?eX3iehO8f\E\ZEVkagkG8mMb>Z<
<[j1TY=2fi3;fFM00N9K46QN6j=X1ZSX10SEX=l4Y9LJY1n:amOk:_bE4D<\;?GV
RX^S^[=C:Zb`gZ?N8:JbPDf;Wb_X^`Q5f:<Tm>7KZQ\`qK`FUWdCTU_bF14d2]32
o:d6k9[Y`F<ZY1ocFnKSDInb?B^AI_haEVUlTBeQTK==;QHTj5kR\I^YO7^J6eL8
o[J1GeChGbFgc7bcL@]TcE<aKXJ;<jEaO@;l_`D9oMSLQ5?ZbS^=@p\UNUCK;j6b
coaIZ]E7OWgReCD1ZG]@@df9?liYadRL:Ad0kK1ZAa`6:V2@:aI?DZ9gb7SYeML;
^aWgU773BTnEhhS3:S0=j8Li??oQ`KF3>c[iClXL4[G5:g6C@7>APTgQZX]PXlp9
Fch9:O3VZBc^ImENLRbhd[b7b[loDdI?FA]9nEG;Zg21cNj\CUmFRPdWhH9MK2A@
0`^U0W1B0:iGIZ6deEj]@B@9Z85]`SVI8AYLcX::M?4ZS<=0JXWS]^o@`IWmZmh;
cZ`mo:4pjl:5h=jIOf0T0Md7m=JcN8e]MC[=D7Uo4E<PkN;f610VbLJSAUfjWch[
G2HkAM^N7l6qnVIX<ElY^Y98EMacFgRMf26@?EUF[ih3eJn:@e;dnU^Akd@nLT6\
4EENWmUhXmPdT9P3bj;SLOdKo9lJ>B7=nmS0L0iWFn7N?6nN>?i@Ue=a\2>LT]JU
1EE5TekUh\1<DVATOCBdq5h5]YJFDNNXD6SYjV\;Un>d38QV^ZN5\BQ1YFc];[2?
7PI1?cTjRgB_>J^B9f9`_B0^9lIPAMZNOjWAeL7chZ6G_@9IKp@8:W:FJ2:`68b_
;On1X8H_VD5fNb\Peka=@:j;2=_fff<h8WVD_0Y[^E4T3VmQA5HWln;n\Lh4ngjh
H561^>dXkejf?KlX:EcL]lX@:Kf]4<;@Ukl35iYl>3@Dn`N`UZ`ePICCJbUE=kiF
GV6Z<C:^Q=b:M?Ol6@e`4QXaH@pTil`hG@_OFo[5]L4J6l?c\g?Fh9MD;E108VL:
kllTLGEa0hDJLDRO7c\9C49=KZ1b0IHGS9CMRD3n0;^XTi7@Zm4EWDc9[Q[:\VCG
`3IgYEN]41VH[J=C;aAe``<?SUUT<>m=K\N7;g^n:@ZH]3@=7ZV;f>X4LBj:9X=p
BEGDM7XQT\1j[O^_>:lP=OPifQ@f^^<?gl][oIiXJSgE_WWIm@^1pFQk@k\]Nn^8
Q24b_\Y4^3GI582W@X9kG4AiGO4bf]lB?3oQ9>g9YkG?Bk_ElWAknORLUAOi4L=4
@nS0SoY33nY6CS20_1CP;?dRDS`aHVWb@X]g1fgR0OR3_A;ZPCHK0I6=cJQ]`I1e
Bini5o_@<[1kSbUK@82^j]MGfSPSRpG]A2Z?:DFHJ=kDA5[:>AAT4\90cn8FA1MB
oFcUH46SDnJK5URIdN;UnSaHPF2db>0L4G9EL@<DfQ3BF;Q:V>aW@V^0YkCRE0RT
><7bgAgl;YF5568R_[^Jg<SM:::YKfeU@?]T:R?dUTn8_UQ@;OCTX:R1ekBWUIhA
cl7Z\Rqfo?\XXE9b^C6[2T2A`cgmaMWINHHY:legSeWhd`gQe\7Qg_GG\UQ\n8o_
8Y[J6U3d59o35BeZJiWNjjodb?mKb7??ajU?^mQ4>e6o]A09AWmXGUYB:XLiRU4N
4oj`Nh7f2<]m4E:S<BXN5ZV^2]e]>ZO54HOfOLk4nGeqc8M:3\Wgn1]CBN][j<W]
DV^jGC6YEio[ho4`2Y5574hiT0ZmUXBJKkbfk8baDlYe=RSSEkkQkd>;PaBLF<EV
@;8nFC48\d3FGiXALcbAOo@n9H^Fk]6?7gT?DE6GMT1lEaNLQa2AZO56kJ7FF4SD
LVM[`MNPK^9]8BG^LR0SpaMGQbg_D1O;fW3L9O[mdi<7`2Kagm<0XoOKofoC;11>
XQFToa>GX0I[CIa`2nbT873[KoBKN]A9?Mgl?SM`dg8[4V3EMGM>OEdKRNMkA3D?
N`]N4aNN?V\;ASKl3fZ@ma:HJh\Jg`k:dMeOUB2HXTZmnlYnie=L8E01kpAjVG:e
mYg5OCoOLhIOb6V3fhI[1R10:]>D?2Bil8`h;gS1IRWbP;4kY<8eORb9`GKA[V\M
VRKa;c6`9CccQZ1\M:SXVJDGJ?MD?BH4dFlP0o4HSP:JU4j[e2O9;l:5S>AKSgm<
0iZa3L6inOa>NU@:nG16dMUdTHM7N5pRdC;Wg@;1;NWa5FC0nQL?NMPCE64l7[[_
0XDFL2OB?4hd@@1G5l\G?\hYBCAeG[f_fY4URPQI1HRBALc4PWNn`HLG[heaUGZh
nX9gFjEi8>9loR^K`fALhcQ9b=<2OTBRSF3TA8?;2f@BD@D[G;[><Qcd9_]XLkNh
nFTp[d]]i\\bK>cNgZ`>>8@WnU]kliNOLd`hnB^ol^^:a]h8^=i@CNFB0OZ`U@T3
cQf2KJK1WV5:ki:j738Im:n\6Md60FfT[]bB;1^GeeYji?=Mak6iP3I8To_^eZ^V
ABW0[hCNTb5L;l4N7a1AA;_VjQS7]F8n?I4U;;oNq1MPF9F@4knCm2;afZAVfl4U
<Z:_=3<2P6cO546O02><Z7B_F@9MeF67UE;M0h\iJR_]HjD@M4mjIC=WmCA3fNKc
QR:bTgXh3NGQhFSXbCn[jLV9a11<>^^:Odn1_;`RNOT1;?V@dAgmghC[MC0]f9AG
Y::nJP?3Yk^n>FVPUqc^mXDjUY\OQeC>:VMf5PgBIVJV:n<YK1RNg:bfB8j@U4lU
JpnhYEUChWYEFERO=;VW<AgG9`M6OH=9M1ef@:8Mj?2^Aj>DmBG;7j0bmOe8NeP2
f0WC4_VdDFbX9ehIKD5nEDad6S9@IVFd6`Cd@3Z\aP]P_faVWaeZQL1g<afR`AF;
S`nnmU2Y@OK9ZBh?AZ7g6:Oo??Ob1h]4NXC>MKpT?0aQC9A1P_^HoSHD>@M`\o3R
CCc7IH`fSEOaCQN`0Y7I@DRT33BO9:YCbThAkln3JQ^nK2o<g?c1RhNU>c9kAn6h
CFE3EYMaEmKJ5_[1V4bKhkk3CRTMC_Om^HO1?1Q[13cBB93NJSN7j_0U?]GADgkJ
15e;aRL@nJAJ8h[qgg<<3CBRG\7LDLPFMm:LQR4RLfU_b4>NXMVoH]MSoXW@o^@2
IK49j[j<gRW[4I]fnWG@TKLU:m@QYRMbP\Y6_B<[aH<V;64>hZVQOM4dK9eeV;1V
nlQKO3`?O_gOc2_dg6Z46BENOUQnYTf[><B>>n8R71N`5KT<h]RLqPNhRH`Whl8c
YcYLMI2b=hT_BEg<LkNjFB9A]7@253iTEc@D7>Y<WJmFF<PBA1LMla47hIMcKWBe
B3c7fh2BRR\Vo=g@kKT7;:4BMAk^>A5[=JZ]1P1mb@^U^XOgo?7Fae]E2X]WX2ao
2IBYhhE_TiTBjJ:SACNf:8c46AgIJqj]Te\4Y[F]PYWhH9b32a;0`;[^H`=JB;Dn
Rclg^?P1bWj`m3GInQaWPNZQX@3mEi1=nUJJiSSRI8[`_=m36KKhRoc^dD557V@L
h`dHnkb<EK[ijH25SCT[C>JnoQalUOBS^jG63f<9GS0YMfmi5oQ0XlmlLnaQUGDI
SZd9Fep^A@=;2F1>3f<GNl@?LWY9F4SQmWL7f7fjDa`bRZOUcJEbeh5kX?nH=:_g
Uj>E4=kZ7VS>TP]CU4`P>GcHLbS543N5RnMncpfjjReUHnklR9i7p8<K2?1HZ@@M
]Cm:d<0hW4P=NIkPLj[Y1mPWPVe?6K]>MoENG4glHEP;kK<P>a5lDcKV;BJkK>Le
aYH0[FPBTMLLCnkPn1QnK047S``I;BNQ6DT\STO6L[@9N1]kQP?F:Uh1WKDcjGkU
;[DEfF?>Y;W>SE2J0bbHi9]Tl`[0dqEGi0;l[Ac]<Jh8NLHDZi\BDedQN@=:dYY:
]b5SKdXQYQHa<SCY6H9AF<o=1^E6<XWA`X2iggD\k\4\4d?DN?o[WB^Q;=>n]h__
ZUJP4@[?R8YEOKR;Zk[`Qg6Q56UO5=7S9`19[e[j\7@YkV?M^gWB5jc[S2Y3AQ<Y
ahJAaQqd_j@I5jG_hT_F>ToVE2XU^`]FHnWJNS@TV[>3=9XSJ=cjg4c4h1]BQd:b
MJgki<m5F\D:CG;Ze]H9?iR7?e[HZo4<H[mUm7_QE0;jT6PFSV44LRHVb5FK>WN@
]ilfPKG[2@oeYhF?1afO6]477PaC^@RODE8ZRg=Y0doj7FKqHK?]J1EjM\HFjLlW
_PLdP7G<Kc\jW:YJ\>jjLc4Z2O;Ia[cXTO<8gJ4U`oBYGF2241gVdSH_4kDKS>b4
@bRH?dl3Ac@NfGKO^LE;Gk4mS6QI[N1UZT88SHK<iZo1O9XJ?^BWlQENX6WK=Udl
@ZNHHc:YI\5jW94R\FKKGSD`qc8IRO65LW?nFeX__Y?1^IfH47fZHGW:Fc78e\_E
icEfJGhO72@=CAjTGncN2TAe?DV9h>a3J`f<GRCOCDZkSB\QS1fkPb0B6G3ZDUGK
9G<WB;1F5BS7MWNHNBEfci<1N49@AI7ShP7odK03eD6G7ff\\Lf9gh:iBdoETU>S
Eq`eWT25_Q5YdLARDEATd3G<MNb\VoNN\[]<ZfbPWA4BIYMSnEF]88O;FR<njA^V
nbi@m`QPoa\I8h>GHS_QVf?nhel\3mB03G[jVV6f69Z8UDgKX`fVR_cLL[3[A[BW
b`JS`;XZ_L>0U<fK?e_K[f8mT14T\5NUiTF>9Q6YhDpoZ38i<SN9SLUI_;98cca9
CSF`Z6=n:e1PH;5SnX2kaFM0_ZBEl3Y9PUFX@SknN59H@ggQUYH3aTOodk]3l2WX
`\5;ZeM_;l2[\dLSjiN4F^j7k[h>U4>n6S29HKR@>D7DFm:^6Sn]`laQQ\X3FoX3
C;>UgXYnCe5`WZ6Sa7mqjc1<MH5K<lQ`;6<LjJWY<gV?_T[2EDcKiEE_O>1JJ?lE
@XINn4WddhYXBbObG37@:e[f0O8N;XkVJAhO:JeF6Wj=ETCRFWc_9LW4[=fIlV]c
3C<0gAAciZF7A^Q?`kUl`A3lBK5c]iJ_0R;2:IS:WgQT>S^iLUIFPGgd[]_CqiSM
>AY;<Yb2Rh7GRmH9cb7Lh6Obh0X;RI>U3k7eEUUgF2PRV4mSeCORFOi2Z5>7\67M
JL2T_=_I2VNmG^86c1JiOEOgLggFNioo60aMc?9c]m6O\3o:U?\_4iZ[0`^]jHSZ
c7j=HGEAjIT\]^BkZ8eR>b6SG_Ma;3o7E06\Gq_`jM_030=3bWVQV]RVIoJ8CSno
O^cNanSLb_YO<6Dd40QG6Re@ff>6qYF=GgVV^Am@]Ll^56a]QS>dPR2OoBEj?i9Z
;nQKdni91Q]ifaoUcQb3nBe;?_M_=m]ePP[^Kf^5@Ac<;@Ccg1\28D2OGmf@lUNL
T9LBR4V^o5NbJmkikT7;B;AGd:j4\b5P]Fh7G:;R;Y;QI@2J\;Al@PO3]=UD^VC9
?9Mmgp:a49e60PMSmO3^XX3ke6c\PgcoI0B6LD5H3]a=_KG<jK@_9d[EgEIV^8o^
Ro0ZKL]W_4NHg5`\>[jmLQTaJ?Vj7J?oc:NhH@mF`=23[H>>^6[9[f_[ilY^OD8>
9PTP_QI2f<]?09J@MmEleVT5h0H\k3Ce_XBYAUD5Cc27Y9p8l;`\MfmMfFlnJZ0k
[<g03JbkV?OoU[73m0C>E\=ZYaj=A>^<Y7c7l1?D?RUdlnc5WbbJU2jComFZBLR=
60`WY_M5VQQ_bj?T3W9g_3MMl8I^o[\NK^G3Da:hQ:YBkW>ki4fORf[R`[3ODjf=
;PIm?J1QgHHo6A4\GM\g=SNq]OMjgbX@?`Q^RmI8_AQ[TiGjNec^939=:JSeF:`<
nfLUNMW8X7?=jc^6El88Sm57E?MFLdC?^M4[ik5hm\Ff_h5D2e[VGZR<2O[5JDDJ
70]JEgkQibb@LdC;PkXLaEe7U5bbdV1a^Rk77fORmM`a9i4LJ81fFBO>1589Jn>K
pcfV?11c6gH?Jnd6EH]5MLOW?io]LLd`;?Me4]Be>RC;QSCMFGT4UM:T_^DYoTEI
6T5VRXKo::\iSSJ;A15mWI:h3eo]5IS?IMVf0EN3;Feg6eYTI8mog1MKm1`ZF=cc
mX`dC4G`?:`R;`hi51D:=cfABHdcWNL5_9e1cEmd_p\fnLDI\T3]7L>^5WERWSKN
ZhHoJf4Hq2d:jP4T7DcLB9N9YkB3R;oANBbB67daXKm8?4<DKH3OZ>[P=h:ORhWa
8E4EA0;42h1<PEoBL5F]J1G>\MBmlXEo?Gbode75:JcRZ52RUS9_L_dGD4I5Pj]f
T8od^<H]WC:MOQ\ha=aIah[JBMn1]PRjo9R6n`E<<l`Tk5G0]p@0P9B2g>8Se\6V
U[4[;50;nhgmG6<05R[^=T5c_kF?icoUYSMXgK3?1jMji8dfVo`l]o8dUB\59k98
YE5@49f4BHhmG6E99nF^6GoU9iJDIGnO@YNK;iJJARYaSY1]a4<K[V@DgH]^eU]j
9H5oD:];8E@Q?d<5Hj\Nc<o<LfqT67dO^M35\LG61e643CNkY;EGR=m@X6FD6m;;
Z7SNVcBDj=NQok_4b5`JnSmN;YoU?7m[_8cFFcM[cReK1?\YKgZVMUH;4pa@N=^>
N2E>6?B3_OQ9=eIefAXhh@H7QCbk_hR@q^4Y3\Th\[PXkh1o=l\C]6UDRe`D<YKM
7`7_eTml6[7hHgFHJ:nnh<@k;WOm2cake^PSPIgDZEeGYhHYjA7EXE>F_A@>H4RM
oOfb?djC2NQ]EMMS_?BKWB^bfi7M@jA56g0bN7AHTEZf5b:Po:IakC?bGAVgLFm<
@Q[D^g?\<OO4_F]DZql_^6L12gAc79bQ\F[:eLZhoGH<HM@S44Y0MnWfo@^HFYR5
Ch;1?QkRCgdW8;=o;XlfN6oB;VYZkbkRUjV_eo2kHAio=F694MjUC_`dUiIPWIDQ
1c1WGoiSnNAC>IC]_ATUNn2=nfYhcE:Q<9YCiXNk@0i_M`kTgoI?DiTeZOOIQ<@4
;Mq2^L:E5S5C^Q2VT@TlPJC3Of[NQ[OB>l4V:7]LFogiG8J;[n\j\]k_RdL6kG?3
lBm2h4U`TbI7Z7kKUW0WlJ5gW9hid`BEMlW7Vdi<Cc8SabT81oN<oJFH[O@NjCfK
ICh6_<eLh=C7=^H_M\DW=n\MHRUiFn@g1MbBAcfIGXPJiU07c5Oqm`IDBJnD2c@d
@;^><2@GBFdd;2@;i\7bFn>5\OFngB[OYjG_K\0QB7fm89\aYl<8mMhYABBnZ;fc
^`31E@D4KiB_XT?GDi7OWdK<\C;ZV>bZX;o5GkIeT]XoI:8T5DN?3H;OVN]OZN_<
Y`O\9W<_]4M7X4FoGbTB`e0P=nLNaU3d1>RDqD>Ng[jl4Rl=0cKiTA>Rk8OKVeRN
A?4o]GE90LoS>h_ATe3TMcILWTOn4o\W0C<BWD0]hMRPgB;0lkOX?KUF8Q1HbWUB
C];o;bg?EFAGfJfM2lO2M_Aoim374FgEldbRd3ZRV1>7OBmk[k[PNONT<Y7i[WN4
ccg<Vha^f^lRMMC_n^JjkqCPmRC<M`B]eMPaJ9Se:YA1OR9lCQ?KK6ieRYbc4876
cgndY?bM`a1kLnjL[MX7oqDZ=Yg=<kZRj<Q_1gGc[24mkS3@FL`PI^DR`G@e;4`M
YGJV4`PNNje0OlR4^Y2V[WDCkg\c?AO^0dkVO`j8d9VFS8RR52G?IaeK7LnSBjA`
[JKM@Yf2ohce9l[02]mL3[>bagSP8bOhk147l8[aa7jZ70RE49[j>UmTdAbEjRBL
_\`Um@p6AI\oBV>j04A4Idl_J7Hf1:>j\[FWFT_?KZ_QF>Qin[EePM5?LJ:=ibM6
;]Xa<Li6`458^72ffF=FK369T\In@j6_B54gZT8^dS>n`Z^Xc[cBE@Y6]@9^j\Ji
mk7jG3aL3XY[C4<f]lS`m?:MW^VX=5G_e^QfSY1\g]6W6_=A5^KW_2Fp1o:6NWoZ
W`j3;4aBML\?<D51?nTGO?j^AlAkQ4daE<kOf?k=[[ifUZP<92Hl]YPV11PET567
a:K_abHc\>\Zj626E=5>nDjDoG8PjHMLc>>5G_\?9O[gMm4FY4Cd_Tkc4V?YanM8
a8AEN5JT\VFV`4][E?=:3oTL>k4_AS3fKemP5BaCpOO4eXbc@mG:ZKHE<[E?h`YP
:C\>fdQUV6:Ge34=2J9GRG1hNiBGekej5]G`JNPRUOL57;LNKgYhHOok5]U?c2kV
1O[c0aeUXbKFB3_n8AQAK3K]`IbfQ54g[35U:@^hofcM3b97\g\Hk>oiMV[hfW]O
oOTX8S:X\NJ>nHd<Y933\SFXPp3_HZ?MYVM8_<N\UOkI55:Vo8Dk5f<VGG7RCDdZ
2<Mif7odm?:F][Ha0VTK\d[1aZ3<E>dV]akKfFa59;g55e@>hL<S3M4FGb<C]91F
<RaUEl:QL9H:a7G4J?>YX3YKg7RO5PVF0SkUgUN0nTC`FVDT0W<4DcFC]TFT[iko
R8d<\FVnAYpbNR1hNUW\U4lf8DZKNa^PBOGE9jUmWPUIhF;`oo7V0ef\62oSb_?e
OLf2aP0K^g=b0]o_4NQ9L0=:jm8aeaBgZeJ6Jc7cPPN=^aND^PBVfgh8\2@RdU`P
Y4JQTI\ceOlJCP][18Q9e0;P?=a[cfo\SkG60W3QKmGkS<LAQE@V4?Z40MCpi]f7
Ud@@?<A5Q=`gO\KJ<MKHBW7LBKT6<3[GQV2M7Y]o3;RH^Xg?Wo<>=kSJPeeDic^K
cenn8k0UH@DVh6Ke@Ao3DZY3abTTl?I5XBj@8Ld1gVRNk@;?MjWkgeUlO]3f:=FC
NNYN8T2n?]QoBZ3Mc>WXDhNVF87BY3^MBk3?lD\JXSVQp5ZPVIhmRQOBS3Q1B6Sj
^:POF2Q5R]@4\U^l8MggolEE@AFekK74kko2RA>_UdWbN5KHSF\LNlkd;N5c>>Vj
^gaDo6j7fjX4b:_8nd;5Ske5`RWc>OI2>kCF>:?M4?9CC^lS<K[nZlL5ng]??N\F
G7;kS6mGC<S3ne:eiB[lYaL7?lPJ;phlXKn?nIa8[CnKYnGaPEJW`0oJJH4@?lVK
G40i7\S;81:Pg:L5h7TBl?MP=k:<F@h>2JE=j6\0Nj1bjL19PgVRi8dG7:8@?d>M
aS5GF?VnO<XDZI>No01d`<jM0i3GY\6J6oR=H:\Z>F;2Ko@LGhko:bdOa8X4MWON
Sj6McL\TL\E1OKpmARgG@DQ9iXMOYL71a^H0Rg@2mjmgQ:2q@n>J9`IfC^;Y^R]3
TKlMlkZb04?akSC;SX0a8e11Q]LW^I=D@nmMM7`UR_ADB19<@a3N[i@g^5CT;l[O
NKl^O3\>H67a@JC5L1i=On\YjhaCo_Y;E?X@U3Phj[1m\V9Gc[[[kngG^4_hROH[
Pk6\WZ\YH<g5PmjHm[FWaJ3Rj7990PU:pAg72_m@aEN>4EV8fO487g5:R?2nBH79
[To`gjO`bo<Sjm@0<a]AfD`2^6:hDNY[JAmH7TIBgUUmkmIXIUO80COc@Hf^7hS9
f7coNX:DOKKV6T>:iHBVVChg9Gc:61B?3`\1MNMBUU[jSBn85Kn3=1L\=H_OQll`
Ve`D`jcWl^NWlF3M@q<41O7[6ogKeJNP<]jG?BJM[oiT6c82QK>D6M9hWcmmgAYE
ZZ;]iNXUEZoIF2L5UR<5Aj`Onco\diOafZR^H\l63bdd`l74Q=^T;XG_OZ9USm3Y
FaUlDbBe5<8VJ@3YJa4nX^278Vo@gT65@KCSDKReWRd3_Bl<SL]kM:gU7NcLWQ]G
RbqZahER0X][0G_SMP5?T`>XLUXm7nV@JmeK`VK@]I402B?LcZ171m6`?P8Y2Vn0
>^YZDdZLg3_hV7mF]MAHhV17nhHm^>MX7m0Z3D1mNKZXK?L81H\aU0T:df<gY2V?
B=VMj0ea=<eh8QX3:hS9AYUbh@_mX1i6VodZ799h]Z[[ijLdjiHpE1?]OTcRK[fV
NVNk]DXYb?8_8Z8TG0P9jd^T_Q2gVkZbeGFLA>C_j=p`140\Oj<\MUK<c0VQ<eYh
eLf<K\@Da1m`hXB8a@aaFj<e7kS07bYT=jQ5i0V`FC?`:OLn]2>V\;F[XS?00ePi
3UX?f]QW^1H@L3@>nd;AiVLID>lZ0cC2EI[4`YXllKSP=^nYmG1V>B`PRMBkJFBD
ShK?@Ah]R@V>b431ZA4nR[Sd^Kjq8HFc:@i4[mJ?F7bmc_Ei``j?nZPdaXJBO=jM
kmZ^4Cl68RFZmHRZm=c2GJPMg3Kk8G<1O4HkGo_SY68OIcoE7KiI5FUb_jJPc@YG
T^KN9]lW1NR7gbLYKH9BAP8@eNoK6hAEb`UlGO8dclLJ5Bc]NOe05n_518aOH\nT
=?hX[<]hS4<Gpg1M`fUI4c7Ve1l:;nbHh2C`R_WO[oK0Vo\STlD9Ya<A?BEVa0`=
[cQ[g6[4]DJCdgXKAM7?F7Qh8^2?S:f?;22S14gZPOV0g4ooW4Sj;ZVBk_Co:@oe
2gBlKOgRE]2e4b;Pm`od27fHiTGeLcD3]kbi54DCbAd<]8Kfhn=eIYE^hXEmDq1]
RXSU>87aFAUB0P8JW>>hkno^YYQ>YQLab=8TM6=4CG\gW_^\CE\_MmOh1MEM<M1C
bY@ie=?]gIIO^OL7W;62F=a`L]9OYKeY>YlVM;AMkPDV8X>l?CMPRZEHGf:8Q^Kh
kO\DPD?W>`eYFh:lo7;Ue^aj`Q<d[NcQV1Jd[b:MJSOeG2pLIgE;:DXn6k43jbIZ
=lJC`k2GhR^\gJE_c\00b9NEUEM5<Y[N70<^=cDQ4d]G40gLj4^A[3`Z]CNP0_k3
GlgTZRD;D?:hIJG;=gC^Ol4hGaAEeQ?6RiOHKd^LiOMYP;37BE=E[5]ZITimnh[f
>adQGkF;_6U]4K_bTYcmohl^iinkROiq6PQ3A:a[\oZ@8LS`X1RTp]M=Aj[@X?i\
Pg0UL7l`O\JEfA@O0FDmb\[<KE8NebZ2CebT359EBRTH5IeP;;]:D]EE7f[i<T]8
b?[ahOkbK^CkS@:;hKLmZ;4aceVHBg;Ri=UZ6M>ZB>88?IUSdge2HDJd0S4@lTJ9
@B1_\2A4WE:4[@[TG_RI7KWC4W?_b7>4AT7BcpVJGWeiYL3VEfIe2g>^Oo9^gKjm
AA`m?fUR52IFd4cf\ieJ>DOKZ[TQPJ=`]:j?eYVEakjXi_>c_ZKQi]ObN:4<IOJ`
o4D8?:AnK6bQ4BO2bh6^P_Vdd7Lm6Kkf\aD7^XEnC1B4GV>_^jEUQm;>Qh@a>aJM
;L\VgUcmG[WV>Kbg:G]mOhqem07B5<:C;S3I]UKC70WRVT:>eGo^gHh_=[^X9i@A
74SN1_F9EeioSa:nji\Ffgde]lS:3C=`?T_M8B=_a0FNhHDSN7fc7HY>gTWKF>F9
1j_hAho5gDELhZULc_RSYL`4e0Ao5Lo`OgFnCo>43A^:j6ESSdWbC?B`F8I1o\WY
mSBJNo7q6Dj_kF]Cc:EGDANMR=7eoVk6Um^XV8OHkRnR>J_5KA9TQO5`^j9H_<CC
1\dG>fG:65T5`YoWG1VmQUXV_O7=dMOl7?_8GhOO[mD>O`N124=CWhCC3M9^hLKo
O7HdD^UAgHTF>G^iGFSma<XLheV[56fR7og\dVTkUdEUgAe2BlZc7DOHpeA_[^9U
nf6RHNHQQ1E?9H7Nh8Rk6;RnfEo[L1D69YRRYa1RRM\LbfZKl93`Q9L8le470EZg
nF]UN?b<;01?R:oAU^9<eT`nHHdoe881IUKf7DYgWF5_^GH<Jj]gV:UR3V4BA4:<
VF[Ba?O4HEEl3Rj?`^>Vgkmci^MO`bTSXXQU>KSW;ph8SG:_XQc@E<Dh4B;On]3<
Ub@f;1jOkfaQbAe33BX:D1TVUAeJWSOXVlnGCf;UdmhHDU8jULT77?MDK^JNL^<k
f28XHM]Bk[;\U\[[9;oL]>0@lY<S6Q2AECUO?;eZ01?bAUoc06TTn:]F0PgCHBMb
bK8VFR=5>A9Y:acah3_;DWS[cWpiDc=be\CNklIf9:1=<C[6c5jnbO=K?oBGn\if
;TN4DjlmVi182j4OH:iEDBcKf1Ei1[n?J\7GiCko:HSbjCnVP9C0ZNg@Lol@551d
V3]3_k4JD`74b]\A9V0j6[Hejnk`bSkB2QOGQ2SW@anRAHmbXD<0n:N3o9<`eDC:
RD:fCD[B6QdqJek7DA@LTcGoe]6SEbG`[PYIa?i;`S1<CE@bN4e:cbB3^cOFXXc9
AX84ZQOLEoTOJIUT:eGC`H4im;oVZZGT3GmlNVQ^]31SN\;jHGQ<Lm@TeNHQn>7A
T2<mW1O8kT?B@6GN7\^U`@Kj<Th9TQVIakoKN]U8?QhVQQ3J=dBSf4W:oTk?qdS>
B7g[Rmh<YV91009UeKDN0Td_0JjVJlDF][\]4R>IH=JFbbXj2k>ZK1WcIiZpW?H1
kDi;J@9WDgXQYmK;]\o=jXU:P0IgNWQ<0G@iXGcI9hTif]GR]LoY1UlaF=<6WlFW
Vka6bP8d]>CN^GKgYOecTM@:c0I7J;0_52f8HoE:`L2GTn_jRkhSQ6OVn>AlkfGC
oMSobl<gliWdlB\c[A@[TW6aC`]7BeSRd]1EPW9H^_D5p3oS:K:kVaSnTG=TG:_M
GFng4R2cP0B`;6lN[m3S26QSIZiAZB<N3];YV1Dc=09@d3fkJ27hVD5K@Hko=[bm
QFJpd<2:DHIiZI=ZB8:J`?0hh:lbBgAG\IgNDW1?FPD@`7VJbG0iG>1k5fj9b:]e
V<JlTCJBMVk1ID1RSH@H]DNNL<4a0[3JclCo4o1OXcQnJ=6fTlf_:P^S6oj0K5oY
KU;aN\QDA0lJqk\FaeE4e`:\oKE`c>:`KXAd;Yo>2KhP`i8?U\U=Z`71Wih5n9gl
\B3L2CXaFSU_o:E\Mc0c6aUc7;dNGJ2T`i^AVQ4lc6=nX:c?W_ng7k1P<`]8P?LE
lC0LL`d5AWF[BHU5d8<`kqX@\>mJ?Co`8QJJ7h@k[jS]_D[1foj6<Ib3\6FD[?[Z
;I<B8b96?OK3:X2Bg4X\INODW8HjTHAX01k;_932=R26G3la3m2k676B\?1A5Z34
6U9hg_5]Y9=oH1gh>7416:^[<e4L^jql?bR?JegXZA2CV29HSX1B^m`gBccE6B8U
Z[??1X_m2HmOA=4blVBSTe170F3L@Q8pgh62i36_ZPfP\EhJRc=I]aOleIC16Oh4
6P`d6T2COnU^B`Qd:A_@`LiU>V`4hl069W\c2kg;R_oO?Y5SX6?>cLUCVa\L[4IL
Z2`1^Qf=PM@egnRKNL<TkMiXJ9e;T]98WQLnCYcRqjMUNCCLnYZCYUdK95[44FQW
oh\Ie_b2UE?hA[Z@kCgB7T_WZa<STLgc`P\fF^T08?cK0HAKWWFUcFR=:aFJbOLE
]8mRoccMh7ehMT@09E9_?NJol]AK_1LId=K[P1jV[RM5X93\lp2jndmYkaCG17GF
U72mFARoZA;Plj=KPV2bl7>j<^JF0XUk:8obKZMhh5^hLk=`Fbj;B[:=6H<\?l`c
]k<PQl2Di2CQnI>2UGMFlb\2A4HWZPiKdK\84;<bhkGWJZmIYWDGFbcT>Iq6RADA
OCoaIQl\4N0fTodXITZKZl>2ImQV0>_GcfFhD1P[CmRJA\Sm8IRFI=fQ:d\IIYio
6MN?[D>9P>jU01<bYKgUgf4CXM:@[>g6LAMaNa0JjXOIEL]ej[P`VfN\l5[<Tij]
IK<p>R9NRic<iaG\C8?gNOeODg__`OWLj_Te5P4Hj?koZRMKSoFAK[CGIfjDfn5W
ienHmM>XN9aSM]T7]m92\am4cgC0^Al1mQKSVe4RoYUTA>\7QE0DhLIG<NA?c`N9
ZbYGTG=PAK]ZpeUPE9_E<jT??1hbh[7HdTh^TE]_k]\5nBT1_hB<MCAN<0MYH3l3
HOT0P@\U6oKJ;ZMONL5khEPBFgKK2?>EQIEQK4hDcqPR<K[odOZlc^l4NlF;dce?
BV:<S<JWo>GEA159Bb3>^Z3^5`<m5E`G<Zk1LOd7mTN9dYBQ\;5c6Moc5T_hH_X5
\WkYR]CED2jgAUhfHCaYO`HFhk8UZ8ga<\^j616fo^l6OS2i\[qjSnY_=m`Bj:IP
]IS8L<W]fh;44pCd9jc@Mi4j7ELk5W0T`KLk6J^9^C3CN5879ROR4FP[kHMi;n_A
3h0CdP=H4gGjFnc^hZ@h:JmlE9U\b@97fl3@aH[a]V\56YK;9n]PKc^O3l_H=[6@
J1EL11=OnVg[hYV073=XZ9pV?9UV<V<F]9cC4TQZe]aEGPbX:lh4>_M@P[5KANom
3Q]noTBeYPoDEL4h@bin1VIFADG5[mc7OEQObfh@7D^f`>3jPQUiGnRE<[4GOn2W
<K7gffd[@3e>XLgHGKJmW?e105Ik^TApXYGkh<7i;Fboi:j<89Ckm>;8OkGD1?=@
mMe<LiOo:c_UX6K78ZkoIYO1eU0?goPa`6C\aWmVPMUBm2]ZG6oPfkSdJgDZQZN7
?<eh=J9<[Kob_lODlJOh]K=`odIRZn_PXOf74K^?q[LKV0aA59GY8mj5`\T4[;YC
7kZ572I0Jbe2`8j@@7Z^`Wha<KC`<]KcYk?4god[EZ8JcmP>TccS`YkEAW?<ZZ2?
^m;ZBc\8`[n2nO8]^0>2eGfHCOONlKn3MNNoUl<f?XLHXDWW4q0LSSBW@Fb0YDQB
m?_TanfmSnlFC^3Zb;GXUfD1Wc?`7]5@eDL:l6RXNKSGB?o]O68VfbO5jHBQfKa`
oohEW<\ICb1n[D3Y3S78UeFL\_29A@4IEf^9Qmd9N?>=Y>K>4:7ld?0P5_p4n<`e
4<75H=J5O4Y;n3I>XfI[A2aeU[a866fd1cHD=;c6<eLgVDkQXcg]2MA2\k3Hm>jR
_KHF8RG3dP=mLMno4i_I]1`KHDTF46a=fNN_A_m`G3755<]iFcK:2Z6[ZEC_g3hX
G3;p:a49eEYFMmm_3^XX1<e@Z\P3co>1^6Y=5H3]a=XKG<X`@_9d[QgmI_^8o^Ro
?ZKLLW_INHg5`\>[jmLQTcckc_`^F47N=Jam=\3MM\50f\1jH@lMakj\\I=0CGm4
ZAj[P25D]VCTqHEgAQY3SKKB2J1[Pe:]F[YLkQ<0R1AIq:dOT1F_68lSUDamK\U]
E0?H?ATo4eZl2?0I<LledjQ0MkK5geGXWW>^P6:\1>R0DZU2hFU=ZfNMaJQdo23Y
@1=Y8P_\ip1m_]W@JNRi];EVWWj>>9XJCV:b>l8DgYB5G=KgMWeVj_C0<m`fKK;f
IdCo2=D0D?LbcGHjOVnh1j\jk33DW7^J1Klbfjh_^fA[GAACa_eOIaFCTJ83Q4O_
IJe<g3Dl[R9RJOBe^6qEl4ggIKGZIFN1=449^6GIZ\0deg=DQa=]IV>05<;V8PQ=
2[2BQ^:>5_2NjOTMfZZX;2APSjjm<mQ8^YDj^N_Z6dRnQGTccUYa[V9SN4\NgWjV
N_IHi=oC@D:gV^HA2l15dN^9ODeqRARnO2Xm\4`CNml@UZD7KA;bT0^0j:=4WU[I
f^iNK:h[YRAY5iZOo@ZELl`c7OFGa]lfj6_;am5IE[WnB2IHPe7]o4W>@U]CAf[^
Beg:KCPWZ[`R8URX:aZK]EN;1QNgLDdoHd7HpDf`D8E=?^oiLjcCZFNL0j^<lC_g
a8FBJb;jRJ]?blKRETfn3nT>`:0B9g]NSdT`?9K6gUIiG;=Pca<;6F5n6bnIXWQG
cKK<d?TjZY_W<lV=I^i=[_3AMQT:AeN[7@YYXSc2g:7H1pb7fJUfXFCMJOD87BF4
kk=iOfoPb:?8do\aQ>I;_F:_?T3i@NQONd0[^QPN65j0KcRaPY7FUa[o?ncK@I0=
MTk`oohTFEnem^mmQkn996:?R5JZNkO6hFAXbNHLCAU@[19Q9AjSH:pM7T;gm@KW
oOUH8o742nMj:dYG2IK9K64ERpZ5aHjZO=@>G7MiN6ToEZ`\K[52ACDam7djGBNQ
0M5ZH3NekL=g=M:=cVhB6DTaaO\5CL=WJLQK6Ln<QC;HQ_]g?iANPNc6@2MKGi\?
1SooYc;jn>Jm3:h]c^Dmb7_hoQFOF1?Y^np1nD1RnCRe=iB6cGDD^WTCjj[SCgFA
^0CDUm?PKP51BTH8m>Sa]L]AlQKB?>HEN3e0NSRFbI^F3iHll2kSh=ebT1bIP6ZI
kOeRnmVBc5\8ALQk4Y1<ZDU^_Q[mnaC<inIco3j[WnDpZ?3W?`Y\DeeCHOC=jOhf
KW2DVNR7k=Tg?efc;bKh3QW<CLBA`OmE>AQffQAa]96^o;H6T;eSl\UF<<<Sf`_^
ObdZhH0VW>I8<^fQS:lPgdl6lE\R^[YCBE@T:J8Kl=7UkBX]^F?nq@Ul\i<PWOg_
Nl]3GKW?`:V\LXZ6bRdScNk>0EPS:DR?IoWJRRNiDk:Wh3WbJJeRF9BP>YHEHQJo
:S^_TLQL9XYMP36f9p3geh^gqJ7;LS^n$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUXB4S(O, S0, S1, A, B, C, D, EB);
   reg flag; // Notifier flag
   output O;
   input S0, S1, A, B, C, D, EB;

//Function Block
`protected
eLbnYSQ:5DT^<`b]PN:G1c0B9hnEjngEWc[R\M_JobW5h9XYWe<f4JF=q1N;?Ffl
RCRdPk_a?lYF[3II;Y[VOjBC2Y2TZk4e2G5Up0ME[HHJb;E3]\mWW]VeL1al81_]
]EbVSLRBcd100q1bSKgTplcVA3m>DM><YWnBP]D?Oe973>8\kRjX5`6`TWeiAj23
SXkN;6Dmfd9_2FSWEjkK]R`pffY2m4ScHf4AYQbTo`:b:JfbbCqMC=m8B>0HlX3>
bJ>:68389>hMUR4MWAp=CBmMK9pBNDQKCplY6ZT59OlPZ2^<EYDemKWZZ2\=XGST
;QW`2JWDbIcS4ILd=_Fj>4NmoXQWa72FTHM_0K81QqP0b<bUS:TkD7I=d=WVBhn8
JG;6;W]W>L\YUimHj87fZ^EIL0E[DaU<N3FA;K^N`G6l39IZT>AEB2d5[7Dk;XMP
BUXYYCl`bc5>UDaE7<JKP=PZ`=1d34T<jaKickV01Zg1<baV7fpgV>?9_hFia73c
MAlNnOOlfeN6:k^`g]id1G\E6^_>3@65INgU=d``KlI;hMSKVLJMV;MQY3c8k>?h
?PgYiSKk1<an]X:Pal1`^GighOePI]N6D3?gmF7AilVZLg<BM;0nUNXaB6oqY3\S
A[T8Mghe6_4_4TjVmo_?>aRA2[=c[:6Q?_Rig9<KJUb?G<j4^BVMdi_lZ7_`4:^b
PLgf4BJ?W5HoEb8\BgCZaVCAVYKVL16\Y]ILJe@fEM`oB^2kXK3`FMQV8doS\80L
[3PnqFaRWCT@aa3dJi4H1XNP9@8h_I4J2ZhAaOI902:`ibKQQNQE;M;bDHZbPUPF
dGSUk;oeW2cWVKa\[YceQahP6<NLVC3oR<n24Vd9JM95BIE4gd6cHeTIEg_94Z>^
HPS_jJ:C9OZ:^q99hFSAj]32BYdXPDiocKWK?bMmljUHGX^@g]lD?efCK9U<EFCW
6Z6HcBaIZ]_JORARefHdOD0O:R_gd2BlScfmg1EZb_kLN^2?gP;C:m60SF_QPlUY
GWL?cKKg:I78B]nEmGZR9<qOH7OL8V7`3n>Dc2GE8^A9RmJ21__3hfUJXV<P=oYe
bL5[Un_Fh@E<\44ZR91qYX3WFMbWH6LKd=Pk=h?Mci3aC6O[@jBT>FPF2`RVX=@=
6f1LfdDULWSIdkKCRQF3lQAnIWNFOHW0JY34OkGKgjE5cmUCC1^l\>PBB^Ieie:f
c0LN8_eo2fSN<\gY[[<OBOK[FY`GqebR8AM0@A=TR?XMm:UNC80P3UWjQm]k6M?Y
8RElOVWbdAO@[c<iAcX5SdiPIC^g8\n=ChO31\\A>TUTM^8[[7^k7TmdIeYXVbPY
mT\@YRTFaZ9P5B3`X?Xgj]1;hYihKfBK>ZBiHpNb=Z]0UIXEWOZ>?_GE<j42@h@5
IcCI27Q<<h[GJ=UTG5_\3FP5fY<<H`7;P3]8RLV:91DU=:=g@\Elh^0klgCUEG=:
8[5EnePk<2LZ<QEac\THDF<4n`nNH;jG2lTachMN:lN<<VpJ\k_dmb^PfM6RKV5U
CgHT_cH0GcZg4Ff9[n7LQZX[=K:AF^G]Fio9_aZhi6nYiJS4G4]8FD;^PYOJDZQZ
_W6S>^FTHVCqAFWMOCf9;?i1PeRDDUn3S[[T?42^>P4Hj?_oPRU89AjSob>^XhYB
b3Ge54QcTGH]APV>Cf>4\lIm6B;`RRNH^]@em=PnP64P6_HbRi\n>V9KNLgM^6F=
k`c0?[Sf>ZXO49=RMiJ7\Afn0:CKKE4^PIT<:@QoP9K9q^P]B:W=B[gNl6IBb09J
EeODk9518WH:6GQ>=YB1>]8jS10IRZdPMY1YbNSJB4nSS^cLL5MLC^V5AJ1VGC8J
`\lTb[XXiKX:f55=745oC2:igKibU\9@WL02dgelJ3236@Zgm0YMY^2_S6PY8]2=
G916_CK6@K\KWp@1`?cUek;M>6X[KoD>g^]nD0B]IekU5gX1akQ29`n9TXGD4G5W
:`l_3`dTG>fmPN@FG>YbHGNIbcm\SRG96o[EZf<RF2Ya5BUR@gDjefHi2MaG^U\=
Jdc3[_Cgl=D3Q0Akh[;lh7NA`Kicc\mFon>Y0NLXV]Yk`3pR7ZW?Zgef_8ffVK5>
gbJZF:83V8I^iB7h@e\gGLhGf@LN6IWTJDOPVKJ;TN^a7Ip3OK`<US8P_KESJYAN
?XQfGHIf=9aDYT1dC<A5CD8nKk`bQe6^iR?4jEdUCWiG3>o3VcB^BjSc>nQ]OQl4
TYV6n0g?UKHHPT83XERAA>4FdWTJD?ZNTH2khicoibj>8DCR=B`8J3EcP7Q7L0;Y
f:mjJngiLVPH8hcq`hVcTmPWMgn4T?TFN5Ooag>Nf>CD5mE[cCm37lT0?L_K:`GL
Gj?8a>HIH@[H`o;X`?@QP>98DfDoVaXW:kW3If4Q_T1OnXEP=Ymcg^P2=<CMW?1b
l\KY;XLb>XZiSgE:C:LG@BCGD99YRRHK>;3P5JQJeAISnA71pY8b^n:0Si>4GM`D
m0do>nS6=bT=gLHI2og0=3UQToclW]?8?DTB[FTT:`S9GQdESYB6]2m_]b3X4P[n
ik4?`KIdNVSEfSAIi5mISm9dB>5DSMnona[5PMBgTXADI=:lNj`;]?Z<TbMIPc\P
OI^\UA=FN8l]nSn8SqJTBo3cAT:UDZ<lPbfeV\1[c@511SkOiE5T0@XClo7jVjUi
OU?C21GRaH6JU[bI1@J<WB@^<>W>BbG[AGM^7mVdE;E<BjdaibWY;BV1V1iE5Fck
ENHDmP`nDEbjn1BSV4WF31F5KgWj2=1ZX6IPIk4;:FLfd8d_2=p6L1hHPh@h]\5o
W=LN`T<[Vh=4;Wfk;i5;Q?n89]on3g`eCoE@00V:@2@fj\MM4Xd69^k2K1P>0hP<
c[jXhkXLmTbdMfKUJi4>h4Z`@`X>eMSF;7N\3B`CWYGI[l^Vb4kan3l8V>H>eSgJ
HZTU>C?1F\AlX<?USOQp5h@WLK;nd>MGU@`KR7Pe^3VdPCHa=Ag@0T^Q8`_^i0lK
^bAeFF@S@lnEF43Zc3aS55\@7?YP=4IS6E;:CE>B78WAe]Unh=g0P9VgOWMRX4eH
g9aHHmG=imHfP=L[Ffi3;DMQgabe=Y=oMCVfd59>[Gmh>ei?hhDeqcmU=CS25ZUT
eKJP::IcGUM]8i>Y0:O>4ZTe5ccN=haJ`7d>S26lC>KaULZM7oC]^ckYcHdNZPdB
IWC]Hen<D5BA5hTM[Z<>k?_d=gCoYH`PK^]:@cI]Y8BjZN1Id:=`QoXcn7M9EP^\
LW2;F>A5bZDf\EbL[Z91eq\ldYml6AFK]b\445=3dPN5AfYE0CKfA?>;;6Wj:6<b
T8??SNj1XF[K;;nWS`^X0c\?\kEkZWTZRceB]8[2Z[:6lfkSl]RCA1RcESekoj:?
M7E4=;OFiVSYHaDad;MiRD7>`\Xm;HT:0k6[XXbQ;d3]L\65oGR8dLpmb>jBMW3Z
CMPF1`REPUM`MPX1Y[g[T;n>M8Co1@dAIJ1a2RYSKU@XUGLBIa=iPG_mCB6>_XO8
fOPiSDIimA44jnJh4f`BR;A;k5E=?NdIgL[MP?;l36iMj1OE:LG]=2b>?IAV3?M8
lL@KY6TS<DPlKo2ofleB513p:3<i?H;1fImhBTq4[BGOZZgNc;0fj>5<VZT5VWe^
VHZ;G>0Bh`6gCALe8>eZRH8_AI59DaOmKHfZ9lH4lZLJ42P`cM4DXL^4oQB5hZ6V
F\6Lh>2B`Wh??g?_BmCcMf@8H`Li6^_?[2\^LFa^4Ke^Of0`gUTXJj>oXZiIim5\
TJ6LBYTp`O6hLlM36;1223?4LhnkX\n5:6[076YTBYg;XDk_4OjYAo1CZng`8SQj
Z;05ofSG`=_AT_==KF[DWn_YRQGnAU[NOS]lH5Y5?h9jV`:?56PX=<Ul:_K[QIel
DkCOJM812g?_gRd\KRY93S83>AYCVL800S@>H?WgpYAQWYAhYG^TK:2L_mAXeDac
IEB3JRiaeiSA:A5S^VlWN?]ZIH466Q53b\LeFgmR9YPKOZU_Fb1[GgXJoFZ;Ioa^
bI;4L_\akYZBZdNOVNnIMLH1`AZFGcK9U]GTJ@OaKlMB[[C7ObAcdk`2PT>11ZQD
^2g@W_H=ap[P[me=MomSdEQIXhC3mTFi94gV6;dkWcNNS=8V7el68KAO:Z2=]PaP
o69>Z_YT:A[aBdW:2=aXnLo4@AXI_AAOddL5f_h1WT9[gUkY?hM3KdZC1=L^U`5V
QOQ9F`Ua2]5^i3mGBaa2<=eN\S9B]4>1?PN1ZbhdThpg6BWNKiC6kMe5Mk>:m7H>
Q?58?l5Ac?INC^>AkP@mH;lj;S4j29>KY`1Ua6HO]c]gjl@WDNQ@Kl9RDill51kQ
np7]0O1[diVJ2AILf\0Q0=co^i3bRd0d;XUmJXIaUZBDIK@51CU[;oVdV3inX?=K
7?kjO9AUJ`<6@nR[LV_cDm3CXbNa`\[0N8DbJo0Nd7BXT9jAd=a?YV2D6Fd48jD8
ZV7_kLX73oX\@?RCP>Gkm<JQ32oG4cd5^\DXCTqcnPc[=\=8O5\J?M6lT>2nUmD:
I:Wf]@?aaB=H829PceTbcf9f?@LbPOnf]B00M_\6S[b^WfXgnF>=^BWjRF?J^LZY
I1><SfDc1PlY=fdJ\T[GP;NEah^8`;b4n^XZXaWPlETO:6He0He:jLijCY=7U7V;
5E6`NA:IGPoY\RBp5^OM^bN[7K\>[>J8l^R4jaB[4dEZDXKLUHVOTT@6_3a8dgDh
<k94?kb<K<iJ]Z;;KS2o]bG1@Gc9`FTocP:H]VWK<Nf4Zm_IL0VZ]\@8d?3UDTNC
??FPG?L\afoLE\o15K5MJI4C?CQ;`OA@@1nOGC5n;KVFCQ38LBoHp]2ofY6Z9\G8
<b`3Na9Jnlfb^XFehiJp3@hKk^o5OW;h7@UWF<:lWdZRkN@8aEPjH_@iY:PT^llY
>:93akP6mWEk[V?Tc[j3RV[@nbKkC\XVb^ldBF<^]VJIINO;\;7DKOF4Z@<F:HEc
\JPCo:EDeOHI>HI6ZmLhOTRU=H6K?KDVGY:CBW1\XlioN0f5NV8EZ?;;ZgT`q]D\
?97Eh6el>9V\nE\0^J\8R_E:H6QMYYMUfES4NcS;bM>]\bDK`mMKNW9>Z4kWTVjc
Y^LDZf9=jWOFUKlHgKf0Xb@k@2fOBUjUhnkLPP1gAEg@;Sk\kb8EVf8\m@3Jg]>8
o5C\o04HmWaL4YUiO?H\lOdGUZD8`U4M5q]>UOJ`FbIlFkV;g<nm`\Ke<P]EeQMl
P<\7dij6\Jl`h_D@;>6k<@`b]TlYT5]E_KDGc>TXeEdPlcjY:W8YQH9T=<IEeC;?
Yn9:iSN73X6KbOnjmWQ:kS<;LFAcPV^S<ZAmQ6K@fnV<S\^Pm[8dE@YDUF\>\8D3
?2=Za@N\nNqHEgMgH;25HkEPfAQf1@FNe]AXInS6;B=h]H`iC7^IE=eoRPAPE4bo
SlW[KoHqk1U>HTmO`[aX^^B[93AZm0M7U3\G1O[MR@JMY9]c9WSfa]4m3An:>E\d
TL2>P1TT1=d<X3ZCnbGaMThjhEek]IRB53?2CVm@GQ3^:c0LeYP8I65?n2a2il3P
nM5L``nb^4Hf0QC?Hl@BgoEkh0hXT0V37ACBT]XnXR3P:DaLph05gI`<REITO8PM
NR0AC\@ZJbD__;BFEJehk5IXaV??ZBBFjbhV\Lo1\hSAVeb:c?Dob;lJ4MOgUK7b
nnXi:XLm3UD:_85hcoPU_c<]e=KDL[]Id4^A6knhPW\aUhE\l_6jT>XC0[e>[3QJ
7nfOcQ@EeGJ=[1A3S`0e`cT;=qA98`E[Peo4l>@GoVddOAE88RB<`DiXhXiVhmN\
T_]I@J[15<i`HKDll51mc4@1bBIS>P70A><hh\gjNS2Q3\jGgNeFgK?bSWKQhM_5
X[HDY`FE\[DNCdFOdF7aYLPK^5Ad<?LHOj6`R5gJk\JjhOUjNgH9@A8ZhIKg;fp[
M8R9k\POG_3=@WJBiA3ojE6[n`XJRJVjobbJ;g?]dQ^kiVDQ`53X]FX2;EBS3a4e
8=jOaU`GF1m5=kN@nT1j^3?Sh1Eg4;]Acb`7dKDo08n>MlYUY?G<Z?RFYQ499NO[
AKl:MY:5@[D51D[=i\O8OAd`O4ZW9<GAPmRqW6@eG>Yf][k<je>EX<SOXJ792oga
AKLN13\;K=Ke6L]X``HfYbd4kOM0a8\OFOF`R5>\lefeBne3`7@`HIL:@PHZgHa9
hl4<D6\P\3cA^[^iA6^aT@IOeJkYLl0BRUf7WV<NNiKOgkT1``3SnZ7Vnonf`nXQ
A]\?D;\Kp0UEch>e@9hSX[AlTWl:E6X=JV:W_JEoclI<::]X?mQXSY@oUK4B?0?d
eD\\;OAA>A\@kkBDa`SDenZP;=hL?Va98H:W[c[`k1m<?FU933NhYh2ei>A[A_L\
9NAo5cmKP_cWkQf\0M;U:FfdC=Ab?6m\WlT8RTnSMYhjQFALMpRUAIlCh@glVXZX
ZLNXdZiNk\BL`SV?lc<7VJIRNO\kUl7h<1kF:04B520d1:`g3b[XBVS<e?KZdaLl
Rel7bG8kkSH>lcl<;:f;VNn7R]ZRiKN=mZFmFk<M^SKDON<QD4RiY1PLPA\^b[L]
?UCoc>mc1kBF:M[`QhfGO7q_VDk?Ibe>;A=k8<KW94JS;1gHQIkj_e;_C32?AGjI
d`XI6gB5C6QJKUSH^JDL?GEb5AWNk?53iJd^B:1o3_@F^Ak>l2HDfjYG43FI]jXF
RoSQ>j:0d6HTl1SP<<[HoaV_6PnjT;3XmRH^IE1B?B7jRbjFk12;=FVG5LAqaXXj
Y^M;F:<Ej0WePjE1F\@XU11GU8MV18CbNbp9?Z0M?;^biIJ^9N8O3Nn;kng<jh=O
E1X5>LMXUWJZ]g36W7Z7jBW2cG_M5aCcC;X7QKe?KR];j?_BgW5H7^k1;g9]jU=m
goaPUSLn@2\M6fU^=`HCR28W>KlMa742;DRB49HedkUc=Tmde;SHWDjFPlcFMPTH
95RD;iRnd7Rqm\kRMAXng_ZW1kTT<hKWF?:G5^<@A1iboM3jjg@cDZ8TD6`NlTAH
Vei?]dSghE;_BeM>m^BUDE?\l>bnXYJ_fldIX^5X\?5[:nIiD5>NLA;K`GIF4Elj
OS`]Q1E`2m0_lLmO@8h;PH]DQiJJXoAAA?=0Z0`_PR1H7b;iDUk:q0kcm14VA;4k
m^7IAhPdV1:1U5b2c4KYZckkSdQkCd@NNhbdk6OdG^94ZE?JnM][E]\CcMOC0BSa
JB?]mI>\h<85F5:52=ip@JJBm;H:Ri^GhJ8Uhk0MmW>AXnC1JK?C?_:gYE<`G9D]
:fmSP0iOUR\RK;<LmfNj@EVKhRk<nWNEoZ2[e?c?:A7]AR0Mon?0n[\<YmNfGY>>
7==0Ead7h<fnKj0FLbj6XUXfRQ0\nme^Pl^;j9mK^`igAgOMX6<G?2A@;1LMkcEV
`B1@qC<EaVb8D=kH>o@FLVKP7U@61<_;;NS6\3lE9qKcadIB6<dWc26_VjfQ;hgG
iZ0G0\Y74]RWXHQb9E0gnGR^UU\VZY5`:BQncd[7TMKeSB@bE5NK=8<`[XL6MYV]
n6OMU6G_4]B?Ih@R_7YPJPJ[<E]C1V[kn6?^W=fSQ=X7MZh^gmNFPn^cOb6Di>kQ
]^OO6:3Le^hAeMXQQg0_CLMje2p1@FJVKkN0d5PCX<H?G6oHDQH7]>;4:]\5Sb?X
QSnJMYAUk^F;JK7fmKe44CZQS1A1`3YDjM5@XB`eH^Q9QTPkIi?^RA6_j]QXeQJE
6?M]EO;5cQBoiY\@aDf3OCHE\N>ciLfD<@\@be8g0dCkJWmDfKV^YP3fN:lJm4fC
iFdmgo:[E9op>??m6D=IPdET@RY@_maa=0HOXEJkTbd]9=^@;e;cc1?:KAgTMFV6
U]Ze;_@08SlQ>]46U@gROUbe<O0c?JQRYg^hN=b`=bd1>;bE8A]AkoOkG_T_LO0A
\03\LQdQ^5LVK`M>m6m>OLo4^iYIce:O53:dN3AOCBjCbcKL:WUIcJhLf_7ZpBoD
DX:Zj5Hb:45DCXZ@[0B0:SUY5UMX6MIiLm4Ia`HB^Wa]]jEh:JOG^b`\QJ`UMB]X
hdR]Z0l\e_e_c;CSXmoNQW05HRLXW\Q8nn9Yn;QX80WE@nQ70KkN29Mi`\oIY0gP
aiVJ80k2I;oNFO^<c6liHW;kN;04C^]5iHPY>QXE3o;RBq<O[>dN5IkhoVbgThno
L3BNbV[Om5PJ]3[]ZhK?K`e>k>]:\J_KlF@jRg[=@bdG]L<DWb=m_iFiQUl8139_
?F?NmR9BegMT]OiXObA095dKT1^MM]LDOT`EUZ3eAJBBc`T^[M`djeFeg=;4V?Zn
nKR3nL9UJE9GNI@aT<S@A80OVc>>KTq6R6?3Fk2SN`Y2<<:jcJnFG=g_o9MY\MH[
lIJ<B;qk:GemN^SlK?[=B5ko\kP=gTaoJH43cN8dAUcE\fVcE3jol?mF\c2i5^>E
X5TR?>HkndNf8[[;]TGV>T0=5P?G\oSXh4SW\Nn^^M\OM]i39J7eXLbXKA[WUoZJ
WkEh3o;cX6K`c`U;0\[jSI_N^3>8_U\XW=@XOMQG9?IWhc4G[KLSlWap90MDLJ=e
PZX_K=hCB2WihV8hY3b43g?ROFK05ibXH6enHFJeYGiBXi:a=Ylg4dKC9im]E\9C
>Jf[8JLmW6Vio:2ZLoc\9M?iJXOj:M`=ICdeFbZMC]UGa=@TeUL6cR_SIkM;`c`N
>fAn9OjmMJ2_X3fTLIVNakO^@dMB72h1O=La3\5@pl90L`H_K0a\BOc09C[h7BP]
=0[_6\VNLXIZ?@bVGk6Mmh1dCaAfBB=X;hYNCjSWFl;[PVo?Wl\DdoQhDF>fP:oX
gY?c`hTN6TD<D6M4H=_DM8BC22KW?IQN_DXEU5LW=5C7JCleElhf4LVE4YocEfA2
MYoi7WAQViJM`C>9SAWK4`J16qZ`QJcU>7o@:6=nk=:;UA4Djl;Ei^d2]VA>YWJm
;mIm@URBi:S<>WU_b_cen=;?L]Z>a>jRn=@dGW?8DRB0<XMCZHBi5?7`]bOfAVo=
3=:]kaGbPRlMJ6ceOFoY<ERjFnVP9C0iNB@Lol@G51dV3]BPARBUO2T9g3S[LG]D
maKfLWi[XAp;2YJP:R9Da6?]D<f6@jCCSg`L@U2SoHOEAhc\YU3H7[VK>X6;GdKM
WRGAfj6B_^4;5[0R]Rg07K[]@K9\eFV_]KcH]b7A9H[6N?hR<LK7EdWC9hjcB3gK
6EYECa[IBGS1DL>?5PE0X3_3\m`G=BnSn@IHP=jiAb^YXgiBcnPmVcN@o93pR172
MUjlalNHAWS:62eO;O:D]MM=oRlL[ODl\fn_fM:WHYgMcmaTGnLXgO=3\F2^R=W9
1]PcWR`\N>Bn=Kg_bXhOGN?jA5lFoO0mgnBD[e6d?KWZlaMPd`[_M26WnJBeKUFn
GZR?Wd^OCJdeN?>nn;21G4W:hC14@ER^OV_AJoeC60e2q6L1hHQm\hh\GoWfL4`N
W[Vh=l8WaD;i4;Q?n59e`n3g`ePonh00H:@_Lf^\iM4Xd69^k2K1P>Dn6<c[jXhk
XLmTbdMfKUJi4>04H`@`X>eMSF;7Nd3BhCWYGI[l^Vb4kan3l8V>H>eSgJRZ2U>C
?WF\hd[2en[0?ST_0TmQMnX4DWFjBp_oT\_m8bkjRjJYmP\Mb;A?[g:mBZ_2]ODm
FL4oZV0nfa0D70EZX4Y^LXm2pPTT_mCCB81XO^KY3RaOiHG=<^Q_Q?F`n;9fhmf]
4ldlbm@3O46Q9PifiEK<c<AB8P9X=kW`8fC`jjY70WaSJ<`3DKmo1>V`Z`RT6N`a
4gXkEOfBFMJaFB469Kbog;];^;\TXGMZ5f^fDFh@HB3Nb8dZ6K2bgIo^jA5<E@aK
lc;EYgc2AqldOP@85e25\iG[@DhFVLiMUJ01:i[UP=H=JZga3Og7S`]X;Wj[Fa\<
hn\@M5:k36ld3lEU2XIBcGD>eJg9kM;El4Ia@B@mPCo`7UIKbR;C6B>_^L23POad
EJnm8N@NVJ<kYJ0Q=?I^;8^XDBP86jTmeNI_^UdQn=VYgk>Man1;Jel?gBqSR]ac
5Z7Cfefb6^:FgO_O::gTd2LI2iQNhJ8]8<:7g`N?JS^k^WGLaRobB>ddPTkS>TUf
2<cA9dn6MUP?aKf4O3\m=d;i7iAB?J3:^027\FiJ>g<cdY[gDEM52KWVjHaf`NjC
E5HA]76XR0n831aZ:aDm\82UeblgcjWm?<7o3B^0QR`pO>G4FW?TlaL<C13jn\\C
eFV^<]`VS4djfYjb5G`IZMHW=WeDPaXY42MH:>\;NG@VO08X`LXA=ChK:P1[ao8N
Ak0Pfk6nhTd:e;fNlFW;FKS;Kg6Wh^f_fB`CSDmn3LW]OLQl[g]f=iDhJko<dA8h
BWGUf^b>DTQ`Eh3j=PG\E6>k`QgNqSnDFFXdf8DgXFEA6G^egn`XLD;FUGDd9NGO
D5GQblB<mM6T`]NjcFcT<^A[18L1kSC4oJdb>?H[gbTJX=3fU::jV_L8:H4d9PHb
We0Bgo8P6=[FfZ5Xd8085Bg@DA64MGdk8TI8O?7Oa[GL_\d[b7m70_:^L8PPEnk4
[ln3@PMnf3J[ipi<9Z:i]JnePLoBhG@2ST4NAbkk>`AgGai?\hf9^L1oB5qJYfJ1
PiCc\J7Y:dnQ:AjQ8?`MPYnW4h0<>9]\Z78PULI8T33To:ANB@fXj4COaidJ3EiA
GQ<9eEXEiT60;4oHh3GW`kf]YhHlgW=2a2mmM>n>UBL5JWEaBSCgVdb;HWYEP=gg
3kV9^o=g9hhmAM]:5VDWPSk7oS0SeUQ9FLDCEX@j^2EqK_[T;;Xb[k[^K[`mbTnd
H0=MMSG5H@aV3X97EC<]W]@9TjKoUhe9SHA0:CaZ^[UEKFLT66WTF1dG_4U=POZY
<1J>62>\@8a8WZH3:Bfn<dn<H^3<eRXfC[cS=Zk6P`_[9Tf34EB4F_6O=PeAZ9]<
49?C6I;=V0=:a4Da[TjShJ551I=CqG<817]M`C<_;?Jff1H]c6nR=U[eUBNc5m95
5BSd_[MEY=HlAJ[o05h;nmnk_hW]>GH>[=ITRDiTjD?:1AP9MDMdb<R2@Qfco;2a
2NkkC:NB2NkUU8Zh<7PemVS`aKN?\]Of2<S]fD0]jAOP8YomI:On\<dO?CaddB]R
6omU`aeQJOM2Eq8Gm^i390HS2ikOE=m@AePe5DL:4[K5;EeeC6`D<:NGibNO=P0`
oA:ob180I6_>X]8P59W0Y[P1g?^3]k_C?n?W:oH<3LVK;GC=f7jZ6>0T8CM8WZ`c
NnfWgUDKIRlYmBl<YDLZULPnHUZ0UVJ5aRMmQPH^cX3gaCBlocFM37Rd2ZLaA9p3
bPZXK2;N_nK_>:S5c:eHHmn6nSh:FZIm<5La2WA@_:nCG2?SE<PJEcQ_i_W9E<<3
YMENS:5H^=Z\6]Q9Th?L7lWaHFl^5ZF7Ol]F7JbP[RnX[XNUH\E]I:N?]Be85YDA
3@0N:E@HG4bmheKl:`VU8a[aQTlX5jnIWV^C2HFR^jOo77UpVATYOLN<Gj4:[05Y
R<=J[i9oMSPoQ5R8@AX6nOKPj=o<Ymmd\R[RUC>JD]TdaPmSVEGcjE]_]E\[3_[9
1;R`C=djH@d;c[R@iPbg<36XW?<SOSbEn2Zc]4Q]UWdAF0RkHkFWMo6>]:KG2W^n
>ZmUBi_?HMf7@2TU]LJ^Q6hoF`iPPGXIqMXhJDOl4<CC7AQ`YZb15U57;ikUliTW
lGUOefgY6gNiYLI75<H]69NBFKS^lP6a5MSXNGE>PSXX7nRZGYE<=gK<KdG<oFTW
2Tl056KhEJ2=XXGSG<7:ocLiP_8jOan<n7e<ToBd>S5>nNIF1ULQVPEeadLXVcX2
`o:Ih1Ii`@MScRWdgp`CCR1@2Z`Oi`Be]1Z<fQc4cBB10E:A:D]eE5W62TkhTe^B
k\>>\62IF79M=;J:H:`0M6O\G9j<G2hLEKEZ28Pm8:0P1Sd6:F6mA6>@3BBGM75O
U[bR:o2MJmiDZ1\=FKE1ZA:I1Bj61C347kc1`UYXj70V5oUQW2EWR5eiQ8n1>dmM
_Pq1Ul`\cWZWMY7Okq`0W[DmaHfN8`K1JlSf[@eklZnmnSb<B036i4aa\4[^eU7K
TQ^Z[1Sjg82YfgDR0S`@\SD@UbO@:]iKW\YUM=;8o3mR4a0]B4kR;1fIQ]Mh7:]F
LN]N;3Uob\EU>kgR^Z0VhUU>kgOZeWQ03o4A56\lP_m3E0]cc:mb<3<jYZQo[lWD
afpNXO\FV_m^lePP5KD=^2BmWkjlnL[1c>ZE`\ZeVc4HGCX5`4YWXiG80?^k:d;D
>64NY@SVhD3:5m3XURI3][I3naMRUm]cO>PP;5??5WCckgCkMdJJWKm87B>K?fkV
XO]Q5<CK6\V:?20J?PV1ToK2C0lRVPGe`g``_2ZO<9`fiUoX\Q8pSnDFFXdf8DgX
FEA6G^egn`XLD;FUGDd9NGOD5GQblB<mM6T`]NjcFcT<^A[18L1kSC4oJdb>?H[g
bTJX=3fU::jV_L8:H4d9PHbWe0Bgo8P6=[Ff55Xd8085Bg@DA64MGdk8TI8O?7Oa
[GL_\d[b7m70_:^L8PPEnk4[ln3@PMnf3P[:qo3bS>]MH8N^On]@<o\AKgg;i:Rk
I8I]ZeD;=CXlHlaoGiEAHR7705e_:O338bLMlo^d`aX7`aUc:cCGK=H[[4\INf2C
B3T]5GB8HCP?C?bGe<[1SBgnlmRi8??I7O9m]>_9eY=1QaOWKT_jI`ff9fTe<f`H
]5m<A7P]a8oGDH:`?4M\XqS68Z?WW_cO:FF^SjnVX9W[MilZMD90[S\IbMF8Ed@D
Uad\PlU3Nb^6SlJS;F>NPLSbiF:m`f>kgFeP<j@]4Dk40LhZdH]c[YKT<A4To0RQ
C5_cY0c_OKH;?\nZWd=iKUhjW4lIV=>\mBCi=]F6930Wi>hIeiK27M]^GjNN;Iim
E90\7epk<3^G0:N>i@Hk^XH0S0;2PliW[C?`4TPScd@WlGm\LNIO@=4cUPSYoMZi
JB8bMUDkTg[^\SAJ@^0^<]Ib?O6`PZ;jWM`OUT]Al@cc=LI<DkS`<89:7[k7>LN\
A1`POP9^\35E=[UJ]g808Vl[K@a^`eJjoYm1A>EJQEm3ii:b<H9S`4DpVZ6\RTc<
:=:?OARVOekh<@C_NH8\_1m;BdG7e4_=>`qQk1k:j2Ze:D?\NRel0lPRUA5ORZ`>
cm\TZ0lC8\f_E0l4Ab7FaCHHW:W<LIWbbj<QmOk1]m>S[?@da_U6NEHa<p`c7^;Z
?O9DhWG;:64\73Ki664]eL6ETcPS6W5R5iJ3onOFkZ9C2V4MZ>ncK0bhkQ=79KEZ
?=h49N6f<`2RS_64A:CAEXOk8MQQ6H8J1XA8CdTZZ^?<i\UcZKE:L30lB]<UJ11K
O0pMEd1NLmfZPjU4o1@HN7GkOZSPlGoFCk_A?\\3@SLN_l@VhYBb8k>5<h5fMWUW
1dd<P60]mM=\fiWYgfl[5TF:@go9Y^\f4@Mbf\6]Ej_oPPkJk6>\`=eZYh6=G]MA
81YZf=A\O]Hq[RC40\nj3W1Bo7GL\^86jgI>QfimnV9Iq`@RP3j<Y\lO0P0eZU32
;ETLUW9SM`n5aO;M<6f_9OGWXGbLnTFnH?c_B9N:XNh0IKobYjRfce?j[R9K7eTD
IGeb:9o]5Di2]nLMSiZ_[GX<5k6eHd:aQ\di11l2F5_WME4E2cM2gp@4<]dBDMVB
b\@GjE9XLR6?b5iGFZMC]Lg;U@^YigEW?=IPo3DO<VKS1dK[HB[6T=CF;\XGlEM]
kThE84W]VYceA<2SN?W]LQlPU`18ALkFgSM\jn4YRCmg1BkaTF:dOB_bHNTTV\pj
:HDKL9:^JWX31KE`i3leS6d[>C^Zd;6V2S_S]Q`_[?6@Z@SMHDmZ@aCflA5E`0WX
70Q9QGaP0N1;m`fU`0o:\NW6LTh`E]]`ZS6eI^ZcbY4VVoNHU^Wh8<[Oj4T3;EQ9
1C[Og`DqeEKHUMm?9@QLK8M9XAO5a63WGLA6N1U2UIG@H5mG24SYC8[nAjB`aDQl
\4N01No6<ITZWlUNC;iV7LfJC^IOS@BJUTYm\JA0?^G4>V=fQL`GWT_je6cm??Qi
;P>fUa1ZbYhl90NcpC51eg4`g5[:Zg[EZ<H^8lbNNZa4X768FohDRnNJOp`=YVUf
Y_V8;2elBgOA2MPSLB5niP@Y]=9@XSaU\Nkf:<XH2lPSk>?E:8AF[>fWKON9:SXF
Wh4D:XDW=>;?NeW_aPO;\o:4CZZLXd5gGK_l`X9ANSDBiCkYY<dD3fJ2D<Lk^4LC
JWp:c01DNCgH9jGW>TXI5_jH[oh[7_M`m@d[i1Ql5Bkd?9dgihH=@@\N9<EcaA^<
a[^ZG0GGgTj:R3YmJWVTQMYhUdBHJF^C`KH]>1PA`;3ePLHYf:]LfZT_f7cg0n85
@0f7c<W\c<gp<Z\ocdo;0;?bPN3NVgI1O@IS8=]CgHf`L?KoEld>WkMSo3XSiISL
RS=XkZC@F1Fm6M?Yk\DD:NRcLJoVUT@QUQ2B4VdZpmBFf0Tg0h_3aC]g3X93A06h
;?9A9kdi3[fno>NLc_4Dg`hG7Cn::dKic03D`Dc=VdLG90`<V1OJEED4V4JXM;=J
1\Gng4_c_L4nJVXB96ZO8TTZKIKb;LPia?BQPABnTGnjdcEWTph]FQAaUmd1^8g@
=oQ6L;\IVL3Vh?:j2NZelM?F[:V?DoCYhEWEIn0W;BQUBSUCC4i`n]:hWU6dR>dW
0ebGJ8IXkoi\U8XZ:@YKl5Ga]iaC51il?9;gYo8=7O^e>BC>mfDEi_iG\dp[dmN>
;1U`?dRBF@A7H_FfiHh3j]n]heN9mCLK8MJc>M_JRLL`Ck867_:eD\Sa_j>dd0dF
PU>>;<;\f=a[2R6XG56I_XAOgA64NCN<LhVc1gl>>>ENlb9R<_Zk\32dBlnQaClk
0HRp[bBQg63kg3_N]PoRDjLHFm6WkfH2YSkb7@HVBb=17YK8JYDnakC<:N>m@7KT
RLYEMagk>I2;17ZHO60>4R<GU9ZD6UP`^5_157HLFZ1f<Tac8Vmfb=9>3XV9RPSF
3id4Sf?K>O5>q`AN67^Q1:CRfc6U<eRoh_[E64`X:PEpWoQLX==VF7f0o<LOAPWV
CZ^3\]A57JhUVe2Vdo0LdfSiG_YXm0G@fYD]Pj2gV>`4nBL1UYO9BB221d=2TefX
<i]l0iQaP7e4462R[9D09E6Yb3_nYPRoA6@ebmM;JSLOOE68J^EcpWMRN5C7dDfj
H[0J]0^iOHEZG10\H87=2l61a]P:Hjm:TNaccF6V1eng;I[38CGe`C`TETn03JDU
dnW72Ke95=CM\H`^9E59RVR11I6=?_hIg7h8DP8:84@gSRcf`N6C8LKlN5[=Opl\
@HD[<JJ;d4<BYe;B7<lIQm:bo`@]=n0nP>KSYihNF[V23AniB?UZNNSO>UjXl@;D
MiU@NUdF<Y5G;d2lN>PlY<X=FVOl><?QPERnPeMPD2V>k<7^H^SANf<[XQ3hjW=G
\15H21pBTTni;bUTaNDj6KA\alESZD\JAfX2PSjPWMd0oN8?Mo@6Sn81`fG_GNX4
B_VL57_L^[]X2CGA9DjkajVL1Zjb89mD@aChj<5k2MTGGAooSDb7<SmhGRYo\ilS
D>^i`2;K9nJFO2cqfTn3LoGQ7Y5KlQc<7[cVoDQZ:fFTgJa[K7j<i]_C;YCgn03j
TNH9c3i_Po\[VOjM6lR4S`BA1XX>J>K<X20N3@YkiX_Qp[G\_m0;P_3Gi]ZMgDa3
64I0@k=e;N6_d18FU<`<1F6TncST<M?ah6T<]k4C6`^WDj\;q=_aobBMc583c]03
1cikOTejhF^0H5^7?UQb\TViZ1^RF0\jFdA:ZI<0P?;U^Nm@h8@Gl9@KRd8QdN0S
gSF^2]j:UfoXj@:a\Jobj:\SDN1;CU73X4Q9R:90ZRODA<3o`_dN=BV1>pSbhYW_
T]h=oC:e:55d[IThIC8LO0Yka9BhUY]^ZIn;9bIdJ1Mm[3WWK?ED[`1f<^`ka\\O
<<?T_VX^B\?bb8ThO>6NaYaWXRFeUKBYj:ejnH2]^UPhVKBJ9]9aBZJLPF_V`OZo
F@qU@4Ek\T^`DmeU4=CN8d6^8V8F6T_EeRWGLhXL7o5Q0;<DPSQ3QX]S`lTl`PP1
6I8l?Pa8;HCRO2mlhJ36B;PU76C0k\WNG8XAFhU4XT?Z5c<iJdY^nQLB;lYZGAU<
iDA>CWUjnm8ql?H6:N63:5=S@dHE4DPDUFFSX;@mFn6:c1>5;f0I9FFE38BWdJA7
Gi=HYE6DYPFCX5@6TF>H0;HUoYPZ6M33^Lj^I1E9Sf320P>a=fGj\TZjP;LhahIL
`;^Gn^O4X7GRokMaWdE3pd`RAlMZM58LXWVgQfhD_dAT`Y;?c:[W[gQVHnRZ73I?
2W@iqMWRD\O?cPHIL_1l9Vbn4cjEPh:j^EeWg[M4:geGh6QQL8bdKQRH7?ZhM9F1
h]DJK4==>bZ1UFeoETb=DbPcjk2?Vm@7=UkWa`W4=;G8H=;M2nnH`\Lo5G:cT23X
;KPWVBX7I@1e:pSLhO;I3gc8DQ6D7<C;1W[83J3I^o7Ao;K7436nZ\YVkOYNl?8o
WcO:;UTARK@YTJ;nl9J^=;]H:m@HTU?4cLCLL;QUo8Y_1b6647CVcfNK9kLJGB@Q
]YeJ;6d5P<WWnle=;KP7AZqkc>J@<c@TMH_ln:MeNiBk5D4VW>C@B1P1WJT9lmPA
[5[V>fNL6:Loc39NLcBmN[jXk3Kni69\==Z=B1F7B96FdE1C0`P1IHRI0J6TbWB]
?6SOCkLkbnE2A3?`\fCKSkj3\V?<:N1qe1`=ObO`HNU^_McUKmN324j5Jh:T=K9A
0<J`acZZiE2=a5E<Kc14BliHln93NWOQj_0]klH>Pk=<XWSio^gMnCL=K]1l?<\E
1BJR6\N?^K58?PD3b3=UHWf1UJ^0jUogUP^7d:SipiZlDM2h7[904eAAKGI9KJaU
6_^kHPR:`VCRoTSKGo4T_TeJ4ECACigBL@_VBH1=;oQnAfifMMmb70jAikKmF`7O
TGc;DqfPgB>`qGD49TB1$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MUXB4T(O, S0, S1, A, B, C, D, EB);
   reg flag; // Notifier flag
   output O;
   input S0, S1, A, B, C, D, EB;

//Function Block
`protected
[;ILESQH5DT^<6LaX6NJhQXdR\7aRb]0k^Mg[eLCi>@47EE1H=HH]:?kdRVh0<En
^aNI7AqU[4kb0dOD5j@Ah:gei`_hmc;GdZZE0BhXVg^jUmpNJZ3GkQ_TG`IUo61T
L2gL?qmkg]?6qP2afo0Id]lO4Y>NgP[mb>IF<<KnV2R<PlYa9]j9`QQ2VWo5:@aZ
XkT5Q2MWZ3m`4mnq1RRcPg^C;KeC\Aef2a=fD7R5?dpT_dcD;7lSQ?`=<Z?^^<Ta
eiE`ee?K>iqkDE4bIJ5FD6YXb^AE5nK><hjbWAnX8gpOfF=>\IqX?WDXlpid<58N
egB_`8LBbP;@MnoIV;<\;i43LWSnKI]<X2mI6YE<HmLGM]0n:JncUKXYZLa<GZZL
J6ec^QJGeZhC@YGGWW_`KHZ4i8^=K><][gfJo62XT617^nAkS4X:J<8Onk`f=d^G
Wlp[YPQAGSC6:c4[I[LCJFG5<4DLi0<cBg4Q2Cm390NNJl@DJ001dgPQoXlDQ;W8
@CO^oUfm<I_ICI9jYPm]=\c@\4G8E6Emc57BBCi<V[Tk=3PcUf@o11NGMXfIPH^6
`?ke0DE5kLGp6lWE`7MmhkXh2g^X;SB[bWFdn@5MQV>V@]KUO[e3N]@EE[X62C\[
Xm08hC<k1l4Cn;CTAQk<@N1DBn0M]1JM8SRaGg04TW45`mKK<;d6_<NW:@h?WMXA
m2ZBCIg3GX8D^_LbVc]jq0=UWXGU7om@oEodHN1[61al?7X0ZL37HocoU]7`ZG5C
YRe6gcF_oj<39=9FmDgVJW3ZfA4nbdD]Z8mcCL[05?Zg^8<a>kL^i1SoB;Q8;6c?
bkN:4d>7ANc@6k@2<KXH`oTk;l<]gpUD2>NHiE:IF<S8jGS`W9L=k=g_8LgUZZXR
g3n@0:610_b^<hcg\FI4[3XJ7k2DQl<70`lVfBOdk`Xej:N_24[Wko_^?b:l@3Qc
g`3D1e`D2l1IaZX?V\J`[QWZ?:ei;CZZA\aOJfqVO7Gh=J6XJckD`g2iQV=]C0F:
`F]J;EneC<M`hK1AGn@hXbcD_P?S;2;F[dnm<^oQm9XfhZZIIVfdE>XIPZ8CZ7E2
f?<<ZgCgQ<]YDO[OGRUgBOC^n3V112A03;a`BSQf]da6?nhpg4hWnFZMRH1F3bKi
VijX^HRgo:gBM_gll^DfRbNSiDp][9ToOH92eH>8Z30?N`7mVDm_FWLd?]MSLPRD
9d13U`7RS5LU0GPYY3:e3:0FdZ:D_P00<HW5JMOjMG01YSYGdJL9dGC8DkViRP^A
72G]o?JJ7<Dn2;3CRPD7kJ6`G>BSS[V`_4op<@iK\6C\HfC`]GHGMW1??1YQef]Z
`j6T:=80h62N;[KhQVnHh?af\\e:Q=mSfVHlkY=Wo8bdCL[ibP7LQkn>Knf73H\Q
IXZHCc8I8804QZm0ck7A`c^D7HeYW=gibRLM^Ad[GTfQp`aVh9PKbkT??h9eX?TC
4EZ\hbb?W;W8RQh?hIgcH^6fM9Jd4]HD]C9Tkd=?_5`^0Z:d2nXN0W_ZL?ibSbK:
77[CnVBDXp@HFL>e?ok<[GR]O:OUoBRW29jcZ[a9`f6AlXm[82h`^nZ5OlA0XU`>
b[=LgVlf<5Cg9Co8O[GSgDL^FWlfINCS483cZF`PnendUoIS5TmYF9^EjDH248ff
W?DP1^Dae1QHg=inS`59\EHk4\lD7Rbd;3=f1=aD\ALS52I_D;qJA`F7IGL<CoM4
8J7KlNiRG;661N:N\9YdRcaERp`>;4g]8j8\la[F3h:PoPADY\:\?cPTjj8Hkl4B
Q2jI53>g[CmL0jTeDVD_N<2Pko?W?B`DOKB@D>8B><X8^@LDQ1]\VcHHNQkg216W
HRmWgG21?dI9<@LCHR_??IHeQ>ETJ4B8XjKNYmSbmGX@HJEo2mRLBa5UUYBh:>6`
6epJ:oD?of:WKXD2^FN^_`K2HCkC`cE]OT8]G01>UOLjE0m;>oXG8h77>[^XB8j9
B8i6ejfCn727_=onHY=D:6kgeML\`G=@Ci]lm=a[2]OT=1^E63:^d82Pe^0Kof<f
3NHDPTj;NE>BL?ZP:5AD<VJf?C22SMW]dKXk01M[^g]qFli4LB3j8]cajf2WSfQR
??GX3G6^10OW=8BCSa\Onci^?BU`STlThY@M`8d1EBjm`eN`geoI`_T@bD@]Bc=D
6^`XDGSC87RHRaW\<mN]0Q806IHLD22c<nZn]5<[OCYn9HbXiLg3HTPKB^^RBe^K
M?N@XfHW0DUKcCKl<gCnqCAKYR;fnn4S14FHVH9Cl_XiJFnNW8P;T=o>4ZoJg<dV
DHH[dFS0keRnqK`b_Tf[7LgIkmICLIU6ROcCJAQTYWbBbP0P5_g`mE`Og>_LnE\:
W@4haedS<AR^h=VcXX8`eaY@hbe\ooUZWCT>iFQX_\7?6X@eJdLXVcI2_o:IhU?h
S8MiL<9JBZl`_7LY`WelU[6UXMnKioGTFF;m<lPZcZUO5LK]ld9YVqcdNKa8`2=6
f[oQM16PPTNTd`NSG9n06SDammD5e2=F<7Ec[2UJDLY[GoeEUU4bF61PAMe[VeH7
jMR1?lag8KGHmO]Sj1A`MZemdJNibg;3eTOAMMoVOIc=W_J3gF:jP[IARN_4<S^[
nbe=TIaA3K_TF`4S6JBc1LMHa1N5edqZF>LHX7W=Y9ahf;O^Sk[k<i@>hCg71eXV
:J5LSU9=SS]:A5YL5Uo9@WT<AYI[ghbMGRN]@bim?4lCAfm=@A?N[:=ZhMgJ_3l0
>g^bQL2i;cVNMH<^X?lhD54Zfc4mmYd[So3kdg>ZSn0jYDl=gMd<<IfH67D=]7WO
IP`b1ihpAaD?Nf>j:<V;Z<O5\U5c[46GBUmZ@LRQ<1almZ@9EXQ>XZh=\7_0`nDg
3ZQ]C:4RONJIDYiB5aQN9cenYNo985O8RUG8W:UT7D60a?fe0FYPoP<Y\4nUL`jO
c5`5K5Y^oI0lKhDbX6aK>Vc<YjFRM4mBlBKZlnYVGRg8a5M4pn60XIPU2LDZYAY5
TDIEPMLZ8bV[bHE2nH3:>`ZlmS@6q;F;JBOQ=N5_nT5f;g2Pc=a=^R5[`YTmi6Ja
PCV:[LYn[c4TN8N9AIUWY=?CMN[nWh9YM76@<;DZVSbZd4\l^Re``?5fRUlL<V;R
8kOWK@CN`DSgZdC`b@@nn3?n4PhfTHiWGj1=b_H6MkYCB4bXiD7H]DJ`n\ZKV5;o
`kMX[p7_924<[gCeDhRmca\=C\AnH:LCX6DK750X2jeh@2kUVK25MkFYHl7>?QnS
J1L2>Z<?94jTcjXc3EPnR3]79HF]JN3CIce5dMA5e;K=g1K^Z<>[PU`4FY_nCYEL
KP2:\QMRQ1aZ8;Q=MdoHG1]8nUWnJEI:``g:;^IIkdKcESqSS6`_;`o:JLY4S=E5
3IcnREK8BWQDIcJ>g?Qm`cXo2fR_dj<2im@YO<]F0KZ6]:_N1JKT?F>BPMCOCj3<
a>:mEkaIBW9`mLn2LOdMV<^9eQZFJ?`UE12_TTRYDc3;ND68Be@X]Fde73HRd7H<
oN:E9WY6BHCDNJJHn5gM8d6qIF:`k<79OHgA<WmUBT_`lYTPWiaQ5K<GTBbQgERb
JcFl<RGNO>?YMBIXHIeRAcXf\mjoT4YVEb;IG1iWX9VGPiH::ib9ZdCBf^[@O4>8
L^;CkLlOa9F7EBXBO7iBnNOmC3CmAkW<?jQdF8K\X:9GlY5A@G8RPC09i4jXOg79
q7QUd;2TT7Y5?=hV>ehPThNdRSd4A\ZGcOoPQ^_eL1<cEd4YbERQ;8@W\U:qM3BY
?l1JY7V7gIZl_AW27YYY9kbJC_ho91H`=ladcMUjWmKAGT6JgGk[J`7h:B@N[g5g
?6S`SHaFCX8VUcULLZ2>NknfZ52aWhf2EF4_Lk4F59LRNkSQS^9\=l>H[EG5T5ak
06_oIMNMh;W9UAXdKhQ=>_8lCi7oFd:@EBFhpQ_5Q`[\8MfLME>4415a37@WIcAF
Zno6edVH=0O0`DUUe>78jZdmN9]Hi;Y`A27Nm[gQ<08l<>Dmc>^E?E=T5@XYP\A<
5EfSZbSB>l;H6F2GC:>cWWSbi[:OMUFnf1[FM5abhCSLBeJj0U^CfEVLNh@RXP^T
\dRPMfjfllAfRp=i6lm>Nhg@]4M]S_a>H<bEd1E4jd6]3K@A5B4a^94i=[kGDO5;
PQ[e_mBXM?WR`AJAS?oNE>b6BC=KmaJ8J9a4fEl47T>ZcTfhF0C@?AlYhkiYAnlG
gBVX62:hIkbjPZ5m]We4XDadXE4N0_JENEMES9C3N?VALWjHWVC4hnqQ>RK]Q2=C
X[Y@GISSjU>c]KSL8nKIP]U_OD=CM6XE[MbeREfY6IC@S7N\FDY_2KR4NkM5RKaW
XS68gKk`8H0`=AUU8O3_3DZObgFSaf[F6702IZISh0>O5^2CmcQ8\\iN:QU0TWhh
TaYMF_4`f59J]>@IR3bRNDDE7YFSOCWq`kafYJ8<ReR:na6@Z5VmFF4kL6JIAWEA
q>2AH95Fm=@NQilB6Q63k4>cekMmd7gP7L]NfFQEdjP4;3j93_VDK1\_c`9;cH;b
k1FCk>=5m1a`lSX0enGD:D9g1eF0S2cp02gHn^IYATR\P[i\6[C7fDSZ06>3YPE>
nPAaUbMRo9[j]14Hd4XcXB`H;3@:QXMXG3YJ7S\X17ImH8kNSESVQ7TUm6Gkm99X
[M<5gJYEcAdPEHoOb?I8SgN?5TmZEX60CeUU_P`6NGiF4O]^SKHaD03ZXbALFJW?
GADOgNTCpbToL4JO5f6b3MPSYM@@ZL?9_HB<Bn]mP]Ec[OHM2f4VFfXCF\91]I[G
i=Fhn:m8XeUGiddTGh0jG8X=M_[VQTdkNoB<Foi\J?N]Rk?N`<FhP`1Hn7VBhSC4
=Yf[Of_;^b<6<o0hlQk]550f:_R`M4?D]XA74a:0=E73\k55PpC^S5kkaA]NiOKc
WFEB2foEaA<9S?@2n<RoQi5:Y\iM25C<g<ORB?fb:W7=;nYT_BKUfMDE1H2kE^G?
MPUN2E3d?EF9TARB^OSEToX4K<=Dgj2H`\@_F`gBdX=YmbOjDWhMW4`kV9=g2KFe
kNUC4=UEmG6V69J:e;J>dAXLN7p47;2;X[Z:UUNdW0`K_;]cidm7[\KTB\7:jHQ8
K?FJJcX^8H7[hTOC=T\G1Oc<=gfElfD@gdTB8jl8U08g8:\bM_e?[AT76XW2Xh;5
W>Z6_K1_5E6mD;cj^VNSCDKJK?]bf1ja0kNRFYbTkXZgBnEQBX76`AhSHQ]BQm;5
QlPqk\FaeEO^`7\oKE`c>3`H>AdCYo>2ihCki8?U\UK?[71Qih5n9Pb@B3L2CXaF
m@_O:E\Mc0c6aUc7;dNGJ3V]@n^YdoQ]DT@]JMQe`R^4Nm46^=DLo?nRPo4<PaMi
i<K;4U8h82OMM1]\;Qk=J\R]KA3;J[cddNHi_c7A`80TpiA8]QTZ[nhO?RD\Ko0W
^j9aOn]QP5>hMm5jHHHad9bAD8W:0WJ?GlRg4WNT:KhSS8?C?DmHXHB]`[Uk]hmY
[=PnNc]Q8Zl_?b@1jl5lhf_RTD]b6JS=cI[i6@4>^_9[JA=l\g2_7IKcn^H<Dh<E
`O;Y^5Q13CdYbZd[WlgCSp\WccY[hN50GN3FAAOd9RD;;]5[e6B:LnJAUJnl7GIF
<B3kdZ8Xhnod7OomkkMb9K8AC59K[HmlN1;eAY_A[CP9U6j[IKe5c7gn[NW6]SFd
d@[>[4?2V_fV0=SV1X@njC5@[Xd_R\`KWeoc6;_^>;W;ngY<ISYcD3YeXNWE2Wqf
[TCY`\IQTf`0?OHFLHaBeO7XTUGfYmh2LPJ9<k]nUDWJb>V:lUHmN5RGbjRc9;o2
d1m<CRJl?c<X4ac4AOV2DAWUTGD5j8Kfd69gjPRPR]m9H5IlAVPJ=Vchd\8;>F2k
naR^U[F1H_>>hbm4Ea:Pek8X<^^kVQECE_DgiLnpKbYWg@BQb12@:0PNG33L[DO7
6HC5\SYP9cL]?NPID<<fPjWXYKHYR^F3ZiCGeO80XM9p4hiHO<Fl?U]O;R;b3YZ=
CHKAJ;a[bYQJ=mXaD_6`]MeVV?:SBnPSb:XU8SdOh@J_kd:9`BjjM\][57U=XY2U
VQClN;A0[24L@?OSZcVoEG3]6b_H\8MR<4Ea\ei8ROmlFD]:R\FUYC[H9G>mXc@:
MH`GIm5OfimR4M\OZ[ZRq\o?W1^gf7Nk4?VDF6H04eWEUGPoUaHGmhlO@ao4h0fV
fSdX:n5O5n7;]Goo@1^6B@ReoNH^^Da\PdI28X<eACR28;PQRM7l1?aWoWBV^c_Y
E>n?VWk:>0YQkIg8AKIA>GK;8Ul?D_B7bn][ZX?=0LXB``C4AI2hL<4]FWTg^q=5
On<10JbOM?Fjlg@e::]0?aCO7GlAd`T0?<a^F?VGBO[lPAUFRWaVg1]mf:V<l19@
SB]SYRHIidm_h80;@@]\LX^O5_A^Ufd7gH_U_[X;;ad:86McHVg@ENjV76hA:WH8
P?6NZjc3Ld_<7U0DJk[0RH6=mk:FY=O`<O_0F;q`9eLCl8GR8SBcA]PQkSMJWHT\
jFQ9f<dFAdhRX6GD3?e6Z4g1_d;h>QO:>Mdo[;0a\jnPLUdgAV=lY?;hEffFDZ6N
jF^ieF>YmS9cn2l2PojjNdn9JJA^Q=[Id]9;nCfL:F2A^59EeDF<8Wch<=IcgX?m
;<Hg<^=HJl1cTkiq59aC5dIXHXK_\9`^?M7DDaYNM9YKB@<SH:ZLDG1jk5oB^2U_
KV4jVB`[PfBTC>gdE`C6iOnU88fO>F_D6FUQFd3Xf9nb4G=hAA<^APY^l<lV?lA9
9da^DgXaYRh?e9Le5NCG8U77J2lconWF6VaZ5ak?G`k3IF<Ud1NKA8liplZIV_NC
U0Nnan>^6HW_ae<S:46lWXcS;5Knka3NEeLD=MY208O4R9eJG2a_mIkCmG:C=VjC
aL;O>lAYRPk6P>dXCa6_@l1Sb<B]aoaVN6<37T;DI]R;UIEdBeBS5RbK`@]b3=@d
2X3YnmFWRP:;l?^NGdU35ek5oAY]1o_f;piJbJL\Ci2SQiNeC1fFB[eekG12OhK0
QO5IZeGQAq[dcOIa4W^H:]7:H1[14K6_l:1C\mG2l4VbJNa1E:OMc_jkFlc`OfKk
F3]Y\1WEfTG>P1QgU1TIgI3]<1eIk6S=E3@CcWfmUABDUGEkRclJP^m41abB>MAK
87gX9S4SfHnSobGj2an:iEXQ]meg1:34KdXFf=2CBSTOUCEIIEpjSHbA=EM\V:BD
0AeeZGRKLDTPSW]]]G?edb18:]\mc3\dUT^cGYQPc_:lIh3X^mH`eZ[U[C7Y1mW@
SPfe<cAFDA5iSAfneNNJ\]LH?ja;4mmS\_3Ra0i:Ue;hHfGC]VX]94>fCn_lCmEN
>h6e5AFZLT4WEO9oeO0OhnWHE>Hp=Pni4_@dLbT[BS62_mQBU_8:]E>j3^4h8XXO
K>V7:N@o9=@U_J9eWHS>H4WU3ahI0b:JE@g]_g6Hdb<]U\?VmE=?Zk4DEApFI;mJ
;QQ]?Pan;2RF>mAU4=CK7dR^R6K[6\?WeSk7KeMVF2I`;GL1g2G0QfNnJ73F?Z>_
6@KU4RaR?6nS[^;\hGO6B;PJc6K0k\WNG8XAFhU4XT?U5cZiJdY^nQLB;lYZGAU<
iDAU9G[kk?>R`clR0976WDPneJQhi4MRM\QTCgiQ=MVq@c4GOYlcS;Z[J1^F=^dR
YQJhi]HqcV:9V7b_SjQU>TGP5_E`<Rl:Fhcon[0oX[:1Sog@KUW@LE5aMUMTf7S^
WCS`M7Tnc0McJUm0T0jbMFa^_@E]P94I5>0ZA70g@H88`50STSPVA>`@M34UUOGa
`UFJ2@ag6@nkgi8jTJ@fW6?Ka1:@[aZ85F10Da_73:2LVb=eAL`3f2V@p_22[cj@
j1;f=FS08]g=mcaH]3O_[ji\?KOVcT@b14W2@gEWLBGCZ`dD1WOT2jleS_`>[LIn
8mH>RmSW\[C=dB[g[7UEY9R\Oo4GOV0<ZAE11>AVJ4>_ib93X\^V=IoReDOJ3E2R
YmD[U=Lh=nAW2TUdj7^IdThn6FXGR28cZ7^RYF6aWqSe\VF5KLjfe<3>6>9:;15R
HLd[nKfLQ4G\:3X0[i0E]7MQK]@[ULMSACKHlL4dcmSVNmTZ5235A<:5N[P4F`nV
ac@4]4Y\Q2oDg[lW2e1<dO<EP=M2S`GHN5E391jOS0[gj3o:lo366WCU\[D:98]a
6o@be^0b^=\k;Z_B\2a4\1eCC`qA95HFBJ^@fdUIR1cW;HoYnS_a5^3gMSBHIW;\
>jK5Lac95f=]T2Bba;R7IFXZ>8]ACVmI@Y6QDco<ACk1V>ALM^Vicn2iISf;0TNj
JlAbm<GigRZQ6fR`MQE7R_@<`G=X^Go4k0CQiDQCBc0G:]LgVRFiHK=<jD?SE=\B
?EBZ0=N75IiqlHoL`K_n7J`_>1>TY66jGa\7`N<`9H@8@I`E1@bcKQO5lgMcGocU
IH`h0Q>7daYMlWKkWXaHaZOGIBDXH?BX5jZ4ZWZOYg@Jf`^UA3R\8nVYGPRI5Y_S
ghX6UF[BUmg759m8?jg3aFf1QTiKk\S4H^KOZeOXHC:8_GKKI:DR7Y>>F4ESpdUJ
ghfmlXL<=0[g2=^LW[Q:<V`V=j9f?_K^2E57XHelJ8`PRX4Oj2WCI:MTEhN2nd?i
a;;H]3`:W0AX??iB^i?J^i8[i?mf3n38gKUUWj6kIC4O_P?YQ5c>E;5>ULH\7Ehh
mS\L=3:FLK>P@Z5^4GYghibMLW\RG3COA3m6EVL7no6oap?1NG<LL2WJJH6^=iJ<
=TeTG1iZA_K`XRV3\9q9ASW7]m7J7G:b5[kFlkTQb6i4Fem[1Wa[Q^4Z9jk9VefZ
HcUZnnE5;@lDSWnP10;9b5`9n[^Q1m^7fVMoRkM7hU>fE;kTNW:WDiXjL4c1<\7g
bZ]POGKNXC2b\iYGn4657eX`l5ZQ_ODk9Z_1THDj1f3fM0nF4iWh25@?m=VeABmN
A:[q>VJ2E:\ZQ2n8nC1Rj0X8PQ8:;POhH?ST8RXE64n?m:8NbP3oO=mo:l=W>Qmi
F1gN>AC<CN?LoQE^MKDKo6XfJ1iB`\L`m1SSC@<Z@kX2FG<9K^nfWH?5WjMHV\_M
@c9@i95YFH`RoI9eU_D_n@@DY^@9`7N:`f_Y>hm6fA=jjdkT\JF4pbl6S4?Djck^
`W=a_35P<YM6IO<<dWCFnmQ6>^el\2PDa]_XN\QTfW\e<YhNLfEhVbS=YUn;H`6j
RYMPndZPcoBTfbm_?`VFL7f:QE^^V5`Bko\n[46Ub;YRSV0SX1hbPYB[_l[jV`R>
:kV>3gBV5FgiAbI0Di8;a\j4<CQAD[Pi<GS6Dq8@`d6a=<M=UcZCcVTF5^QG>EBo
;h;:5CE3;8<IFeX;i:Ti^MBAgJNm>I2_UJa5_k85jFA1kGlX[8\[lGXN52X\Vo\c
:6db5DBKe5\IBY1X6DYbePOO_agK:?aNU>eK3A=_1g6oAcl85Z7N4gS?ICMi^>\6
6aKiZ1JMY@?j8YOjKm_]TLpZJ9GPF>mMd_RI88CIPG[2_1:eU<no3W382P[_0@=B
83cDUVU<J0\D2C@0G7[OJTWZA]HBm2OYZIL0m3\EQGOi8Y\hl@@k6We1YdJ3Ud[;
9T8ggb@1a03jRUCk7VZF@[U\b=Jm:W_Yd0Hg^BJ=dFIU_M7hi14kJ;7_QK]N]l0k
DIU6`LDpVOFaRK3[Z@@19Um\8IFcV>dcU^EDYZInm4cKYa@VjKf`8Io^L@^8N8ki
Th1P_?5PV^WeWXcE_SdIQWJH@<F42TkPk0@Q`LIJL2[gDFi1l=Q<VPQR4FQSdG8e
c73>R>Q\HPD=4\2S_TJ4I9o5eo>egl`=kB;XLd0efFnYannaIl6ddcf8pY1WFlY0
S]_;22X2CFHaS]^<ccI8a5EgQm:@5`WEDM[fWbH`?UBc9?PkDY_;j53icYRa9d24
k?de@334iK_a_0oH8:W8Nk8gbC:^[T66_R^PWlg[]b`5F7cka_Ke?FjGOHokQ0Pa
a?7[o?dd77Ya^I7CZ:bTDHG\3oJ><H5cc2ESI>MDdqR3893`OE^e\YXKKC\W@8da
JG5L:3X=XP9D?\N4XJmh78cX\hdL@LOe5X`<Emce2ORX^ST6>`\@lggh]kk<@UTf
:c0R`HVZXbfgj[[kNcdVAB\L8J1XOJTWP]eF7fE=V]j;YZ;P0k\gggMVSbaDUge5
840Z7HCTj[02if9nQJXDBgH?fHp]WHOSY<M[L2EEiK2:nR;B;jWXM9>A`>`3j9RO
\EU0;lNeXZnHOFWYoQ3V>j_[JKpE:M\mYk\<a5[YKbc4Bj[GmS`CnmkAgPSNO:K:
HoV:<>oa?F`fLd]nQ2]fcH<V5AlE]f@dlfRX6H[?Q3=R9jJY6Jd\bod3@P\A39PN
;LKmXW4oo<2O[CCQ?Nd_?46e\bXlKQn\eSeXlP=`\]fCBaB]n=M\ZdI4E;bmcl`[
8e6_lKHA69fpEFDF5N2m>aGM`<?\``kVmOB]DMVK?V12POmJBf?idXmT0XK8_83X
nEdg]GnUg44_Ejc8915R4GOl7fQW:I\lb6RDXHVS?k1[VUBO_^V_Q5[<Lh\9RXDK
T<Dfl<4=eFiVnFTB;[?l4O<P=o5jJ;?WIg0`XLYdDMA9;IOR]_KO<kUkcViQqGWV
N1@helDeQoTc>N=eYn2e=Y69DI343DlAG@3i;k14akR:E=TQTR11P@2`oA`BnGJ\
J3lX8B8=NJSfOUS6djWe_Jm1NOF4[5V:OC6bTeB1\9LmD:j3WD`IFgOCOfY7aU>S
FMc=JBT@>T4I;cchhHSA_J1l[59?o3h`f:PLJgHF53^GOp1<_R:Bm\g]oR?9nC`F
j<hYn;7YW^:[j`j@fdke?hE4d9M\X4H3Fk[BiOOJ5bJRN11<<iS003f\7P^o\Y?O
jNI]OHD597mFjniP1WLgN5D;NYLZ=kP[b>?R?oTd:D1mT\7XAb5RU6fIfPd]jIh3
S\eWEZDAGfJH52Sj9ld0k>l2@LU<Y=qbM5na9d`bYC\kZEmLInG]jc?k\^k0J2eo
S5_bfHTfeWN90=fSQbVLIUccanDXo55bIS=AD3hFnhjISmUYPF]0KN2G:`1k02D;
4W9lFnKDYTi9N4Un[=XILbBkPdic9Y`MkMWW?<<F99Hm_Z>c\8`bIJ8GA18`B3DT
VK?j23;UgL3^=NOqQ1Vb4c;QZ<76DndeOAQOi<LE;KHkX8@g;0dZ;`_SX;iam>4U
?35[aI9n[T3H_mb^QZPmflRS7oAN?U><gPo=QY2hTXl]Yb@V:YPXl9QNRVXRcSAb
`NZleLg@@\TfFSNecW1SV[]N7NQ7n\CG0b94Pa=hTFm:]TMMYKDd[Il^`RdH^QCk
pL<gY7>_I[n<GMOO@j34nl`ioW54P[;PA]H93`2Pa5Q@\i[>GKBXmBaXjTM>`PQ\
5LH389RflPB;@5PTlN]4N=8?a\WcZViP>L=@NHJ4VDN22D:PRZ3]`lC:^o1QOcQ7
^=6EJl9VCP^13o1mE5oJ]0b9U\@CA5R<:6f:3hA?l;Qj<<^ERpXJ:66_>4;3:=l;
hjK3P;M<[n8_O<VD2;dlL5B;nY=E2MkRaIV0<QRZMi5f[G0OC@XK1KILAFk?nlED
bI6cPJkF@`XPQK3^2<f5n[nQGc>lEN_1eA>0N?D@S;imV8S>03C_lMOXZCk_3d^c
ldN0`N26D?X7X:QT?o9[SX1[8_kIT7LoW0q8Uf5f:Fl^R3gbfcUeS4>fn?[mP`53
k1c:JWbS2H@P?:JIHWE1^f[RVQ>9m=j9:Y^8d`qWNH7;4XG;\Y1L8K\0G`P\Bf<[
?_j1D3BdF<l7`kFbOHij2JLMaUjE<gKQ^Ebdk@lWCXnH2T`>4:fUkbGFGn3APBea
h>W?23b6i0[FODGV?`RcKkcEmbAoA5;0N`[OAC;egHoQY3K>m4I1W1JGeAZ>oD1a
[WJ0cfZSIk@fEYl<[IV>^f`qR=^oc2;1X\nLg01om0G4XmeS4<H1kf?ITQKLGoJd
W1TVe<LVTj5keV?O2b3^M>:VRdTfab0fnElI^1hm?P?65[cmCob6;I?L[mZihGX?
m;;Ic61<k\\HG8keFhZ7XT]45cfdJM4WnQ4\;lVDGA1hb1IPC:Zm;1On]KQhU<n[
cDP47g6;pTRZQC3CDTJ0jd;Dloo:36eMn8A2h\fONIIIH4RPoUS]>kooYMokefcd
5;H::<HB=TiCS=b3KH7VfnQSjaR:`\OkoFGA[MaOZOL4Wn99<=\;BH=[LTmRUTJ]
>RZ;;Q;I6BcIL[N]^HKhGhKP^\fh2UYlWFg70E9kSLF6<[6f_nbWn]0a6pAhZoZ2
m:4jX@VcjU9Sl8]Go`?:6[Ne\k3C4XNY_X`7KfAjIP[h63B3fSHbKVF;?9AdMY`B
Bc5m;D3LUi3Zl8A<Ri>T<hNX\;]m=71QRQ4hRP6RIJLF?_E?oQdFa:ERD?e2H^9M
`K5iY3Q7Qi0mEOBOfj>NB9bg0PV78?j9WFe=LW8b>mpI<\81_S?]48lLdSDo:HfL
5=LASclLM3nPDO95:C8QWm3eWTJ:0JebRjgVYfEb2TPI49bgKXTF2RUQHVZCVHJB
51ihdlhM63a6]Z5J8MjBE6817R7f@<D^Bm8n]I5Ognm0IclVCZ[F[3OMFbH4biHa
?iCh_]mUb^Icj`W9<W@H7H^o2aCp@c]Nh46ZIIiTF<:h2A_bUbiBCISkW5ZF<[cH
Jjm[R4C8@=1N`an;CA?>ba@\k]aA@1NME>H2MT2S:7oljTDL<09PU?C1X<ZSZm2N
T9KEaN_=5;of_gJiZ\83kJLCbEN5Bn:^]=0VMWJSNCakN\YX1CH0UB_:o`6Gbf`Y
HlBk=D=^VnPFqQT8MlkmdJlTXIi?k3gXH17b4TZL:SWLL:b2J``:@oSGmVeV1PlL
F7LHe57@g?f73Q_mAfI78V5N>1G3fbKX2R8_Q5Md<6_L8C8Ul5RnEjmLK7HX22<c
JWA_KcN]PERU[`Bd_JUPfVniQb5T`e^=S^_[R5M_]dhDfS0Q4PN?Pb?b5boB8pa=
>JE3GQD3M3Z8;nkFjFdL[ID]eWEUl\``SPSPJfj8lcpdQcD<HCWLmm2o7FTmkY6f
i8;d6Gi;5E1L]ABXoZ[Lb=6i@f\T2CFlHD24IoFado;dHaEg@X?U0;:UBMS`EY91
\=caG8UQeEl:T42Q044Kh:05GW8@Gce93AM;E@7mYTF>:OS6\`0UYcFoP9dGnB8>
`l6aSea17n>6e;d0d]0WfGI_gRhpcRc6mVEl2aBCDBnHI6lRM^\TFUiDlYHNK4bT
oYAYi6O17ZTCkR[4eh2`ga1if0\ccjfCWW]X@MSRCVZ71CloN[XC8:bUZ;Hb``AO
7Ch^mTF:eLP6fG^^H?BT@:3;9ReHjcLo<9F\@HHCH9H^7COicSAR8Aglk7I9im^E
LL[FlTDBnJ]Yp_<MakbiUYMHCeZaKeEHaX``cF0l>lIk>2FJ`f@0\:_P[8fE1i1:
UUTYk7dMZN?V8_SjJ3FJ@TNj7^DKMBo?6IXqHb`^35Jn5\8SP8G4CCFBoCV:h7UP
]VY^3>DOLDlR8^5=J9cB0b[]BiN_=@\:fWH6>h7kecc31M8XIlJLF1U`E8fD@CDD
2kSHYWDO`Jf<Ka@S>2RXPG:]3VN_l>UcCM4e===BW5R2pENBd25Q<kHA0l=C4lX3
kcC<fi?9T:b_^>jiEP1m=>B3TOAN6`HC:RKd]`b@Mm1]Ueo7aHK1K?[nO4EWo45U
ki0h4ea_:T]kc^kiMTR[2RRP0O5?:[Jj]=0d]<eiGPUQd]aoTl_Plp7O48boU]9B
bF`>T:mL>CWV_Dl7kXAbnL>4FkNni?BZ^P5hafi]ne2GOZk;`2_Xc3[g\A=?S\ER
ZKoC:CG@<OVH`_3l5K`M=57BFf:WZakHH516UgdAd8DH@4acW3QWP?D4LnmgZApe
o_VM:DmZXaAflA5O`0Q570jLhc^^1;;DX2\b@iU;=e3M;>c;^8<4R`NC_^ne>bgg
=E;4UiWh^HVMj[b3LE`91H[Kmd9PFQkK^2^?H5oeo;@AV3JhfZK:4`Z0I4n9Y=;;
V>n1kRLqd5dcjXo9hK2K0Ya\_GNNYd;ePe4kPhTF2RDW4m6C8_B::D7RO6oYJX99
Qg1O=W6eb;=WUGo32bL>Gl`DJVWPM=M\MGUFLTS[KaD0B>X[ilF0eGcXZ[9<3S;c
HGNO5H6PTiY2e<<DpG[;SITiZ?5eGI6gBQR6?=e^QJOmkD3DKUDHN1QW1=`RT;BF
lBA;o]>71d_5g7eL7UmZJim6ZFOYX9CYGNh9V9B@oH5SUST05LiHFAT1L`]UGm7Q
Eo9ZWj^71>l2HDajLdL:nD`6hqo_N1dP_f>1JA6XA895Yg>6p>^_=C1]YLf^a<FH
DDVN=mTV8=UomhlYT5Z0n34b\3BjoBbM`NQ?Z`eFn60YE:4WEZ]BO:7FVi>1kAON
U5X88kQJUSQI2U_Wl?n02\6<H>M>jUW47mY231Q>dLem7dE>Z4OZIl[OKpb>CI`]
42nT7\`h6El@hfI8>Q0nBbW:cWg_9f\6CK=>EdNRQ?Zhn7fKeeZXJig;6\<UR<mW
^G`>Rlc6[7lZX_Q[enA_7BcKZNYA9Qgk\T;YQCG09ZVQDM0Ul3d3YOQaaMd61jaS
^XqgOIf^UZWaaUQ2?C4YJTkRdLaRHP9jS4Z]MMO:_nYBDIW5TLPGTMlahWTXL<j6
mWTa9WheD2Vj=E?`]=c1C79BeQRhO;mpLHFIBZTF1Io\aMY?5aCf?ST5>NmoE<Yf
4X@8HK4YcH_9NWFE4<<gl>ahOE@8VFmQ_Hi1RDB8PUhcnndEK]`oh[e^LoL7i_3V
[i@XQ1cgo96l6L;ZZ`SQ77ac>_S;5i9I<g@94JfKq]YWCBccLeJC<bJNLQ9eZo0U
8nHFMQ@;];4\oiV;fQAnf`P9_^0A@@?oVCRfn\JKT\@jL3:3mV60?1`>IKZ5M;NP
2YP\?Xo@W>G\X0n];coN6]<IlP;A]jmen9A_@m\HmHdS8J=bOqf@X5^Wb=1:aDZQ
Uc@gHg\23L<kPFUnDj7=o@fUP6@4a7;ak0gJK@DPA:gPNVWEZ74XTWC;F[E;9XLM
;0RJD@2oT1EjSf0Y8__JoM\31CTJffWVCWCIPF1bAb^Bo9ZV4HFUhgS3M?q>]dVo
g:1?cnlS2ll?NTn]CDf\6GUlIFfYXRn2C^V@F6>AiWk9nJS@h;XkD8?Bgb6UNoZm
;PIf>I594aWghG<dQnWg]\Gh0bo>7RmoS]bWK>J:m]GMk5;]1SlB]E@0Q>m:AhT_
23EqKL11EV0Z7c@llCVScY]@FVB2][KmT_kj`E3BQT;UhP@B`^WJb5lCBa==k]J?
?X@IFodAdPm;^55L9mP<=]RR4TkKIAT1_eUl1Y38WQI7C3]h58[T4PT_1^fI_O1i
Sd7?V8N6m<XhpA7<nGQi3b9i;cbh<XCCiEc1[4[jeDGAMM<Zo>_]fFgkMebi0[;>
?miqn@<_UK`E3]RR5Y>W^nf8<aE:iHT9c:nU2\Kj\`mZkZE50P13mkVOeMSOof^O
A2fQ\E]PH5@Ta[J\ZTT4:d[j2?QM9o>RL:kiI=K]iWGg?HRR:<01F9KEF:S9K2X=
\Xcd=ITF7<U<qD1MU8[YROdNK_`<Nk:N:ARdf]=IlUGQ?5NXI6;3<FffE0jcljfD
G^P>FY\<9\>m5DI3dQh^9[L37Rgd7Ec3jgf67h857i;Iol?XnIB@CF5f7ah?:oj4
f9=>InFPc`?aQ[g9RGDn8p304X3nABMeeK[^ZBQ3=M=g>Akaj2]10M?SFVBTA9D^
DLELJYA30fXien>P7H2:`Z:8?NLZnZ_J0ZIW5\YPfQXVJCD12o6;gc\ZF>IH6_=B
naWBG>kOXE@?b^EIE\;fKbfTC2\ETnp?>QV?ggH2_l<gKQRl[;E?Xen0XDO1dLE@
JmeK`9@@]EP8VC=SH2CQ_InX[el8a?E1Tk>ojLba`]eMP61SIP6<HFf^6IbpA2aC
OGZc=5ME;YQl88334C@FA05h005n2IHCRK5K@c8i3oh]_VQ?Q1^b>12AXek\UcO>
:_N6FTTQAY_eX5^4442gee`ZW2Rf[VHdNXi`@6BYLfT^W@1GKT^:V;_;9GP=g\fo
g6ERq`]^4UPn96YXU4YnbMc;E1@Iab6;RQ[Y?QVKKRgdYW3kU=i>:_M@KCiZCh:e
hASYMPRMjjBYOYA:Dbb_fIZi?>UgBZjO7fAmi>RK?`cbfUi>@L=@=?XNj<aPDT89
1CSV90P3VQBk2p;g^<WjKaP58MOiV:B@[85YD0jP80E9m=NF=PUbRFn7MTCOZ`U[
`Lc]00K;RMbHMfMVdBY6eS;Te8P;R75U8=?I7Rg@=3coekFe=jG2i<nWWNkEdPBZ
IV>U0S\J6cWI:I;iW97GQcqY9CH=MQ6ASQ4TUcGHC`hUNC^RQmQ;iAIQ]bO\X>J\
cKb;[3>;nU2EO@dBV:Hmn914EE78i<?^9hQgbOebgDeVC5?JQ7PCTJ3hab1B;F:\
[6[?;ZRSjSoYY2nZ[k@fO@V`c>M@b@fqXA?07>:J_C6oHBW4h?mE3VZ:\YED:`RI
\>DnbCK?>GAcl`1b0KWniJ9ichOUi3Dlaj]Q8;c5d_7TZ2Cagh1kM<\SnL9Yc\eD
<FDhKRPG>In1hV=F94UaQ>HD:[anIY13P<`ULV;Pp1OgU_i7CZJSHZQE>9kXbl<8
VeYW;ddkg^TaC;S3qnD<nlR;=BEXmFYWC7Z1c>CQ0Yi?E?WBR;9ZlSOh5S=`B^k^
INJGaUefMSbWn`F:6V5EFLMIof8TV::EalP<Pac\GT8S2@QNDJIZg4kVT@nicbCa
STU>1TnfVjEGP]Y_@dmWjVD_YqUjd0j>eCHh<i17EH^a7eY0PEoX=@[<k=@bI4>m
aUR0a8E8MII\eZUTK`Ae?DUfTHGaS]6:gZ:6hE_PH4Qj]5Yacd]ZBY5^?CCRIn1E
a>6S[j:5fW0DU5__KlJ8S1XH6[c<dB=DL8qHCg=H@QSSJXabXI[QgiH34Xd`0DT;
3a`e`LoVD0OV07e\8jAe3b2M2im4^n_GTb0dT`jfU38hX;0=16Q5DT?@l_bPcECl
HlWEaLDY\lVBI=R=[VHC<gAOAC7H=]EgaAD\K]\^GjJqULkC[5nID:iAE?AFU_do
T9g[hIH^LRnWf2c@WIaMekjeB1GgQZCS_BC60JW1n104J0Qi7k1Q`Jo9f;9S@bS^
k;DB0LP:qZ0>RnJpdOX^U5R$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MXL2H(OB, S, A, B);
   reg flag; // Notifier flag
   input A, B, S;
   output OB;

//Function Block
`protected
NcLTFSQV5DT^<YmDL^OdY;C9pAgJSD]>cLCjQ5MdR97E1=@h\NFgik[;m=0>OmG6
1q]GZA28G6<]EO\LDUH@ZbJ]`5NWJ2<5REnI9n2o0qHh09jRpE=<b`n\3X_PnOeA
QVUeWRG=1B3lEE^CRV`IJn1ELWmo\j@pcc<Pd6ALYP:_g=1X7^SD_1o=d1pmcZK[
GGp\GLo^Xqmf7<:XEO6<F^3S@\ne;1jgVlKi8D9o`kLO2h2KUD=_L?UL@DRgIP^H
]HVo^[4AX;m>Ri7oQkbQfJWfEGh[PMFejP8CGMYRhgXY2_p2Z:1R@jbA5M^EVgBB
?6Pd6CdkkTWSMkiDoRco1@OYOlR@^EV3be:98c\U^ee8Z@S2j==Z3DCDl@eMakLh
4R<VdH6O0;85EIa]cINqke3`bO=cKC<84XgW[UBRa0_3aA2G=O\mmGUcpbdA_DTN
AE5Va@f:Q7Z5@O15Bn5[;hU>EnVBLG4;i8`m20GFU^`Rknl\f48oAhkkkb[W_N8X
h9;^LVBdB`oeNLIq8ac]nB2]TTVKmWHN3h<K=T^e]Ti_DV=an8<UYY]Q89h5c0NJ
LWMDmjJ_EDX\aeMO84IKd`G6HmcW8FGOVWKMVDQGg2XX=9=ionEXdU9G[kbVei3;
DD1p5`G6;Z;hJR@a\P<6ETYdjT9A<Pj`ZFlh`o[ACOnV_:@F3BMdR5iJlRj1a95N
>DBk555_[WVW\Gka;T=aXeYGOI6TON2=9iliGnMie``hH^7k=E32IBmpPI2j<mSU
Be2g`hEgJ`JdMYWbkL9LA2M0H>:NO^`XAAmVq7TLKOUhCESBfVj6Lbla>61ZnPY;
W4jH4hjFnG8]Ye9g>P[LnR[1NZ`k:SWB]OD1b7M=aQ<L3H6Xf1`k59bMN_`qSZC7
i6Id2QM\mm\SLVK6kID85C9EQ3ZcIj74FUAHDhfH8jMMgQbTWJ14``CM0^?1Shlc
?TFWJnbSl5iffG[3ENe^XS7JJGNPUZL:q<LN:\lQCj=mF]C0jgbhk^B08YOcTVPf
Q67ea5Tc<;5?S<gb5\i=AJeXVI1oYV0]P<8eO6QPVZhQ_A@;EQGOKhmLJFJI1mWb
kCKk\p9GkXeZ=C:GVM:<dJiXF4dT4R<KF]:MKJW3P10D`AdE4gIl]g_kLieIL9_4
]JLii;9LOY6KX;KC^W=fjUj=6O4Vp6bBMBSp]8ZFCD5$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MXL2HF(OB, S, A, B);
   reg flag; // Notifier flag
   input A, B, S;
   output OB;

//Function Block
`protected
e8DZaSQ:5DT^<LC`5JXd_i6>77eb8VjL3FhAKPq;BC9akF4jV]a>XVWOSO2SE\3T
H8?aU>RT`fC7_k1_3hbAD@T8igqB;RfCbmQLEDNc;LO<bOpS9NGkRpBlHTc1]bAT
a_oJk=1f_XBVj:<]QXG`;Sgl45K\]jNP9UIBq2jmQ;gTcI7SHWa=NS5\RX3KbY?p
HnYJe7mRRn`TPamea?fk`;TXF6[T?eRgMIZ;XTG2FI6b17qPHUTl27q<OVR:?q0J
?@DBo7S^KV4DES[lHa4oXChb<[H6W;l3P7@kJJLQYJIGG55U<JcDY?8h[^7UO^0n
^aI6]0l2;>AO;]gD>H\?;\<b^52Y]Ueo=Eq>Vi:`a;blV>fHABOd3gOm@3C1g3]e
M4Ib^>Sjd]QiDXb0b;YV[=J2O7UR3?DP8mI>LnAGf]BXoK^a2e>TDGT2WRij;Q:b
A:Ll12:pGlK]l40`A\28dJ0]_O2kTj@25MKbpeS;Xa^VMWWm4\9XFOEK@d[PE]=M
2iEhQ:b@McO\hMili6I2;SfE31oPKVIBla8W[e9iWTeVG1JA<l?F<D1AR_lqV5`g
<f6PT=Cc_6lcLJoQd`2dCU1JBHRF96oUZ`4`W^CY<=FVL<V\93fi`b^hg\e?V2W\
65CAFf8ZXhAmUc5\_bAR1`U4gAR;jY9OULWbFnRR20Nd5KAq1<h>o<00A`8`AhiV
XVNUDAhDbNU34ZcN7FF\f7M8fBU5AHL@KC82@PO6S\Iiaoam1f0]gF`K8INCVo5c
J;NiBK?bK^JZbdcE;^X\CMnfg7i8?2:1iW8qZk?=j@D:8b<oAmHMeT5bg7fc^lS`
OgVCm@1LCKj9eDZ2BU\`X6^daXd^BeI0HE=kZTA;aCDhYA<JYiLeOnH]IYp_E0>n
7WIYXVZ1e6`O9M=eBnaPOONngUg69nm@Hegf\O[QL87LD[FR4GF42[HXZcU_a6I1
`b1=C3GLFa0HGROl`e2A^=3YPXZOnk2p1Qge2[^5=BWh3BAOHmMi:D6m2V3R^Y3`
M:?BK;<[3ZBcH9G9KS7E6K0NPS0KFA:I1L26fUPFUona?nY5XN82TmR;Xj1UWDiS
SW2FqDBDW1oS0g:MA?lTj>RFOoWGZNjYiEdm05Y9J8=:Q^C>fZn=Tkbkl4Yo8jH2
1GK]7DHEn32T>W<@Y4YN42PL94lpnQB:k;pZEBTGm=CaV>n4LGgcJqF]RL@7G$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MXL2HP(OB, S, A, B);
   reg flag; // Notifier flag
   input A, B, S;
   output OB;

//Function Block
`protected
;QnaPSQH5DT^<;VM^?jn7@\A2AH3oLP>3K8?iF>gKmBY>YV;=\Mp[1Maj]612B41
Zn<6N1EH8ceZ8PZelRGDe0EpO^6Xal<kICR6M82eU^@Y43hp1TSLP2pLC\ei2mQG
EoO362;T\LEh8LS]PVTNd1SSDUN0N8f0bOIB0p8IiVCSD<KFK6Z<iXoILH<D@YG?
p_eO;]]YqNMHY?OqET6h_QDblB1mLR1_B;E:WOjVYJ\Z<;oHU2aKo^I[^bcdgEjA
>i6a_`da6if37kgAEG;6G2=fI8H]RO468FP1eiYi3VDYmW;gZ[?NpA0eNL=Vk9d2
GnO2PXE0S=Vj3n@l1<6JFiUH`]cI[>kj3=m8>Fe9[LG]\cZ[cSd@cA\8XOCDoL7N
4W09@Q>SH[eQN83V^>BDd_AQKqEgam30\S\;QR62gQ_c?5ZhZBKMVnbH9LPQ6\P4
33Xcm5lRRHfUP@JhZVd\UQ5O6OET4bbYcnJahP^<N>]K3i<^pfeLB:i3@=BC]C8]
`Kh7UchngM2dH=]cc>iVXELhGRNM0N\<<FmG9NX4>FO25o@?4f4I@l<9cR=Kb0FO
NnofU9FV;@8Qk5RcRGOEnLQjYCD0GL6;jIClp9_eIKTBg_S4Nd[80KZ82`<1YGD:
9VT81>nS1SG:EGSj]ond_J^^X75ch>G:hSJo8SdCihB\Cqcj:IBIonaLlgMS;h9S
Ilb]E:M1KcF043>9l=<PnD3:1dgRlj:jNWa=gM]PHn4AMFcQTPcnoWiRNSkUaYDA
I1BXWbP?EnOC4EK]ZaDf2NkZeU3_9o[R@qE`4FHVoOML\7nCEZ>CQJLH;;Rn`lBb
GC:jH>j\G3RUVS4c^Je;I4LN14]J=e<OGaEQW[Xk[LoO[o;WW@^[@i>lp7[[8D]h
`mDjF9i3ADFi>f1j4aG9jgJI;RCS0cHceoUkXOek^>UkCcgQVnkVC4Df^7E;76c^
U1L:LX\YOgLbU_:UPm]P`[>]flGPCqFBfPC=lR69GYM?8GR_EUAjFQMai@Ag9U[<
Ac;b09d4ZiY>mUVPUo=7jhTEWk<OqCgYZIeAVXF]4V32mQSFVbLoWQW>dfD^m>Ee
Qe@FfM:loeBAKc8Efd3<o\ER7dDS2C@9CchTG\I_\4:T3<G^gJkPKlASeVUn[I1k
OpL`JNeeeB[S3WICK9U6Y0OU?dVNPifS7hK7R=kU`jTFgCVk3M]T\bIi:WZ;c]3:
d\LbXPH[g:?mIlVAhJ>TDQ@Ipj^[mJ2qQ>Tn1A<$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MXL2HS(OB, S, A, B);
   reg flag; // Notifier flag
   input A, B, S;
   output OB;

//Function Block
`protected
;_L3`SQd5DT^<b5Re=5m?1^;jk@;OoAIbAoh0[8M`FSQRhU2QF5ML9nSRbMB7MFD
qFnNSkK5ORkMNU4aUFEfceMkb0M2MK>gE^PmbL9OAVg[?omOg@RD6q220iZkRbIA
`Y\4liOhP:eM7m[J@Q[V=CeTXAX@VqQH_ZFbp`Um\USPV\:4Wf`U7FOZ9gnOD7G>
dc2>P7Mfh3o0OMKf<0Bq8[hZ2X1a1]j6hFAl^gEJOLFDTXq[Q?VX=lqc9\@U@pIl
?E@b@aE>J7<?n:8m3A]@:fUT8[b[@V4ZkF3P44783Ec@KHB1b]^1H0mCK]\nRTI4
InjMISFWTiH_XDmHVZVIj[7TK4iG>XS:d\qKL`9DLP:`gWj]k\<[oki1QjM2ebgF
?RRbW=86:O[VDSiQ@_lCFJSR`b:Cd;noh>hK>b8LO6M7RDE:ESB@T\6j5RAP`FEQ
c^`844iqamm1hXamPROaW>3P<D5G:ebNefYcmT\<5mH:`8kJ;^K]KRa]JHGGZ;Q0
EjF50AF2a@:X\I;o=gfoH\jXkogTTTpB_`6ZWE]3]Pdd]df?<B`nSM2_mJ\l`IVf
8@Dq1GmlS_hX^lT_IlbeXR<C3OcEQ\AQSBF6[<obbX;_dT4RCLF]FM]5eN3jUb2K
AC^91o`h^2HKTCcmYGD=TIRI4]793TA4N[FC<UmS`\mWo]oIJRdjhUnp>@=AHM3K
d3LX4c8S5W:Wj?URJTV=Z7EX;6FXEZ8Y=\M5e8E<Y=\Wj5cnD=nce52E>W5Tf@^I
8ibCRDNBO3:d5oE3?7BFCCEEb3M8DoF=UgT20dl`d]=qHZSN0iGUDonOcD<lFSN<
]4D3loll24?8L0X?7C3;kl323Gk<RLQinBNle^U1KoZMHIG[RfUO@0GO0A:AP6I]
4=pJoLkHGmdj>h?=QTD;QYVBmj[KNk@SCf]OkGGUGWY]5lDfQ>>U;aCk=jT?ad<d
e[NJYJ9C3\3bZGe@KaE\eHAkg7T3GO9RH>?Wi70qoLiB_dZA_9dc<kk>o`o\1XW6
H4c5bCoUN6k?a^d;KfEAC[VNK494UJNcN5WL=eD_oZkl42>i>MjOFU5cIl_h7c_A
KB8TWJ@<Zge:q5eggkmoaCE84nk[NEJoc`;Bi1Dh0=GfZd_Y87_OG]<km^d`S=1X
B7iS4N>CC`ZD35IkbPPCK08I=bc3D41PA>DpdBcRc9qSaUeY^H$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MXL2HT(OB, S, A, B);
   reg flag; // Notifier flag
   input A, B, S;
   output OB;

//Function Block
`protected
g9i6MSQ:5DT^<R=X1lio1nO?d^PiF<9KWZigIDJ?KDAi62oHW4XNK]j`Rn0^ij@W
?<6PhMF;B;\kJf=pk2c[8WPomWo]GKQI^=Q3YUkF3_R]j99kCG`3Q^qJ8MM:jifa
eYU4Hnl461CQnnd;WZOmg12l5T\]8gU27;685^T1SS=3638R7of?Wa>Knq^cf6c1
pFMf]TGlC_:ooNK<kMEZ_bcmK:;6o4TcAYhVk=5DJ]EC]5jq=0Rf8X3INd`bCk2R
_=39O2CU=1pW>0bBe4q?R8VZBpB@NFS[o[90LODS:FndVV>9X?OS72VZN]DJG9?K
N`ka6mf1P:=PQEAi75^V2:6`ZIBA]hNVW16Nj82N\mMKJB:W^Q8ZoL@Oo>NDd:pV
:5QlCd\[jiKLX^9Pc0b8IpUIJB7a58POYS@dP^_c21f10Jg?7H_TleCnAYi7Q>jE
X8CFS_cfig3\EeVkHNbWUbUGm0N>Pj=<W3Zb^>Y3ElF<Fde1H^[hf_H?3;pAogKZ
5;KHo]@@a^eTEdI<jU14L@TVP7XNa2Ui^CL`G1K_Qb>3e2MJfL821oN4k:7AFo7>
1BiX9M4lKKQ=c;PMYpGCZYB8XHM<D[iShCRJX=\aH[d`AkkW`PYSLFc_a_D1YD_S
GLSP7lFOgd>AF00fPoGBn5SZeaV<SBR]Ja1J`\hgSHVP=I37`\XMhmKo[5]f^8N9
P[Ge3qh>c2Id4M0V>V:mH^khAmHSL3agW:[9D@B?9V4kRlF1^UdQddOg:fM5Xh>V
7^;PSfh5ocbhAPmFKU86YNW8AUYX\0aZf439DVD_KS^jdGS;HJY7@XS\=p?C[aN0
G]mmM:SM?_0ic>jNcE<e`0ho<_g56j@E[AdMDZhI>GZhTQW;8Z<IJ\@0fC?L7B\h
O=7XcOF@MbhU^?=bp1>\cX4R2_2;3Uj3V4=nd5^B4a3aM36J__l:icWjnlbe^6@F
[44^V77M8lZdAMgU`1Ae?bh72SdPe@W:g\Lm[ST>QTm3?Z<Eb>j?[qIL[T?Q\<Se
5Y2IFi_GFAQIi\2F_6B\^mpBaheML9ak:Hm6T4_OobU]bB==QgoMQ5SCediZ=AiD
TAdg18Og<JaQiSfXIK;1bgCBdcXLiSC1f447X6BRJdET3@C>h01k=Kc\AIlq>B`c
g`K[oLn0Nb6M9mbnJNJFeG7`G6979k<Wh\S5Kl6Ajb\;U@:TBUd3ZZAcjlNj>k]m
6<6bCn[>6n0fFJITShqVB:OSiqgfnhNG@QFDcd52egnBJ;^`15ggqn`9VA8a$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MXL3(OB, S0, S1, A, B, C);
   reg flag; // Notifier flag
   input A, B, C, S0, S1;
   output OB;

//Function Block
`protected
j:0U@SQV5DT^<OW1Ni9E=MCO>UlQRj=0pRaa^Ia6\W1c@2m=TQDe2NadBOFD8d=a
f\nCO<XfC>3qdaJc_IBdU?NoeMqde\QeMq9_ng4YO48Wad`LJ><H<?>?BD\S<iYc
2J6H9G7OH7R8ZMe_QocEZnEJljMSapdA<03K3NR35cbjc4NE7EC?aW;Gq\8YR4gS
pPlCQ``p9VgB:_RQO3=3baWoPCSk^aMU1_6IRfAne[`9h0Tm]F`i?l[m:FiK_>:D
iW^5ZYi@HQ`9VcIdHUOYi[[_oe=70jL:0_Tn64S]6B9:PEH:?c9Jf>C?<GlYOlMX
;]gpIEci4W1geBU3ne6M:fDlk@M1?NVJT?3YaD^3>EhQe@@2ab3<O9VJiBHHWc>;
I^a\F0=`1;_el08<FJPU>da]neXBNN98<kYJ0A=?I^;8^ADMP86j7b?lIh^FP_9p
nIXfTJAdN5JZ:]SSn@ZWC79hgURLb0XQZ8qlM2AEXM\KC=51:EhI;2DH0G_SM5jD
T?LbeIML6LdnCD\J2a`4KIgbRLW;SH[NAj:JKK<SY0T?SCN9G23BgEfMZQd?M5FC
HZ2^P@=mX1i60o]Z7991jRQYj?=:>?qBVbF[PFg5?QbblXljhWn1M?j36>305\]b
c`]kg?]WS1iU=MG^jAHI?mUH<P=InMD>k`:>G;F4P1Zm^75mcXPPMn8O6>\BkHBN
a@YgZ9ZEFjIDG<JjQgON<@Xbb1q=;OYL1h35J2ISF5eg53SF\AEi5F=hAV>dW\16
6ZOG5L[<3LYEccEK_YQb\^DNFmad375?hLOB1F4fkI;D8X]JCDB<G1`_AqIHUAhY
0NQgKPc`:432]88NQMk]?k3W3K<De:B0>Q?@TZZEPRQ5RbHM1[5ml3RIQWoCLQ]O
a7oJJ>4ZIQ\VCA5]QC^R6_7j;2g12V9<Pd2IDMIH\onhG8n9VN^9Bf1GLG^C[IhR
OYB:AX[cIb5?3bP^4qe;6NnEIL^I`Ei7[AEo;Q4WXTY`i0nBlEYmXJ;OEngfWPe@
5k90MbP\dnaKE2<]7FiX=[FF3^D=k3=;_6:@C:RhfOU\UjdX5oL9UV3BICj@SdQI
R?1Y<n<i;@m5@4`n\l=E_4RFcMIFYB:Xa3:8h=9Q6jhTBqY[1cK@O=LZ`<KHN3YX
7YOm=@okeSeE:EJfIFjn`ZCf9bea\8Ida5DM@Lk8iQ7@g085UT13PZcM71cQ>Bfo
3]U8=KgnFJ4`@OUD1B`8T5B[kPX;SG<<oHQUmV?5gdadR3>5HTIZB7PJmSb0E?[D
jINHVpH@V\oA>ffDEJ9[`i\o8Pgg;nn:LU^KhEiBGg1?HU_1eCEP2Kig@EWl\?9J
OR3h4p3oU\X\LJ7HmiD1YD_1GL[d2CM6T9e\9Ei\6WY>MZK:>fQjJfH2N3G^og\a
H[EKA\OhcY[7TMKe^STf1LXaUc]VKC6d\@lV29`fe66@HLhW>gD<EgbcB=M1GkaF
O`V>l<>X`FQ7o<Ij[9hb615^g=ln[Z\j9plSRJcO;CCX38F>6m;?nSn1B_5jMBP_
`[D<HU<oNHG2FCBAKeMW8jkFbIXZ]?RHEffaSSJk2YF1`;gGE1K3;`T[Bm:0d4eh
jKGD<R9mRT`i>LJnPK_LgJ_Q<6Q1LEnIAb>aK1i?nAMPIfVGEPdOanHoOpOlg:o8
ofKaVLFN8Ucda___AVVfB4NfejDENIj6I6YY`G;XRn`VRMNXPVle\`i[Dc`]So9M
[i=\aKCN5mXaHOYRXSP8AVO`DUnGeAUB^7VZ`hC14o6A;Flm4M42?dG1ZY4jF9JM
`iadHNZ8<Zb>6PG\FU=kaqTB18;34g4g^I;4Ff]Ij7YB@O]X4;ckmoaS?d6WI54L
3nn=fllhm9jg>aX@8TPRQh:9MiG@J_fCmNVPLbO_Tb@g@dXTS9M>YO;fco>cN1CB
HoCj8V9@860ZiRomAaNmmTh9oZ0PNI8cV09Y7TZ^C:`?^qN\Z3R[j\T:9j`<JVEM
^:e6\9^N\KQSV<Yd^[8R4S_GQPdf65_a8HG3<@I54RG]0g:9o_`6UgEVQMGhQQm5
?GDo<JK;I`=25ef?YOBCdLccQTM4[mMj1JobF;=Y>kl:FD;bj@j6[5176>C2E\ZT
3bc`cPlAiqlM56eXbY9[KIQf=ojD<bkdXc30hnmhIGDCDc;1n>XD6:\YkgMl4e1[
a[O@Nn>64BD`h\eGIX_JWAa\B]EA6fLb2ePm`__kRqL_PXPg_1::[B2oahhFR52R
8lmP]3E?U5d?JdDTEE`Q>o7:MDJZJ7J^fioXj]17bf_ciEGSjBJY1BE]?A2S7GVH
dP0b4jm>k2m9_S6_C]^NHb>Lb^=VQ<<Zd<1<jMZ8i1PLjogNjS]mZp@ekdbL\\fl
LM9nB^PAM`Tk]N5X>=HoU:[Q50<T^<MOd1onBihLJg]\1hLMcnJ6F<J82o7]9:SL
FeHiLD`]EgKFK>kmcUOKVi^3e2:<b_O7[[<oYlTTZdBLZK?8eU]lo;K6g:e1X_][
:p[0^YCEi\55ZE9TYRS2JW8hGk\^WVQM^e>3A:R?MRTf37q6gTd4__UldJCdX0Z_
d_4F1io;FMmUjJF7Qj`W;MVeME:L62^C6idiBl?fMETa?:Y<<Q@3_OMYn[`o8m6D
Old5hF4YE@J\iUd6SgR>jCZ5CFTnM3LO6\\9k?4P<Z:Z4S2\W@@oEfZAH7qNYZZ^
f\l9od<d6G0o7?]?9S1b>?fCTB1_U<S4@QbE0W6n1\Z]PJa\GFdneSijO75oV2Fo
BYcEOB9j_J_TNomQ4]905C_@cg1?Y^e<ZlK;3m2^Y_a?fZ>iSYjKS2bmEL49^cUZ
<l;QXVqU?]:PU_e53ZA1P>2f`4amU]Z;G?Vf6_9he>YA4KDUJXP0bWd<9YnDfZll
iK<V^A3mc:]G>?Vn^12B[KW5Xk120UXc_1C6VCqf?P9h`a:7HXi@9?BFkf0e;bdh
LhT<>WoeQ8NNCmAa2MoAH^S7Co^j<f^ALdmj4\@We1nRDf8lUHLJ0KL:l@9Q75A=
Lh9@e7fODlJ_dTLNCRj8]IUGk;`XM[Ze2SgiZ9hF9d^bo>NS5:pSkXi6`HNTU6]]
RLJP`MMTfVY78dR7AAD\;a2Y>;jO`afXBF=Q7PdV\i8E3joEdh9<9mXYYWJE;3gd
f>CaWg;JA\7A8dHldT39UJ;BiPZdKNOCafHZW@6cE9P2ObZiOAnLmPIfTL0@ghq`
6_\f\]b8^:dGo7mFIECE;Nh8V:1j0Zh7]j=djlgQG24@`=[cQ4T6[<JdZ>iC0N;;
UI2IPE6=0DCPg32J20>E0CbbVb:F[\F4:eif0Bj[:^X;<eaab<i4g]2JNP9R;oIK
jgi7EH[NeRq\SkM`Vn:]2U@VC4YF44[oI58[e3jX?8NTk][1E<T`2ac0Gc2M__5T
?Agegd\JKCH<75dh9PlA4?^HT`mo9ASdOeKae8MDnbY>C1`j;e[albbPlcY9Pm2Y
Y6oaMk591H1JJ=VBKJH_lYq0D7oDGfMQoCSDGMW\8eYmeiA>jW]7a6RRkGmfhXSU
S`ql`aceP7goV9PQb>[@@TfH_Un^g5i9D_C[]Yjj]S3F\1fine?M94N1OVS3]QAY
b0>Co=8\5CR9mf9bgS;13?28eYn<g5i^;KdR6S@nDOSm0UNG0F`mIm2XNdBOXB[D
EiKi:91d2NQ]OXpBoJEL9>C][_P]1kAU11Zj5<1H9:dmV@]NQ2F35P=Tf^<ZU15a
>=XC9e[1<:iUQT^K[W^c>b`52K7<g6mS48;M]9:N9:dT^_5@=lK^JZ_?<52ZaVY4
_=9I3K=0^PPG3FdSe`bmMIFgVcph]Yl0fmUj?J2HJBo2eG@eVS[hP@S@8D^28Uc@
;Bf[BIhWEZj:Jea`T]E=o>N=BNK9mcZ[3JlF@RW[2KLN<]_Z;Ri9P>mE3;eR;BCd
BEK7gk;1DaoSlCkEK5BkT7N^dc4FUBMe??hJ9:pNXO\F2_I^d:eI`B7=2V=`>G8d
9YWFo^nGo2`M_h1EMOa;TMZRF80Ab?<`>1o4n8kJ=nEShHJ:GWUhjR0V@k:E6F=n
93PAnHi`@NZ?OW57AcmXOFiF`K3g7mLeYLSa>7bkaleK:GmU@ApYno9A<;_B4MXl
O0S0R0a8fb^G2eLLZXImLcCUO0XkFj\UF;YJTg86k`<NcKe@T=2LY>1RmFWK2nlE
WcG\H:2^dU[MnD^hmpC_DYmP^;JKU546kg8@ojZ=CTc40X`nKLIo^a5WWDJ2BGn<
858hVd]@Cg6FbRiciW=KE^RK98AHCKP7Eh02:GUS?F;4>J9]U[Wb5Y0QB1jR8nDD
ZVWL0DAJleZI2phR80hO^[3o[2i?9j]@=:RIhj>jd<Oa3TUIO8fmS@J2Y@k;;ZAQ
[Pb3mOffaQjUAn1;=CagKO1?I_lbOX0m`8HI?LDj\EdFSgNf@JdP1I^?\LLEIg0n
YPR>Yf9aUp<aSCm^4c1BlWM87mVW^Ki1dYRghSfaQHQfJnh^:?>oKD[Q6X<TMdKf
07ND=MjS:1380piG>iWN=HAenBJXL@@;<[=SScTg58D2C8ecic`Hgjj=IU1c[1f3
Z5Mm6Oj<lS6n7:J;>Rj\PI3io4<5UNWLn2@CU@:gYlbcfhg`O=L?IM[YS<SaEoPP
jmhaX<6edqE@9oJ1YeG;==M[Ia;;Vo:e\PQG2angEcL8oGXMiXomUI;XbGDRG28A
08_Lb[l37JGeBV^Nb\JAOhjUX<WZ_X>9]haGHaY;58?kPgKEIB2TD6;<DSjF;T?`
H:iTLpO@<38^LLR2liR`UG=LSZdl^6=Z3c:EUoAe8[3h1[joF0EIf3OYn7K>2V7X
=i3cZIPBFT=>cW=NXBXBK?KOfHO7QhUj3eC6q`bbn[Dqg@JLLQAi7>dgSDqAJ3nS
];$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MXL3P(OB, S0, S1, A, B, C);
   reg flag; // Notifier flag
   input A, B, C, S0, S1;
   output OB;

//Function Block
`protected
g=k@MSQH5DT^<Hkh>QdSTPbJf9B7Cok;l`T8@C\^TSiTJIqaD1T`Fk9=m@C__XX8
`2nl=7dHhANkFWVh55^4O\ok`X]A6l?oJ>2NIiZbAg7@k9@k1id`eq]DC;K^3292
G6EdfXJ1=dhD;LjKo?a4M2]m:Kp\=8OaDq\aJQJ=`_Yj6kZUM8VOTbHPFfR1MjUi
3G^N55Y;IQj`TTL6ib<gLe1g91]OSqBB;j4a8Qc]BYFQIkjSQXKJJVb`pWO7S>]\
q4@EI]Bpd=\k9EEg[SX;Vk\lmj:URCJN^e;9:EY[IiLH`c:I>VgW`<HmbN5MLa=K
F6XD>g2gahjn=b4oAVZ`Rbdj03io?T08meJce^Dl@>T1>?dGZ@6b4CM=QRXEA8A`
o[7pNTEl^`hcB>7dF1aNYM77X\9\ed7NeeiB8>U1^783<:hH0XXE<dM>4aa:Ch4E
6^d8Zj;WAe>O]G[5]1VRQOO`oee@<dTmXXi_NFL5EjF9@>enTjD3>09ef]I@3gHp
72kc]`Y48l6ANQnY0i>=81CWj<BVR5b:<@C@i6fN0jg`O:V4aod[YmaG9Q4E6ia>
3=nlABqNS?lj9>Oe?SOBkHFZVEBfL2k9WQeA>3m7Ung@Ana3A5V82BPlmi:4fI>@
:i?>RPm@S3]kmD191na2dGIimnLY7S@ZW6e9h4QefQR>G>GS?^ZckRUH41]hFXDV
ELq7LG3LH4N0318H]XTi@Q4YV8ZQ:`4aL9>BHWPjlJ5[AGSNmZ0g1a80S76WF`9>
22]Kn?>CgHa;<Og7:MB@lGa<YRBW:e9lcf]einhWenZ5lWlifn@PY@oB5c6dIPpN
6d\8kQGXbj3Q?9m7NK3Q\T?X=^nUH>YebnMda7[4]:gjiF_XjNDMnNWQ[c[HHYcD
WOJZZG9Dk<:d8jAZW7_`6\;LG6nN0p`7XWL6N[EfB2:XiK>8WD\Lihm3BL]ZM^_;
]2l42iI@WYS8_91Mg^[Kf1[ajD5OaD75S@B8`:RjYb5]Y^Va75HPiUnmFXT_\20l
\;a3AiO=iQEH4=;kP[Q:ceJkdE730Ai5;5A3S_0KaHlKKn04\I5V]plldTl<`Km7
8U3`E9h1G2CU?e^5nHeQXKNOKMjPGMm8;i@iT]=@loH1`k1=DBIe?nlYBhR8bIDK
@1oNFPk[<5oSO`76EaeB?V6T[nFTP=_INmdhB9L;\VN^O<3SgAaoE;mbgEP8hbFN
PK4C=KVHFl162l=Odq;bnhB@F_C0_MZg269`Hj3oR23Ui0QS`A1Hdnbd=b2L@c5d
oegA@PO_;;=GFE_kV``39J5\>7cId]jVi5O4H<<WR][cS6[^jR6^ac@Im?Jk;Nl0
d\UfYLV<W[iKGOkT0S`3B[Z7lVonZ3nX3@]\XmM2WpdaDMc:iVML<W>l`;3`n8d<
:IjB:1UUR4<_iURlY4jA;joPqlPSI=l2<Di8Kl3[Ng?YehZL_Y[Uf1bMEPlk4ILY
7gSJeUE3?bNLXnb61b\[7VL>\n5cP_4fWgJRnAC]OldcjXkI5fAT]1nEV2\iNcN;
Xf<JMGi0\DCZh<am7T1H39WbGeVTlT4:Z2Kna4hGjBn2omcNSOIWp57`g1NV@nn3
cGLG`L1md3JS^XPg=jX`;MD>2B9B6kOhJ=^SI7NPMJ>VVHPR2f@lILL3mC5aQ39a
0ej=dlf\AeOSmTgZakCh@_T:F]e4>J0>YJm?EUA90XO_o9MLm\XM\GLMDbmZ6Z@^
]Ckg@\bA53QNqU]TIocn;Kak_hRM\o5ij9Qf6`SCE3OKAFldF_Bngj3aE7g5_EVm
7oHlX@GoVX=OE288aRFd0?D@GRKhOXoXVh5_di45_3IIfbU[FnaVebAa]lSPG7iB
66:DSPF4]k13\B1NDdFaPHd8Xd^JChGf?HNYV7S8pNO8^4J1=ZJK_FHGOfL?kgD6
C;@8QMSie<M;hfYQmYVoW=CnBY>3SG;ATKFhQUo2o>Bcn2MBEl<BPo35;dH3W]a6
]YjT58X]nK^IPYB?:3jR8:j@a<8=UX2X=VUmG<DPR<B?n5mdgn<AdhWAWeHoBAbM
qF[<Y<Mi`bNR7MLf1kU4mTXMW0O6SfAb[\oWW[`Q9>Ff[i\@R^JZXA01<D1Ui2^9
0gBE3@G7_0_W<?]H>];MM<:K5I1]Yf3EMEIi_V@7QEcfa4W8;_cad3ZWL:m@GU1m
iT]P9oG2=l]g;kcKYKm:J4ATTPHLpSol@CD7>KSnPBce44UDEA[h@QV4L0cFVPgk
iEEUQi8I4cSbb\Df^Y9oYhG:Vk]KW:4^lk^N0_;O:ZbFIe121\gDGJjmC]lXpMb5
iKoBMb15RoNJ^gZ6ffh36ZT9SC0\oX<;GBF`2Uca[XcME9MDf<I@98EH83QBVgkI
VQb=T;Yd6B[8gAP[@SEnPm<^QIFWIHQ]nN^X3M`hm3e]c7_W6E4R^`HFBlS8hUBY
nDeXJ9BAq72U26iUge4l;L=6S@`@?1R>2>Yd?[hCOB^hEKP?bjISN?PB4;1kn>;N
BHUhP:;oG]ljI`44^kdk]4nY6B>]oeS>NJgC6bT4I[95LNhhW62n37G3A;DdR]BQ
h]g_cik;e1K]Z3D\oSEGp38nL1VPBHa0[0=4[GY@Xn_I613;JMDaHq4goodiRVOl
HES:J1ERg>;Klg]F4IMo`4ZB;hOcDN9Cni0cVbchRAFZ6FXbOe9djGkLi0f0V[9J
P=3=0MG^_>Bl?Wc<VSYZ5AKQh7NM_K\Nknd9n88i^ZU3YL]9<[ml_5NLk=U]o3<^
0qG`I:9mo?^@jd98fZdjG=UjIQ?\l[TZjJLh29]R7ccf53T895IeKgP0=:;6agVj
5dhX5Wj8hA0R\h2LN6KO9iN7ccK?N^1cA:@HXU9mb<=6cfoTakWhof_PUlUM]0cM
QW9<:>^km^83?pO6?C:_Mc?i\nWZXCSKL[2^8>6f_84i@QbT1?YZCW>N_2`9?[RZ
I;cKT=\[Zoe`4PnahJB]Q0g@k8mWReH:nOc5Fg5QV>TWcp]ZY1d:e_]lCkR^0IMM
?e9amdRg`Pf?eU`_O]0;\49<mYgVKEYAfhe\V@4b9eE5GY^2TNFKZ_`HjF5L?SS\
CLV?ShSg8C6FSa`cY<[SoPZn`?9=a>iJUjAf;k:CDDE4A:IT\N@Q7b4c@qc?a>N:
d29>A<R=5ZNnkkV^eKLnUM5NKg9EmZO]\LSeYOdkD8H3acQObm:Nn<71o:8c>VC4
ea`=NYCWA>_IXn7na97nS]WOUaH;E@253XoLnF<TL0a=7@HKOl8]D8H?2?:Toe^m
ON8ZgpW_[o^cD1L_i;[\m752S4J<cWA=NGJm1dfQY8oNMgJ0i\0TUTAWR_d?fg\f
TGVQW8hWSg7T:>BIQkhW2mfA3:XTnUo=KPioCA1P;Jg4]<Qa0cX=Po1C37WFWlbc
l5ICelWMIE7KFR3RPp:O2=K4PM]5Jnkg:k8hmo;YGh>27TD7>VDP^NPUEB\<ZoOk
1C=2LOK79;E:hI6:<TKKiF2;C;FZ?jo[kU^g>T62HXg2Ii;F0c4^@kL^lgXEXQjW
4cFg_90P>h<;Q@=d<\M>cS51JOWhIq4CGg\6_OcPfa@ckT8me:g?cK;V;S8A>mXd
iTAW>5S>Q6cLdZXS2^fkHYp?ZPWQ_640`X`D<OhSIQ4Fk]>MJGEkOK^B[fWK]489
H>>>9agJk?Q5]lDUW4kGdlg>gAfgOX;[i;cLfDFn2Zffn;9NJD=42`T`DZSMd=77
U\[BMPXmZ2glKobYmD]3\LSBC2kSCA9]YIpi^PKDRe_5PcOO8^N;43KO>l5Dd5`;
8AD`fYY=AAFYUAS86Xfai6=6;MWHC\62YnKZjCXh2Uo[C5C1Vi3@_]Pn^3ERdEg`
hWQNfAQd0T51QhUN16A1RAZ@NRV8RCWK5^5cn8CDVmQ@ilph`bT7L<j`L6P?d=PI
\oSBEj]1M3Z=^QU=2Wg4WA:HBgmo7R=6OAoLHmMfMWj@Wk?1InDEI;kOI`MHIHi7
4j7?1@1CM?Z6d6WBDJ8SVjEfo^EF<RY5JjkVCa^LWQR8XLlFc9=1LEKO=UqjTOnF
Rfa@[LT\D;C^eJ]V[1:SW_X;0@RN9Ag\RS5Cdj?<@0kBCSEVBhem1Ch]X3Rj<1VE
:eLmogjQLh3MfZ8EaAB>WDiojL<X><DDgbWI:Of[NXTRb\N8GnTO57UW`_01XW5X
KoGTTkpmQolGY_K6C[kiKdB2k6S04ZnUb0_fbUCZOI\l3H`WcUi:OQ<WNF2fVQL7
jVjSEO4jnGK_n3mjQG108JU4F^8@4e@aQVZA1pGOQmcK0EggBf`Qoq:o:6Q:^m_]
\HCJ^B]AZkoeM06g06C6]Se^9^ClYIf?I]MBAMQ>=e`E>OBFd?e;kXE71Pk]56=P
ceXGRIPAo4FV;=8g06J:eNB`5m<bn@NI335CLnM0o_il;IX5Oq;Y2deeN9=\Im^=
i@n>FUH=G<5@`Rk`EE5>GH:<``D@gLbENoAIG\dOdQMQ>RVJK67@;LCm`fimCXKk
6PV36Z3n_HL@fbZBi_[]3nW1^BXVFB7o1AN]A]j_S773aqkbbTW3ekG2Y49ei:QQ
`Z^FEIfgOgc6=AGQKT0mmZhm3LGZKZ3EjKd86KUDNf9lcnU0S1>a38diol<o8VFD
f\IKCG1gO2M1Z23k]^_FZVfjndEJT@[2Y<lOh4AI5qbgaG_i60c0Yf3INVLZAg[c
@ejB6K^1j;A:]4<k\;R5YOX3Oh<XgmTT:MfiI<TLXdO`OnXHOm1>eRJ^l7cj8L1[
IX8BnPk9bm^O3DdHI92_6=BGVI[bdLUiCW9Qcq[;4_N6VTl57JdY8oE<EK8J_>oH
C9neIU``fXjSbK8ZD1U1P\2?ROG>HF7C10WL?lJQ70Ig45E54?1Yc9AgZndLIQHE
l4@1p;Gme:DpDBQPRgi$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MXL3S(OB, S0, S1, A, B, C);
   reg flag; // Notifier flag
   input A, B, C, S0, S1;
   output OB;

//Function Block
`protected
AbhROSQ:5DT^<6Qhb\=0l^fL8>3dh>[?LWiU`AcDdl=d=`7L5Bf\CZJ9Ko9p0cYE
NoFQkdEAkJ`>aLhGnSEAk7<mY1T03?njo]7;;^chB`SgBSPVnDNNqZO9NG_d`2<G
^38N?IfU\n[9BqXCTLLmq0Sb3TXMP;ooe@jFLKHMi>9WP4g7Qk00CbKZlAE2gQ]c
fHc4^oPH;@iBCEJfqTV9JZVbb:72@EBg0GAEkAmCeomqb<K:LYgq>`kPD?qnQanH
FOKm\mUX5N=9FmC0faK\k5<TLJCZc1]LIP>AA=<i?1liYQX>;;mM3cleOCeo02NC
JCo=GblEJ8K=LIe7nV]Rk57XgB1GKogMn7;7IlCD4@_FfC@TV>jYfHpUP]\IMgjW
6@:\UjKF=2`A55i8k_@aOHAE>;SIdaCH16?\Wnb;I?bUR9X]JQifc0QXY88^la[K
DJ:3B[[fACTeC3Q=k_;?^@RS;ocC7F@lAjW::iSED[U2:m1S@=q?1c<]ZSYB@KF6
nCRFdHTRhhhQYnJNGeVDHbJNkYoS3FPa44Ej>HkHM<817EH^m7A<0PiA[E[5PZK4
RI26E4I_j[TNYEOdDf?_O0lT@MaUf>:Un;<i_[J:Ve5Jk8qSM2\19eggBP_ck:eD
E\cUlSbO2:Xf@KkHC_@AR]M2><_KJBLmk9]Z?KIeg4`N??7BOK1]U;@M^I@8_1mD
Z6oDHAAh2CXe<6`QCKbTEW>XLo:_GJNW^0I[SY8ZjBqihmJB=APS_QM_<9C0TPoX
BNG]A_HO<l00^;Fb6`9q5oCc5XW^;WjHO4I]ia\;85SMDNke:cWYGVOnY_@]Qd3K
<kS1g;CPd]SJLWQMn8GKj7E[N9o9>QXG@c09?2GUlRn_L]o`jWpbHFY8C?mS1@mj
n?0TBLnL9b2G3cKHFGUMYbiZUclUmER[eh\HINk=1kGFijdlHMQWC3h;3K;2Wm2A
OgWSY1VCObKaOZNYTH72KMh`;MklP>_`NJ\kaQMheT\=O_\d5[d?ClhgC_o9_<^9
J`Jk6653_0qn\EK6Fe2L3_cS_U4[5E0>\`2U^W:32JMf?0VF>@N8oZ`SfIZD`=35
G^1mbi>S4k@7YPCP8j;RlC0hGdcB8lWgeVZl<6fJf5[G05`l>;c^@=LQUQFF?5KP
9:B2[kI]2[Y>YmHfCe@CdXO3KRj]Ae;J\_pnL1adTeNFLkk:_DoR<e>WHR=K^Ro?
L3^h`I5Q6J@@g^kRD[[8e]YVcAF6[mQnUPM^02\]CR:_:Ub46@89bb_OTR4T0:40
ViAnb`:M@^5D2TmGZj[<in0B7IkM_A`LK\mm0a\@T^6PNjfIV<ZiiE?EM[q?jcn`
ONK0Tm_C0kPZEH7R`XCTSZR]O;@fOAX]egT`6Q^XN=3R<h4CgdHKBB^>k@2SanJd
Y_8kOjc>cIaQ]7KK3Zlc@4?Q\4BSJ=1^eRc8ZbcoLDLNXMPWQgo>>7SJFRAKa\FH
0LDNU:U296o\f>mIGCpeJF2NhQid_T<jGi^JJ\JMleAg0I83RKDF6RjX8mF4hjio
_1OFf=_jb<7jSTFV8RWUOkD\QQB9F5ogH?X06gIaMeJ4a7773::O@WXfMmbm9WQR
RCkXXA`0fB[^NiIC9M=QO\D5DFM2ABeM7dgIjVL71Sp0KC:0RYGi@7T064PoZ`ae
14=6F9^:B5?QM?_2D^LfPInWVAKDIG5<N2_U=bO@Zd^;neNM@qadRd9_[CKd:=2B
g4@DI9\DW86;GhbMiZJ6lemGVD[5bT:7XfaZD5L3AQ`;oY@OK5Ih[L<N]E6H<;Ih
ZJb2ebXj==D2cD`b[Yk;S93G>ob687S[;N2b6A[3A2:9VFbK67ohmnE]JJ6_HK\T
M64nD7GARqYSlfiNK5cHCoHXFFTT4IbUIaOWd@61J?PVPk<TjVbBL0=[=[?b4ao?
PBWJE2e;\O5\H[F0hhoEgmiFaf0IAN=4I<5V?`bcYd;fMJCa4A[jUIoiVEe<;cKQ
2`lPeSB`;DM\Y6M86UHjbZY`3AcdTLG@<p?GE0LmGn[56jHbRHk=Qg9Ro3RDLW>\
7\XSnfBBII45[[V0=^083V1;WWLeBi7f8oCoJ05n<Eh3=bohNE>FHZaAVd<RURLY
8=:4f@XB;FRhnhBMCjCZ;<RaG5SgKKLh9S:oAGO7\ddEY>AbQ]BYE]Jb2pTW74k=
;2SZ@HY75QUP\?C]=0\i[@RUcV3K]SA@QaEN]m]0Vo][AUfaD[24WKJ\@oPQb6V5
Ug23dTNJ;3PdGNL6`5E][qR54cM[k29gJGLGEShg2@YA:V:GCjJ2Hgi[oZnW?KZg
nRMBME>hkDd?HLi[W[5=g5EkS:ZMTd_P0K4SOTPk9DgF;B_;5C8o8X^fcn]0l@SP
Ein]WeY\c\_\An0\@6C102kQo\Lco125\pLhL>;E6^0o<B1J]MDO>@C7CmeO_1ai
MQ2^2WHoOe\ocVAfM@b>Y:dcY9HHkMLT]Tj9KA@R5bbRWoQ36_R0`Xc3JnX9R61J
ahgAP2a@5=No6[3CBlfT=ghXCec5<7bA2ZWUSnGIUdcWIpQj^SQ:IWI_LO@42;Jc
NJf0hq:84hN`B;a`7BjQIVP\JS<dcOL_7AQ=a^nN>OA[Je;6cISP0A3i=:?K3@[n
?1bQHmJLh:]3>7:_CU6<CnHde_Rd5HTgbBbM[2;F3lO7BK4H:_57mK^4NH`29N;Y
diOK\U<W24DM??ke7pcgcDMUc9FGjGLN[m:7FRc4[1lmR0>MZh7\IJ9>0;JSV9JW
h[0>24L\W]nG`:;a1I4<[NXT^dLgF4W`V5hl8ac]FS[KLgPI`f=l]Um<WYNEU1YI
E>^?7C`Fnmg=^X6:Y`g=RkiWK>`U[pW3D4K7>cS=oESY7mnlAgcbRTbTN7>Pj`5[
T\N3XDXMYQo[^fnSa5Y6gn_ka]mb1KU?S585PY9`02Y=BQXfZ9[bWbKdIZe>bp>8
j?6hU=j:77NNEH7U@Nc[U;eSF5E2[9SP04h;IjSIKpFT@AV3X:^F\FSQB_N=Gn_@
H3b9deg>IV_Wf57g1[8:PRP4=D=6DKH:2[ZJ]Ff7U3Jb@n\kHhY`GPfW[>R<6XY_
HFD`[B1T7CdDKA<^jJAbOiUoFn3K7o=M_ko4U_blg2F\=n1_8phF_h=hD9U1EF@T
jY3gg1flA5ZE0X5Bfkehl\[1lhDX<F>>k6?Gb^m^R@:[HYkVeYBI[Z9fRd;]o4eU
ZKEfNVHJ<YeQnHjZROOm>`SJll`l23VLUWL\Y^MEe]>f=E\Zc@h;cJ4VhpGl;O[N
>T?>KXnnOP`:^bBZ6G>G3ELVoKNUU2UKKeNXcH=`fO3gGnT1R[jN2N29CYBSL>[S
A:L_=c??^3>V\^16<Mh`bM`hReD;<<Ve1\0cf]SUUGCR:\6KQl5XE?:LlPG2ABb\
Hq@S:o9;_i0KjkF^8XQ@YT`To87elGYoX4l0a=P]P5Dnj><<eILX7GWI7bRe\bDe
`_NPRUOLX78E6EP@01Ook5]U?c2kV1O_cGaeUXbKFB3_n8VQAQ3K]`gbfQ54jV?F
73@4Ea_I_qmm_Fl;V3EnBIo656D1m8dUB91TWETE3BQT6UCPU_`^WJbfG`B0=ck]
J?Tj@>XodAdPm;^54Z`9Hm[]@>kfA5S[6XUfTmkf:Kc]QPRfEh^ImmdmUd_BfH8\
]mW1Vj6B<6mLAgOa^p3nTo6B=M8[YIf3o;HKo^CPk]b_dCVOTdU;1dEDadd6Db1K
N01<SJ`73He>?F0G[;jKF8@^A[P7D>KAj6mRG_G9BNZal>VL8LWFZM@YUEfYjCW^
4mLf<MHk^HOEZbdf5S35ORn\=qCgB1lQB:eTJ?B;>PUXSmW9k[;8Y^kN8R@h[N]o
So<MKEBR?qcKhlKgfd\Ig1_ALY;>bP9O@E7TN4NCTO3\_MSc;OnIdWDhfN=7ik@m
0C8_9UcmmRWL?kbd1gkA;mZI<W^UFS7l>kdlnKE\Jn[Yl\E@keJ8^]=7lB<dLJBF
DTBJPQ=<WIcGW9OS4q@S:o9;_i0KjkF^8XQ@YT`To87elGYoX4l0a=P]P5Dnj><<
eILX7GWI7bRe\bDe`_NPRUOLX78E6EP@01Ook5]U?c2kV1O_cGaeUXbKFB3_n8VQ
AQ3K]`IbfQ54jV?F73@4EaJI4q@8WONmoL`Y=G5Ih^:__7RRU[D7l>d0GQFBgjWK
UF=XRGSlVb\0K\CkDkhOT?XXR3nW?EAoVY3[2J1eA7:F1KDO]Id?p[_cOlMI77LC
]hXLB<BG9cHmPkPf;65b<RXFUVn@F2[2?m>8iWh_@gGP=eC\fo^[^mi37BgU@3Ml
]FAAchZ5dEhQ3PPbP_Aj<BSn`;`iH\Ak2:^S^40c]>[^0f^npHQjRj_`SLB:P1nT
ejcOcHaf1Zok]A_mAC99R\9PhUT=;`aCaHKAJ<1Qk@jEh2HhbECUi>Mh]Mbj2leG
Lh6\0^i;`2o`2Kbf125?2;IDYWAmHj9HbO2hb\8JPNc0pg:oJH>O]9\V@BhPeY18
D028\MA]01NfmZXJQX:n5R`THK=olKhg`B9mBH7L68h@@>[:77[ASi87[0SUV94h
ooaJ^SA7>L]\[HX^D\[goF2?F\HJ?>07nLHTAhI<pc]NHMcH814hAaOBBUAK6fnB
BRDA`<QBi`MdGJAUQLSClkS7=JG\e:b[X85O4`O]o;Y?fP8mI>LnAGf]BXoeYa2e
>TD5B2WRijOQ:[<4DKE5TI>nSE[D4jl2K`ejp>c4LHR[GdocZm72X\jd]2DK0PjT
5ZF<NUkk8gjK`dKblPY@jV`@0G_A]kS2ok3B]mD>;Ae:cUlDGZId0QnC>C=lPM2k
7HKqHkUf46p27a1MTZC]VY?`Y1p^QJlamV$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module MXL3T(OB, S0, S1, A, B, C);
   reg flag; // Notifier flag
   input A, B, C, S0, S1;
   output OB;

//Function Block
`protected
Oh3[LSQH5DT^<aUM`k]4YS<XAlc8KVQ_ZV6m:2YmB7lIQV9k3W_^K=FhRIfXMV>e
bJhaJe@fBgqFCSOTbGJoK<@=YFJM`NojecSlePgq\3nTRQb2NI25@:iW6mOHXaYF
l`\IlP:4iKCHg7pla_Kn4qR85EJmed=GX9P@iRJTLcd8ad>^ABoXkniHAJ?9`<HY
76Bk89`6Hc\f]f@WXpFLW7WfMkIic;2Zdhc2=8lg_]Zmq\A7`;kOqi3=KF0qheUL
9KdoGjb1l68KYB:^S0S0Y_5[;Pcd:e0LAHZlTb^AZ54eeS]PZZ?SFi94]56HCg98
OcWAkkjFA3KCnC<6o`ULj_e:69M`UO_c[nRmeA`oaI<XZ2^c9<]ed`Tp^K^^ai35
31<UmKUm=N1b;D7n\6hF3Hna[4HiVmGSV\iA3EO3_K6<oKGP\Mf8QaoXH5PI6_DU
2S0KZX1[^aeZk0aY@6EF>E5SP8OkBa:h?T65Ig106geC6:=0;20qgKVWgQSND:;X
AiL\_513eOaI]2[_IJdI0PQCHkJdIS32?Y7T3RZPhd]gX\iV6SU=?3KQ>5LlTF1\
LB_0NQjCklDV\2X6dSVkUJM>Iim3n22@G?J1?a_[N>J2nP=qO5Y\6[BfI1@2F:F]
I?hEC^e3>?Q4jSp5PBe2\Hn`7WfiDkI7FTa7B1I0G9MAU_V7EhN?<oP3L?9XJCf[
;0mji:ecZZfEH@4XSY8U=@=4UikJAWdZ1Z>@WXY?GWeggLH8R24i2R?k`W3PajlB
T8B]:XWS5]qF:JfW^HYhk2BWhBjM^KnTo[hK;8X8gT^1KLVnL9T`TcWaI<VE\M72
:UoD?n6>`kC3IOM^l>FSm1aMjE:gcfkRAOJ:5LWTMqiDN7E[cOUL\Foio;\^4QfO
G@9B3IL8_NBe[<Lod0fY0SYkGm6C9@gTUT\02Xg_[=2adOoQY5W44fVfhBGV9]3j
C64:hNOCK8A]GHR;gokHlEYZB;T?d28:9ERN^j@g4jid;eYQjZ7F4YH6_1KXif0e
_:CHAqH9TTQ:o`O\5UeKkHe24a\M;RAFVVc>\GM8SS0mdmCnELn_;]p6>`O8CY=d
C5a04V=I7cAn;XT2X5KG@kE:Id2PQm?_AH4F`RmnK8P48YAnElo4CKBNLhM1;YNX
a>?iEFaH0Q;j<C<O[9NM`<?^@I:LFM>Zh=Pn74nZG`eYYATcclibc66J8XhH;GLf
9dXUoG0j\gOAogIZSaq;6mEn1OgT5I>>m[a3BF@DDo36a^UZ;>?bj>bFm\J394_0
Ean<M5eZXJ57`1<VNIF5jmD2n;e4O\FXJ@;3fF3QIdEjHaLk^dN@3[o]i<6U5CAK
5BU\9LF@?o@4WjJ0ZVY3OF`8nSSO:Cd:?FgEgCFU?IA<4XpYUKJT<:0WK7Q_Nal4
^VZ>K`U?MEK>1Tc8:A;VL6]10dPI>:d;FC8NObCNDQD=T=3AlioKDc>eWNTRI[f7
hH5DP<kO72I12?@efSkgD:c6[hHn_8gY@@4X8m\]Qb=L9n@4QMBiDk]72j@Cj0jl
Qn6n`22_l\qS_nR^O^YofoKPl8U7c2JO1CIDBFX`Z@96f0:>EFUb1FkC=:?FdbE2
nkFiDP3[\RHe1VZfH<F4J2WQE:MZ]:Y5_1ChXF\>XNcON75dS@\mJIaohTYfKRhI
oN<:TP4o5S82XPURH]nDKjO[aTXEe0BTT?[:VCpWYIJ<`P]@mnnXL18ZU0md[_CD
bdOXeaLQ;QDHMLF150[=e6lL2D>ecPW5eM6NI7^3bJBYM8f>S[_B@9iN;GX<m]R`
ChmR2W:nG29Eck;_RSoPoEjn3[5d[?F\7S[d6TYQK9_UMXZ6Rb7=@lJdUKLeeJJg
=Fq\fjfEX3kPS2KNCmQi\EL3IkF5]C>=BSNn_ZojenVAUM:q`8_:D@63Lj6Z_A6;
8XdjXho`AMenF:ZMR[^cYJ:h@M`TljL@oW?\eS7hSKcj9B:he\><4GQaoFbn\jk:
SGON>Z>^dU<Bl:9A2H7W[l>jJC]hf=5=g4\BLFS<^CRPNDG1CGFOkGcPoKf\?[M0
2MMZ5nHYklXqmFjf1S:M_21?FleL_0lJCaVoUHWk1GGAGN0JmHP5YQRZ7kJn4eaS
U5W2?KH]4fIe5d;X@8TcMoD;5_>7[J0l52Q5GGePJbgcILIQHVeP7CMo7J9i;4JJ
@IGg7Q@]G8UUV?]UF8QA`L0_\=JN^^m>7Tf`Q]epD:cdaa:Bkm8=0US_X]]?Hi=U
]S4ciF=a6G72?:8kLmO`l2<4T39[_B1Z=b0fblZm7<K7OilhRc:S^QhS8ZH\K@@`
0NL88k`q8Bk`FNo^KOSNT\j4c:D3:4boJB8_]8FST\^Y>:>8P85@:=`Gg;7ZUCd8
b=cmRb@]^UQW=1hR;Khm[QRLQ^6^^PXL6[@Hin?L\n]nMMl6^<P=8Lg5C<lG]:ML
hiJIk3VjTic_aG3875jqi?OFL7]MJ\]ZAiOYl?L;47CFYQ>Xh30[_n@^PQI[K>f;
gd3CVaM85[RhJ2n_gTYUnhdTE14;FXhNHh6SDaegOEkGcE_?d`e23QZ9]@SR4D8j
BAdZcFm1?Y[3o>CYeWOD:dC?4TNjCe`qkjAc1IMV8?lanECIESKPGLY3j6ba5?>k
Q6gVXF5JcjY?AljEC8]T:6fH:9Zg8ISQGZ5Y=lRN>l1S@FE:D4@oPlY4RL9`XedL
aSE\mobS>YU85EV_Wc^ogQV3dNK:K0AT`Kg3LFZbF\]pY;bNgiBI^7mI1E6c<AH0
6gJOJX]9NlPF0\I_Tf]j1=5h86faI=Ik:Kn\jf@VVhnSJGJcaTZJaa;2HOB`]5O5
d\AAjK4CoW^EdCCCn^XWDYSYbL[ZKcZl8TV;XDLT\m[T698H\LDUB1JqP:J<e8U8
\@CUnemQ6@iL`^dS1YY`E2K4F5RdJEp]FYaJ?\@UCmjA@]B5k0Ge6=YXOgPNPdVj
gWZn:ID:ab4fXAROSfGYR8idV[eW>THoUGjfDlcI1IKLY\5X7mUM\=Ab:Z^]2WqD
HQJ^j;lIRmlH<P=I\MDQk`C1[=_0YY[1970WkSNXfIe\KN0Z`K@OkFIU8Ik7P=N6
<Im77J^N4?:jg7NMO<@X58[;[=8MlZG^^0ckmn=6;SkcAH`e_BO7d8^[=9oX;mbR
e]PJ?@86KZq_hbmjoQ\;;4WX2EagZaX81`0AlgWAYgEF1ib9][2F=GLN3?g<2Jl7
PdC0Ge\_na]\KLLDT^V4H0GNH5iBI1P>k4JQlg[hEH=L`RE?64jM0Q5=eEWY]MFD
b3e;Sh4Q;k9kdQPLBHM\Zhpb6iUTlk5A8:SKK6E<ko8T2<V=8D\c<0D=P9bc>g22
g^o\ZPfF:>nCZ]MbGiAHES`WNZ3U_lgVS@8l:oE:X[2?gfFI8OZ]aaY\ZKZNnX_3
PW[fO>OECX3nPCYjhePMhRP==ZidlN]U0^pT?A@Vh[jjH@ekl32Aek7RQH81KXfC
lm2^PT5HNULnNGW\fJd5T;n`>N3]4D3[>lcCWTXN<?29^]SaI>T\ciiX_Tg2KW1O
h6dkKfkH?X\0hWQTX=h:g:W46a>8<Q2hZAi5jAGEl5d0<opik6lR_9^_DeSHgTbc
4]JUXV:F;:MBS7H6mL4KIV>Ua]Og=DhWXRnmdGLEclhZhTJcg6Hc6fE@@I?Y:L=0
LCUYnfNa;:MV0lWHhfE[mhUgb<k?i0N`H_=OW_n>gj:n`[nFbH]P1OOo7`pZW;;e
i`hOaL_QU=emb4[[aoDR;E<ejE0d7>4_Ya2?Cgc`E4`4a^l3J675<hGLG_Hah0BA
U2?1]\8HK2ci]5AAoceR;EE7LM\lJUWIj?RAOJd5fn3Ik<cENX8m<faOej7>n>O8
;]m6Y3qMo?g9BP67\HkkZDC6<hYV:UHEdJORbW_UTL861^UWPN:?YKIY1Pjjff9=
F6h4bme1V;2GPANHcZ]HP=@@:4Oe0O@6dj3<_o18CARNZDoETUlM6QL;`:G^\P?L
HI?M?9B4gnPoT:PT2EqmljnQhBaMbJBLLd5@;9ah;jiDceR>ko;``V@9EgcH=jA1
9eUZb>p9eHgKXkVh18U^0OV[RFfn0IMgJG;<:ATcaS6S25>:5Z^TARkVA87RU<4F
b\WZ3Nl6]<336:435knY7T5fCkYelLd2JH0kaTj_jNkaUPXQ1>L[WGgoJUYfTS=`
QcfZ_mn55?ko:i4g`=qHo6jFPKcb\Uh\=F=>oM6C4@eVob867P^AT2=o4Fi]JH<?
0I;YDg8;ZkijXC;XQoCkRRJ0@;_FhLGKC5E3;3Coj2UEbAHR>qcjVERn047fBY`4
gcJWCQnPjBo3mOJN`DDnhM7Z]k`Qg>bn6ZMPAm6M^>jFPFVX;j1:5g9l<noE5eK[
PTB?1T@_Q:T3RI59:KMZ9PDRD9mce?;Iihi?Nk]GJO5YLq5;NfGGOSg9k[J`7h_J
@bkg5f]6V<hceoaO2;GfbYVgMn:oUYBJRC3:K`<X:FgTlm9;7P62ln;QFIj8>c=E
G<TcUD961=IMNMh\WMUAXdKYQ=>_8l\>DaWJHBlM<p:9:5e3]8K46>4_05_4PeG1
<:PgacjIWL[80n9eo<2^6jM5B:TiLYe?lYShM3hJ\]AoQN1eWFINgK[2agYlhJYK
501gh8F4@N0<T`n0LXij^hh4hXlcl27mC]=a9q>5d5>o2TUi_8N@nX5EGgV4KDIo
2gLPc=iCghC8@L[PqEniiDm6hLlNHkRQPH_i^dQ]?Gao>TQeE]B;?=;Kn>EL^QBV
a93e0`SE=<>K^QQSXFdW0Ab?_Mn>ECA>?;C`d_GW:ia`aaC8EUfmHE4j]JV0gC=[
E:;XI9Qc9fV=q`JD99MPIGGhMTQdSlPZKZkM^bQ2Ii?F]B7nljB>D;e9`I<:4E>A
58W7Bhem@<<?=hYcJh\]>f^:1TN]8QLh=bS?eN:8Y29pcRFeEBp?leM]Hm$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND2(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
5EV\jSQH5DT^<?0MSW3oglT:W9<qg\nJ1::I8;9DF1g^qh9MidIY[^^1OS:ji[Si
;;JmSl0pB\eZjDp5emWnR=D[EWkLg7hiZ0?E_6fa:;SMN@9p4T20@ioqQ:]dEnp4
Q6ZeOZ7PFLM[n[e]ee[YicMFd8M2X=FEaoFmDTWn:Z3HM^i^?7SX2W=ZI;QH9K_4
D[5BVR?`FQJZ2ll9MYqLAB@n<:1Dg^DL[3=M>RaKOhXi7DkZkR5]\d8HV<8hV_ph
Oc2\^k?ig4h4P9Cfn:BV7]ilgj;TOkLeD5eNAVLM]eV2Rilce0[_U9X`Tg<[JBYh
;a2H_d4K8@lWkki8o3pU0_7ffm$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND2F(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
gQImWSQd5DT^<CJK3?LjBL[aRJA6egb]mOHnfDQeq`^EDgHiLai8ceC?0ODq[<Pl
ojfKQLaIK2W7d;BOQIBUU2q5kf7QDpJXX[KH0>emOiL5PGaM[K_IAo>88dTK9fq`
]m73iWpNZBZn4p`hE7KP3idN;eo82Z0jQ@4<5pO9m8bOJ[og6C3J=bn7\6L\d\33
Ab<::L_PeJmWU0\^6O3\7H57KP7W[[oELa1bQbOcIcJ1?\NgY<kM8KldaqWXf=j3
>0n5OXnaN`acbADh1k;KoGKmA;B^0ho_\o1aRDX\XXZnFiWC2dmmmZIXC7W_Yo4m
I_OFb;jeS;KhjqH:Zm^j9$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND2P(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
_>:E0SQd5DT^<BFl[Zo0=MKA64MU81ZB2PDC?67@`PMGJK8bo;;[16p]ZJIG^eGM
?`haalH]1jh1[4c_L\NfkQ:iF]5PQS>CUG`7H6i92e0eYffTIeq\0SebQiZhNbge
=QUhX2=N?8oC<Ybkn7HVW9pc@0N4OqD_4XfO`E^BMaV6h8C7LLR:_RT?>Yh@SIpC
P]AY3<p1LJk>nl62Ze5^Le1LkU4BSaFcS[3pfJHoEXqK6;fOIm3FE<8eLB>i0b7I
2YB;LYTjUf]=8WciBP7f=YCBjQ]DFES;c<VV3<M76iAKbd?lX5^cEbYSX7Y3Q4qU
DKcbln2V_8]QKQ\5Y\[9VhlDR>50:>;3YA;J<KR:DIXMGim`GD]i`kHO5JOLFJGU
Q7IiG@@1;SS\FG:\D5p[h7MJIC$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND2S(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
a]XaMSQH5DT^<gI:C\TD[C0U8\@knJ<OjV=T[\Fk4TYNJN2J8bZ;i3?[AmOkJKWG
B3Gq6`dLjnid\T]jc8@:18MbBoeZG9O:1Q_71IL;@I]=>TKe[gJcIm5B[\1QM]mo
I@\gq6RCC>QR[2XSk=f_4<Gp4aENj`qHo6j^gdQF;UA>C5M_WS084MP<b75^1Ihq
m4cAg2LqQ\72L^qKVP]e@gG9he>:[c^hoPFmn\=EY3dSaLpYg63?ha^5DQ0:SPZY
\QhW^;4H8?NLFI6dL9QPUEj8d:@IHlKA7_LRlLI92:^DLT\YmH0<E]]4DeAK4W:9
o=p4oNCcNO\XKWLl71?WAWdgJMjfW9j3j>lkhA4S@i0U4Mf2oP3M@cE:MI4fR=DG
E:@4cYiHD1:9Uoa>MU:oDlq><8Km6E$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND2T(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
8QKFLSQd5DT^<h=`7m]V^npTCck:HdZe8gEh\YUY0jFPWkji\YP1gYk3GU4k?oBl
\<K]OONQ6nH305oW];A2_KGQAbHp>TZkRl>`TjgM6<D_@lCIelVdjiT]kRio8oQM
ho6Zq<XY2D=pW>7A=69c0ZQ8R?aG<^o<jAlUgb@Gn<\1qEjc1Ym\q3h:9[GqPTP8
NcX>dXj:^FM5G`khT[TjlbQ\^ZLD=Pf=Ac6TMY1K2Q_7Klh1fc\HG5Jhklg8Po\H
og:NLX98@2i>C^jp_\QQc2;X\1fLQQZjgEe[0OQXS[YUBQU;OjkL8COjkDJ1ZQf`
a7p2jl@^TZVR]PY;^4BSSc6J=0o3C6@hQ4Oo4@E7DjVSLG8P:1QT?PMmVXS\KfG3
`Cl28QaA8bYB>H9FXl<F7OqDARo<`b$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
\6aITSQ:5DT^<h8Mo=g]42XmB?gRAh0^=77p9nl1o;H]@cR2ih0<P]M_99WGB9cY
?6R9o4JqhaARfjd=fdNI0;H2bLGqUbb3dkp_TZZ;I]92gE4j0>j\OG8G>lY2^`NQ
WJM>Rehj;ep7DPL\DZpcU`CLmqEoY>l[M2`FT0:PXGf?LO9>INc_K8IMXQgeh^E?
>a\Sj1i9YYO26ZSgK5fegY4o:HE3kXnC;NAHG6o8GKh:gqOojimlBd5JS0W2k;4g
d@gjPBBF`A:`TRgRYTZ3Wm@m1MdcdWU9R`WGeOD7F;H>YVO>gR^jl3PJ^06b;bnQ
^pjAjdEc?kQfOY@3<3LnnB8[<8gj8YdKTIRcD?lB8iDDGR`T=`^DkFen4<LhEUf`
Wdj6ZL_?<goK@BW_bBn:Lpi7HcKa^SPW]SjCgU_ab<9>6YknZqoHe0H`>$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND3HT(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
5\ILESQ:5DT^<0V]IJeZ14PXWb4;W;7VC[HE@N@WX\i??]nKpcSbG=_\[>hmRmPj
]nYV`>]]0kPOOPL9Fi9X9>oD<>JGR>bpig\k2ehTm8md=7obLLYRKL27BVoQo3I0
2W2[bMjGXh3^bj;nSPYVMo]>Rdq9Y=2@>pOD]l5T8:IKh>A9A0X8mi0dQj1R<`_0
Dmn4Y53?CpEjcT_]Hq2e1b]OqFmJd;AIoVP^TV1ZNRMaJ`N;1XUA5TAR4OLogD4A
_Z2>ZnU4\b2IY?J:P3?_bT6M1FM3DjYZjiPHTK]RnSl3p[0VJ_b`27CYJ@RDY;oX
ZV;=:OPMFXVh6]0HiU[:n@lY:m2;6YW<mGX1T4^m@g<oT[WbT6h0=3CIlA0fjAhg
pDf@81SXg@_O5LTOWlk\6nMg<6\g;NiiIY;4eGFC:eHXF>lM>EWjldf>AJa]64_I
@DQlo20JkEfVHbJ5UGGoq@6A@CP]>cgV`<_6eKjR=;1L3VdEoV7Zaf:b7aLPdYef
PaNlIGU=_=T>Z;kiOR[_]11qZL>9Y`:$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND3P(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
S8OHCSQ:5DT^<jabdLj[d>j0f3]ZSmm8f\7\M]CZ3`^X751IAQFJfjoQGBaFKoqU
WXk<@YenPZO3DU3^[=6UTC<`K7I:hHF[3ZS=oZ@@Hj9P28=a?H]ETP@pSMLf184C
4dnMSj@BjT5TeZ8P``nG_5kBMi]dT0kRmH2q3TRIKMq?Ch2;b112V[78UidHI^`m
?gR@oJk\ZXUJOn6Q>Kp9H02mU7qWd@DL?pfMb20ehLLf9]0Qd@M1<ES=?@LWUTnF
59c:l]ET\g8`o?3AUXIR_GESOloUCXN<eUfQEU6kXJSfVVK[;W?Qip0aYX1\^4fK
T5^0SCNI^JlZXYC3WT8S[3@:Z=[PZN:oaA:1e>E72_VH\oSSSbbVN807IZ<;Z1SK
:La7[YK2XpC[2JP[`:>IjNda=fo6EB0=3CZd1GL<jd:CcJa<j^JPg`nb:3`\FKbl
fOH8beh`VZC]0JBk[S^GjmKc1HN_;p4A@fFak5cf6_iZ<RM8o<gcYTR=@=Fjhn[@
B36\K0@JP@o^Z7gEBZgJnSNWM9CDa50FE=BYb=pkc9LGg6$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND3S(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
VK9L2SQH5DT^<Y2DE@D4L@UX[:@3J8d5\f7]LeFTU?1;W@2gSMC8Ba@9;Jn\Pmi=
;TU@iD0E_5Elp5Zg[9ljEWjfD^jZE\@R8<`Je3MIX^aTHagg4F2KBdKI^?gC>1D1
1=hoU];HKEN=JY7][\nhpG:Cm7ImE[\PA`bidDQH8VEAnEUm1hkT6_MJK^V^4gdq
n27J8GqC_DYCa3=A:gZh7EYH1=[UF@1XnbD^lRHWJ^ECQXqGk>]HL<q<NE[F0qk<
P6@15gK[\=TiZM<j1hDDVaDo2[:8c_ME4iJn=1M7S?fcJ<L9di;:F5DJfaoE48kc
F5UEcSjFmBD3Q5];>qT]2neZBFC;i6a`:4lLMMHgP`IbhT3R4H5nTWHLWfK]2FVe
8X3OB:8SS@T02LCX0^TGQ<BA=nN;\6l8OiRm=p46[4=l=LCU7V3S:P67UbSgmFY]
[8:FP4Ag9]:_CS7J`H@D@_BH:2ggOM:l1KkFXl4AmHJC5P\UF7DBCBSm=pMe8Th`
1$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND4(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
F9MomSQ:5DT^<9Ia]lnVh7daB5`1[=qGNAQeJ><_a275l]l9m<70ZN6G<c4_F?jk
\M2Ko?fkgA\GeM>7e3N1RpHoeKI;iF`GPlB^_4f]HlMQLYiInO`;F7le0A9_4F7E
f]9P?Q3KJXWQW0j_\Te=DB?9kdG5\XpWl<RB`qZC0R_l0KBlaL1a8QcRniF7?RKa
aE53DV4@X\\ibIVX7hR6qlCYTTbgp]nhYU@p6g0fd\BBkhgQ>V[YlKbFKh9dTi[8
QhIFPl[Z@2n`D_=Hp3F3>V:Z5cl:GZ<G5m_JXBh8iiacal[Ej;:^`f1f2\oQa]P<
PhCjNg_=l34nI2NaJP;ld9G]=eZ=gQfh_DS<h^<m5mUJq:^lab=i7lOP0=BH8[In
oL\IA0:i0;FClU7>kSR4UD8:8>anc0_k<_1YEUD[<W?AO;jQf:XO?7KbC]i__QmM
[Ho597GGqR?iNDe<o7\RAgm9DQF<J;^?WlXJEW2k0E@ASmZnaaE[@h<gVUFA1UJ9
=3m?5YS`6@X7YA356B`77EfNPhFdJNZHZ]B5qU[C;oP>`B2Yffi8;c6Gi;KS4Y]V
>2oFRKV:6MGoeI>gjh\2g<<d=5_B2Oi_kLCj3[mmiYd:XG3J=J\PbaPMV;2EdlSK
pQNeS>Je;J`eGE6U?F\TUdFnqTK0eL;=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND4P(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
5kO7hSQd5DT^<4N1<\YAP7mYYXE5:3k0dAJHIdP5Ef^q?W3WO\CdUBf_^OkIO>oj
d]Fol8N^;bclOJ\1K3?ZMWZqE=\gHLFOlClV:XMkNB:=hQi?VTd;=JcB^34352\h
eGqbio^C1pGh6HL0^Bl2>NVdNMl?_hO0Xi5<nBZU;YjM23OoIcjFHm=dqIRM5Fm\
qf\:?fGq8dV<NFdL26jL_P68K2>FO7BPU@N\JF6hYEn_e0k9mh_?DC]enGhRl06^
k?9jKid=2[fS4c4RfIZC7FQKFh^EPYSjV_fq`]1A1m4omBR@X>^M2Y0@<[_:hF^F
<mmiRnJU\j?`>^Kf9JGL3lRGcD5[`kCoDG5=;jSb\1JJ10k[OFoNSS`gVXDi`W@p
8e=nRXaPS5:[Q<AnJVG?V3C::3Tf2EDBiN3n\X7Bil6o\JRqL\bYHII_`9EeieLV
Bm0TlPn\8aO<An_a1>^hda;o9DaZdRj93<B^^R5QYCe`9:V@18YZWTA^CPkebLcB
\mT<:kOUA8Gq:CKWjiJJ\BGDhBYHGYRY3NBOQ<@Ui@N`cX@1>LVNiaCQjhkHkZlc
HfV@2TCbBE0KgDkJ9`6XC\dg\bj2k>4PeQSJZF]q:5k=OY<$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND4S(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
b8Jb[SQd5DT^<05Yo80deYFoHgN8[Gk^WZJ7Rk@[o`?3TXmaWe<f4@MHqo8l:V<m
P]\H2WYNK^_FBYc6HeJ;VnHCpNG@lKibaOQAa:H1\2i>`eYBnLD[CcgV`N2lMTV;
Kh6Gp5gK9Ejpc:`NY_fg4>Ch1IMb;E;UlXWL8Q[k9Qgdf\:P?@L>E4Y>AWp9KQbB
gepbLlFL^pL`NTiYMc^XZ1\Fi20ZDEBb;dfC]8T@E:QNBm?J51n@1Z;ZFidF6\43
f5^DNOI`:[Ll[dOHgZl_XjVJV6T2@qFkH^^3]H\cI1J?lDn<RfXTl<DlmPB[1iQ:
4QWGf_Se3n:=Ejg]S`997JkmoINA8VKD^bCk\B16Lf]Rm\^nP[HhfqA1^YhmmnVn
d;MBWNXogUCKBMCga4@>ib;_mS=[>1`GAT?khaA<j3;nU07_d>hHl<R_I52QIBH\
79[DhaNA5640gpH\Lc?T?<dA_;hmQ3fAU5iC^N9DK75?\Y2^:LR=EK3IkZcj1m18
^0OOKT]4aPk1<Ea^NQZoX9HU2GWcdRH]5fP2LjW\6pPO0>5\1$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module ND4T(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
nkKB9SQH5DT^<\bY26MOY6gVADE0R9e4Efh\6V3<2_5>TEi_3E^le:IRPcn77<En
^aXjJAqES@=c]\X=Y__I^lR7dPNWcWKd^BG25pjk0k6m52KIko_Zm^0ohBXCZmM\
dhdUK3hG9=Y`2>nI>pkoilAmq5Z]9EQ]MdYoiiS8Q[JjadOmoBV9_CCBD6UU9eY4
GN^c;NmqYAV>MIHq:j^?dlp\j6mfDnVZ:;_gA0lDY_GC1k3Ea?9\;8_bcb81EaUB
8FcIoEgO]ZPR`ZMjMPT8]_:W1CSn<A365:4aSc;Zc^VC;6pI4gmVO\<gen9ZB<H:
a1nNcYU:KjFfV:FSUoQ:[Ui59:dK[WHG=n@SUYGS6R<`Q:EiU>l66CdWS]K5ihRQ
=Q9X?Cq6V[Sf3GMI>IF[PbTbV[jQ8b^Y@18WFHARRF>@683a3cX7g4YW0N75OoQ?
NId7C0ZI\]G]hVnRY4_8jH5@VM`ZFDkoI<qo2[^3iHJEhBHn5g<GJ8clPVLf69j:
cpN_8nGVfc`Og^b^ST^3TcU8m7gNTn=IF?J@\:LSDjWX=dV@<3X;jnYIVWbI37K8
PIL:VS=;aL87?BV=bcgc6_X66n[4Wp3^>5<6^$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR2(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
5[6]OSQH5DT^<b7lL^OdYXSLp36mX4LcX90NP]<CP[3<^4>Ubm^b8eO?gpKVR_e;
oBR@>M]=U3T=pSNnB_Wqm]1fD[?Q41WW_jn9I:lgTUiP=nb_DN;;pQcfG3JHp_O]
WjRqS1ZLJIMCcM8of[FhBemHb:Mhg]:<5;H;V;iGKD^MEE5LC@`^Jh<Mj5QfZEH`
n@KISPdJk4:n3MQAHKbD2T>q<AdEa06`5eK^5Hgg`;L;WJIKTdGSok_M`eH<OL7<
3]o:2Nj\FIF0]DfP@HAL9Hmj<K?RjY3SBdBi0c7OA;mq2QYM_d`$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR2F(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
b2nLdSQ:5DT^<LH]HK>9>ih6`K4><Vj[3FFD1Pp7]H;EQNQh:LWN_nad;9U?ILM`
ab4hkh>\lVD?2IX46pZiVRmCI:=EFYTcQellRVKNWHceZ?<P<97bqC0lc0cpg9Q;
Tk9\I>E5Q>@VhHA>;CYbRi8B\o>Tp<n_J7aFp<oU7aDq9SoY0b3lXFh8ilKVQU]:
kU^djLl6K69ClmkGQ3CmoN5?11MeK?3DR;X7[aG1Z[Vo9D<:YnacmFkB12mAgdBp
?5eCIH[5VIZBlOk:Wn;WV94ZiHi0:V^W[O>lNdb:0=ZS3RPA[mFENmlGIl8O3\Ln
?nNE;9CK]1Y@\7YAk26q?4AJC0=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR2P(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
D[_k2SQ:5DT^<oLR4TT=6G^A_;jgWWSFUR8M?`NNI]Bf>YV;l\iq[<f=KE<NjXh5
X4amfCiZ]T\n_\NKaWZ^J7JF8[NZGoDZml=m>9ilQ=N7GW\<XIS>M`4Q28q6nimM
PO__C<[n?q<9?4ampQ;c4[@jkN2DY:Qdg9j[K8GL]Y2XA1a]CqNjMLG_ZpcYIZdK
ISOa34@>XS\[NSn^Qa4V@BQnK60;Q5pZ?aJO1q>gE0<:V=8nUPENOASPQ3d17IGg
YMO=2RA_:JTmR`EjaoPB9ih5ASlU:0VK`lB7oJ>I:_]=mK?F9JSgXo8FdpJ0AKkj
NE;2\T9cj?ha88m2NML]@:Jk5NY]]f5b[>Qjc5kLQYH=8ejD@Wc@0lE\V?J`fdFL
lc=RChY?W@1L:qIH@f3cf$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR2T(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
69FP`SQd5DT^<oHbjee;Y;BgLWF4[jJ?U=VN4L14b3bkJPIOQ<1AA:VbRbMB7YEG
pL_e?<gUbA1W85X4181C[QJ5K7RmTO][I5iikXWl403bV=oqVi8V5;nD`GK6ndLJ
<fi7VR0X4aE>5KG1\bB<h88Sc6MLT1qWgo[h=pSZnKUkbREH`?d925RLPRXHiE<h
ghJgYQpXV4Zk9Tqg1Uh9mpnM\M`B1GeLG8Eh7Ni6_2IdiX`daL1ADC5Zkj?__HbI
dD]l__7UfWb92Re44XV91Fnm<E@e19nG]8d]0bZ`lqiIDY99RIY@VmKC<N[HZ3Pj
35F8NIjD67_[ZLPCh8nPbNoESJh3LYE;a4KPSQTSigiOHH:G_h_lFoT3SGSLIp<f
DS2=`$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
_9i_XSQ:5DT^<@a]R<[NLYD2`1PNi5T2:Na\U6\XUSRU1d3bKegi9>_R0]MD9I@8
]jGhijF8B;\kVnWqKVc```;VG50DFU]CY7<Ed8F8Cbo_4AM97aPTHPfZjl\UpOMl
669<CC^;Hch5i=CYIJS3DRda<=hYMp>0i`[Gp;IQnkY<k<5iX<?OR]Q>Z9\ZHj_D
6jPHFTK@cNahpZC?`iLmqQVOjASp[nInhC2I=HDY_PALiIJ<LfeW07ofY]CDcSk=
k7=NB`4E=;E7qaCk7S\cRm:HNk7>kIR6h3=[ihCD;j4gWkd;@>l?ZHRa[J_?ISJU
a64_LF\13KFK@adH5=Gh_djc[n09Qfiap`F1VX@^_4[_cJafh2[5Ni3EVP7R_?K_
BIGd`i::0C?[0[iZf9gh?Nf=BVLL^4ACj`ZK2lRAkc796gL98@BSpe8:K:<ZQh]E
3JKKSR<X>^C6f93eK7mD3T^BH1GNgGPQJX9YI[0UO2>I^O\FoG6A7eA8K?`]hcma
9oHdWJX1qL<D4ab?$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR3H(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
WQaV2SQ:5DT^<^eiNSWO<IP>>UlQRd=0pFlOab:l47j`b25flo@c9pm<QXQ`?M4T
OC@SGFhIk2jYBOnUZaaReV3G[OSXA;EK3f`Obq;ojQ6kq<fFVe\mCR\?Hm;geG]V
VdT@YGWb3JHZ\B_^?mgiqkgi^=QTqj?XhnOp1FjM=L^:=59^cA\;:h@H9LJf73\O
aZ>RCoDO7:BTbGiA@ESkWOAMT4heA368NX_K1`3<?4naIATXAJ6a7l2qlmgNE6P3
SF?7Z0daKS?Dhh]EYK=WL9^9WIEgf_LVooH=8B2oc=DU@QWB4^4if?ool8kkF2HX
bn]hPGY9f3Sp]XHSNm<WNUEfNhIoQgk_M\88C7[N7XlbVNJ]Vm9_C]MMj?N4fMfS
Z56[`O7cUB=:]Z[1;n[FDbdfdV`jVdeq8S=J\ZCCHn;f>]G^8iI1JI;1>EEk@?k6
N_BMlBb6;HOUObnB?oYPEUb`^G:@5R=0cmRA5A?oqc_2lFP=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR3HP(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
YkGd2SQH5DT^<B>XhTcgKL2aLOUQMGoRefa=?C\^TSZj]Ip`iVbMOgN4XM\g3<XS
\_gC?Z0C944^X]K^3K5@oI9M2Y<9U4bLKA]bX409T8q1c42^Ei0:0U2[LE2>[f1S
F7MBGVAF>AjV`Y\NI=@^l`YQeY703\[SX9q3?_;fGqaRdS=S8<AS[5REbOo02d5e
`WC2eN4926Wa>bKiApG>jUa4bp11^kZ^qo1>NJ^XI9lD>1cI=]imFoZfqEV[PD9J
U`hU`WW@\Z02gcG82G=[`A4>Qh^^No@Cm[Lho0oW3d?m?Sk>C;N<MEN<=EYcD[>A
W]<J:aSao=PnqZL5WgJ^@D8`^K5N\`omcZJ=3CJe=MMD>ln=`MVgC29gLAV7NJ:>
4Q;5mU?QDbFKJZTLgCI9K181F<BOC=E[qPRHJcDgGiPXCci]5g8a;INE:m61EiXc
5g@deg3UeiiJ0mP3>0NfQOXPBC?0Q9QGaP0N1;m`fU@KJM_;@][JpW8JMhn6$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR3HT(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
YZBYNSQ:5DT^<k>:=NR5BIh6WVoYNjj>`R;bMbfFR6=?aWfkm1foCZJ95o\p?FOC
Ql1MUZ_j4a[nUA\o6=oJ0e:<Ec>4D:8b[]_;gK39M7fimoZ:F_A_GQ7p`;QLNId;
11k`eBD_5gbjhH8JFSU4jISbd]m7``4^je<:aG2A`jKZ]898YePiU<=Zkgpbl\G^
lpbW2_?JjgHLBN_NgAWT4l?4jjaZcM1[5ZZD;J2aXp7FG0h?fqjk\77UWXT\i@OY
i]R55VXY]c9<ol=YHmFf237`=^V5Pe>S75Y\a=8dKB^k_^6MC??HcYl4poDF=c8q
o_jnc_fAOQY\a;?X3VF?Bg::aW:\QJ^:YgT<F7<hj:I?Z`]G;ohO^i?TDCHQhGDD
oX^MlG=2f4FM7dXh]ETqmF?VCdUY6Y0AU?I`KPLCSLdCERY1\`0]Mg86^3Y0T\b7
CjHN_cbggY^]@5gb5gdMmlSFKhf1TYR[2giE\[Eq9jLYQQ@`R[0123oDZaJ1hn]j
:=7PGn6_9Cool6`3<_3dJNqG9;`6;@VY`G8dHWiDI\;PUS==OLj[W0X1gYW`GW^Z
YI[7h__GUh^S>T61d0E4Dl6GIHcDah<0iL>j>WN\2QpN9hOQ]m$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR4(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
1F;A]SQd5DT^<QU`TA7IoRHe8[U_X8:\:6kS1P9Mf]F1QSQn4WX0[E@BZIO5ZaHD
VJhRJe]NlgqUi=PI0n_Mcfid9@Mac_6?E73i16hnFUX\9^4IU?L7GA674NXqo3Ch
Qi=aMSXN:iQLiCcW7J6M8_cBcZ=hGg0Cbn9NJKWjZJ<pMWSF2Tq\@S3IXEK5;KMS
RVT^UOmX]Q:i_m8=548U9k_SBL<`;?=1CpoImRRH\pfQSSU@pjT71J0_A;6bYiVI
Oj>:17OSW=Y_Hdk`j7B]En:\ei2Zc0NGV2<=9>O]kBf;_jT3VFMP79KV0?XND[9f
lgaeFdanq<_`bZ^T[P>flRZB8MYaY`1I^I58?X>@AX;74:Gei@9j20Ndb?@WEPRX
gUOjDGloN<\[hfWR@gdnc666;0JWpb1oH85NR8@Ph8PIIa4F4a>oMHGU5@OVIU<B
b@?hN8UaH7H:jZcfPI1S>fPRFPbX<<cbI]\No^>k_U1o^ZS6eEE=dU?;p?:4fFiX
\OUd4m9kKQNg>Am1ONRT_U;=E3_nc\>Sp6Xl4^Od;OB\e?N:0QMYifkTe;^LSJVn
og:WVF68_kmGBUVJf:9U:Mm=h7fNFBNXC?6K;TSXg5DE1Tc1Ui4h0ZIXp>lDS=GW
$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR4P(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
MNVFLSQH5DT^<KeX9V3?glT:hDDq=^4KSY3h_\dhfn3Q;^DZe]jIF94S>SRgC3=M
a^0HN7k0qW[F`Dd;Q1XcGo8nJlQ=Jf4c5nj18QLSN>L^^B:U?dXaVbZ@Z?7D=L^q
9@iGXjphKAm=7ZgBF>b>26KV8B4A7<On1]GSJCETchgi^YH83K?=dqbK6lCm5pfh
GXJ5OF9^4Ue>]3aALD8?L2pbl\G^lq^H`D::fIeAiKl;fmgg\3CWN1aVHLj;=oId
H?m[39RZi^o\794MC\8Oi9\SLM;Dj<o8[3]GocaF\n<J<PK?G0jVhqUOO<AR^4G2
cPJKS0gK^HEZRjmVT=M@kE3>]FlN:\mcU;LY37@J]I:4dDfW^@V3IdLYR5360D9U
>oH?j;PWEgX4gp>@jNd0a9o9GZ>BBFg2M^R?kRe5I?[4LdAQl`QF]Q_BZGk>FP\1
@2Kf5?j0bd;K1[?m3mL@b>0CTXDH8;`P]B?iWInFfp`d^O8P06TPlo3OEVai7R0@
;fMf8Lj?DE2CQTKFgMUZ=C8LgT8P2id9UNIfDgo[d;`hQjWXRhBlCMEc[23NgLXW
QqURij;8a$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR4S(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
ITnFaSQ:5DT^<`>H3d?S7U4ERb9oSl8UmOHnfY0Aq[nljH;L>CibBA4\:FL[`>SV
HW4=@a:RD;1_48h1q?0B4h<2gJMO7>;4=?gKFFhnQdJX1ke<WO1QS8W]Y?U:?NbX
ccKN=WB^bBJY^2XpB\]Db?p\MKG@h=F?T<1coeV79TAn65Fo]2J:7Dd9Ma3BHGI6
0@b1^pcIN_?^4pA6bga1pA\732c^<T>:6X89ZK<Aa>LcQR=U20meYn0ae?ka@B1^
Jh?NilRkOQTW=<D^h8]ImEKFdiaLFb9To;IOlDIjJRn[pLee48;?4Tm2iXj<QolF
M2Hd;@jHgm3Oi[EjAMKV70DQ1]W@_0iSV?Zj6Rb0^AO=lLX6O?_7mAdE2_IFa_Q3
p^UVSB9`oSEo=F1oMNG2n\[h36]6ULOmU@3E@2f:IWj6S<jQ3X^Ik1N0IWdACJbo
]F1hITn7?j1E7N?DePHAi?8=p9]]`6<?89]R@YcmoODRT]U:99F5NoIG@H5cN?4>
@iJSo907SeOhd=fZM7XVbbY4g97Tm<BP05[M3m1Z;]JcpK1\PJBG$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module NR4T(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
4[^l`SQd5DT^<cJ1L0c^9nQfYi7D>1P[;2V9^MgRjafZ<K8`o;E[G6qZMNHe?Nj2
iM<4J>EBhLnkRAhUdiYQl:AQdRKj8WGq_Uh??l\@_<f=bh^D<Zhl3GfV3L=bc1Z]
cLPAS`a:hR487[@qdSO[Xjqj;bkTQ_ZQOIU30C=LjLn]LTYAnlVe566Ig>_GDlB:
Z`MDdqbh6i?DYpO^V5E98W^eTGDfg;WKJ:COH74QdBKV@5@dqVDEM\1poJGg<Mne
Ta[mBaDPBoQ\HcFhZGoET5=`^2A_gEA4GWeeYnAG?^kH7UahjQPRi04RTnHN4\[=
i\[1``Tc;oVoDHZBa?GpOfA7G43NRWZ1KMmS[b91[VbcFDW9ZfHW6E:hU=IT;@8o
8>`eUl<d2I\PFokRkl6CPTcB;3>9MR=F0JR51L=]h`:;03QqGUQ2]J`T:21gPhOl
;7n_TfRWUeh<Vg2N>[00l\@P52AAgd6_8QD=ff^^=TRi_=VJalYCiiUJ_ON9Anh0
oohdI9iNXh=pgad=DcO^jaCQi]3<l1KB6SOSG?ZFSoQ04gikV?k?ccch4o1<0kV@
8\0EJD\UQIHdla]VBITMTZ=]MT9LfCiQ6hAl5@`pP?@Ki?U_WV0=NYaJm<;b;_P^
9cHM8=nV\hXfW3gcE`E_J87q8>[A[=@$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA112(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
bHET2SQV5DT^<FIaB4@1^M;bJfVUa_O3M_hhDimRV1Ye1g5BQ6ZZ_J9aVNO8JKWG
56Gqg_hZ<0W7DM`eV9ho0:9ne?IkGjX7NJhn136PY:KhnJn8i`B6ClB;?b85qI7A
m2hk9eGZaM27[MJNgkK<pHP`?2Tp9c3QUFHHHEfeFN[7:50in=3DdEaYV41T3XqC
TT0adg5_:SnGMnY:?F@5X?Fle2j]TJFYk;[XW<kq167WJe[0heaeN];io<dMJLGU
egqF_C7l6_p3h^H5TmVS\dVLT\W>5EAH<4c>2FC5J<68TSQ9nB3_dJQ9lHSXP9S1
;pb9B<bVqC0@^a_;UdcjMhkdjk`i95N=_R;8Q6UT1NBIgSn0oIQm77IEc8oj^S`1
YG;6NAf=XCjmYNjjcoSJ]34;_0E5<d`OkPG74M\@JFBFG5jaU0OG?iITbcd`iJ2p
g1@>WBf4L`i6JldG:H<BiC`ZOT_hG\K]39==oLT@YI9joEHL[Qbi?B:m=CgJK<]l
gS>VTMN`Y2HT:jXD8Z4YSDJ:lDOc_]aEI9==b:348=MJ^Ro6BkBP:4qeR`MZL55=
JP?mo\\84lc57UTYNC_CU_R3A;FLl?9lIh3E2m=`>X>AUI[\cC?NSCQe_CWF;68W
c;U<;UFGgSbBo@1>HM5_;^:OA8]LUP5T@MVJKnRT989?1qmlOi^4P40kk]UKTORh
N`0k3B1>1l^h\GFSHkfT\njiQEHPAJQPC[<XfL\FHc\T87mFcMOY]]d_X5>hRY4^
T]36qhTS?^YL21Jao[JNYc@ZThJLQdK]DaTUc3ieDg82nINE:l61BLX<U=>GSUIE
=4UiWh^HVMj[b3JkVZ=fLahGeVo<k`GTmAHfJ7ib>jVHH`8INiDS8OImJ_2p@XH3
m2^jZ5fJE[Ff5iGYYfV_QB;EVhD?l7[B;RcR[5PmoU6eEP3C?:2::k[1]OiY@k=D
S9XcbBicjD`4Ff\N<>FDZ2=9nG`Mc7Ul>=0WR;QhUgZ=Dhmo]lq^A\fA@]iHb06Y
OpGP80D5iG]Af87?^GZV:;G=:PLl1TGPWA3EaFhRi:a?E\GI0:dlfAJNZY`5BFcV
[JGVYTV^oO>O;6g__JalLa38ADZS`X>ggR3EbO:6di]68]]1nPM9^I2Dqnc`7fn;
H[dVbo<Nkfn@:lZPooU2IDf:?P9AW>8WgGK_FV[SbHPK[@Cf8f1CTI?JLn\;aRN<
Mnd01=f:VT?Q?5dpXIo=DBqnkfaie6OaE6XcG1]\?BSoOAm<`g2AR:@F`eam96E;
jK]F637m@Y9El=BLdRCTc=S3l:BgTETDFI4Dh5W@:Cm6NdqPQ1;gBZS2;7CTW9Zh
IHa8:]gZ[o8\A]@[8hlBCl`OWVAocoNjMOmQgFMOP>CCkU1KLGc[9PFGaFQ7kgY\
2PGCR^pTNO9bcT$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA112P(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
McaVbSQV5DT^<h=`7mi\Tnq:d0YNI7RWd>RfZkbLAG:Y;c7X8221=Jm83M0[X8UJ
RFeIVJVlj1_cNN?^nCVejd4YIM^pZobbbAJ>dXVEEnD7F9LR1hU^Q<KED4@d\BNJ
pX9f54OqSX01gn`26?\0:[99_<RR0TX:b\Fd[D?aElpmL2IQL1ic\nl4bbL:=[6R
1Mj6d<>ZOdLoMdhEKRZq7LG3_Yni;2bgNITMBaXNU_VJDXq3nRBeXap>3^:4?poT
6RkXTdNIBOM;W2Z?j>b_=3\g1`N7pj4P238og58X=gcO@=c^NjAA7dkPKHb3Hb64
`>ngGQMeXlfhbML31ZS5?CaWAd\b_jn72h7CFcRWb0Y2jjH?9?9AEE^g^<l?`J63
`AOVIh>;:GAPMADMeD=q_3853aL1?@hCNf>j^\B?[2;Pb4cAD_beYA3OnJgJIh:a
OmeU=aBTPBOclM]5aDAm_AHdWGfUP:9Z@>PG@Jo0N@0Y^Z6CE@5j?Agg^XSbeTR]
Aj`;71kfflq8l80R>ZC;mKYaJ6XoJ1co\=:mVVj<d97F5N6EUGJ6l81g3Go?f9Ne
FdEP3cWZY5_8WD0k]5BWNDmc1^1AbDoCjcYS\gZBOjO?5[Q[^6L?G?cREkIAo[2l
1q?j:2fHhn0hISBjhJAG^3BTZj>jQ7QohjJ6n<8>D]6JTY<;[<7LfZ]L?UV>HWKN
4h?e7PL[hkD>Ml`Q\NX8\09CpVQaT3k=5D?5<VeFT7Z<]7B7VPgD388e9Z9E_2G[
9`[::^34NN8<^7eLU?M>2XUH2V\U]Ym;_NZ8:@XOG_gYGk2Qg20RR4h19U9EFfkY
cNBRlFdC]dM=4L?qP\3mL_IDReE9oi:`jKQMa<FGeQ2^ZZY@mc[CTeX90U^Qh_o8
4ok_ac2ZBbaL8G]gPEcmY0Q3g@_fIgmhn]C4iZ[8[AaVU1lKUcLiLlh@mOb7La4T
i2MQDSq^f68o?ADlFk7fDDih^@70iZXc[Sf8n?Z4;_^K`TWbQ@=emMEYHEOJ3P74
eRgn02P^73jQb3;O6UEY?N>P?94OW;hOEfPHF1fQ;3J:\lNRDV7=@iEQ1Q0mVq3:
F3>K1nnQVA]LX8?DCVA<MfI_n1VI<_FnF`m1l4_fm_l7S<U9DZmT`I2a^Fi>_<3U
M]7cgjU2UBjMZ@^_cb2=qP7Sfg5a=l_7h4ICic]V6na9gYGVj@9PLoJU_1Bd`i;T
nSU];^E3DFS=ULYlecEL7j5=qmg5F5Pp3PnOHbf17;d;QH[kUTL`J65D^TcbZJ1>
a[Ci;cIW95\m03HSGT:aXhn_5W]k;9BOaBFYWK\fj<A1m?co>ANLF00qHECk];Vg
PB8KmN=HNX>Ye>8H?8VYZ>oe85hS8\OEQMhbHgTbc6]\GVUeDc9>lW@hZUm0[fC8
nLA0?P:N_V_19l_qWY0bEeD$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA112S(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
DSagRSQd5DT^<H5i^0g9k`PgRog_Ah0^e7hq`]ob=G`C:9BWHC2]`W`ULD@kC@oD
]eQWZU76dPPGkLfNDfBU[d5SXjCV7Y1qYCFVXL0L_Iaj1\eIq>8]9Enp2PZLK=eM
FWj=TZD_T<JEEHBXRiAJBUM2N1qQ>@2COEfXPJ^[=ekBKT5c;9HH6o>ccAb_LZO?
Y0cpCS4c<iJdJ6_OhKaYNOci0Fa]bdqneGBdLfpeNHd]D\516=IiR^On<Tj2YpZm
09LWp7_3j?BJ526c_\^KbFmZ6M>HN1a3m@PnPJ5<PL3A?92`;R[DLh6@j3d0eY70
D4@037GZSU2ZGAYZ29<8FO_bkQBhLh>2DXS\\j5<0FhB4`k2>04>e8o\IfPp<n]n
mllo<cjZ7R3L18_22Ia7NCeT:j@c7fCY51A1VV8NiH2oNL;3VmafLK2bdf4J<M0h
jco3dJHGR0^oCT^G>Ni:AR1QVQnD=fCgdZnSJU=Lai@93g`OhgqnN:UQZh4oa2N[
:<1NO;6QI3GW4TEUHa\DE1dI_I:]7XmOR:0EX;F?T=6UVo@WO7encUODaNl19a2U
Vc>0kd@22fFCC?e_549YE_jW=ek3eB7\ce3]BJV=VpH4MU;Oc:?hD9[A9]:l<9lI
h3k^mKE>Wg:CIb8`1:D0Ae^eG_ARC72iG>5aT`Oh1WH3_IiTW<S`nFHk0TQUQTX?
p]eL0;2WQGQdjKeodco[jIXKjL5Ci1QlOKNkfMHEZ8WCTd;F;jWnQ;hCfUlHN`6@
U]\LSLV;]9M:2l\5>g;VOkAcl1[n26ZjjJNHjNQ[CC[2nhk?T4R[jHJqPh?UlY>g
;fDjD9?R;l52\0gmU]9IU?KNdmXTThN;@E:V4>D^8kd6oTRA8OXLEXG5Pk0OYLlZ
PKTdb[da`GeUn;a;F?g6NH4=FmO@`I0l]mP<[`SMACMo@GqE@PQ3o^XIa;3;ia\7
^ZbAg\Z90^?LU_>;F<lKiG9`Tif4=;S1P>QN_c^GR5]L6i6EBX61Yhj>GLcXcMBG
e?DO_VEKjDQ2m?o5FeciYG?1[P6TDo5Al?:]Cp21e503M]3=`N]SL7^m;2:@HHek
qVB\8R__KYVaBZKEljMa:j;=U0;eR@cJHlo@^]JGSU=a1=lHkD4acT7MN@@m\KO@
XVgLTHc7H35PL?G_=k=BoZ;q3BIJKPq>Q82aQ_F;CRQ5J[36[FfV299Qe5V31OIU
Qm4=Pb1Jg]<TJ3XPbd6cB<j];gKYE5FH9gFF_R03m5bP_df=l@kEo7p?`<V=mRRo
_5Mj@mQ3>lKQHRm5VeAAcZ]i=b<8=NMX`jNAVebhQ6j:gOb=0[<<XL^c;B?HE:l6
\1i@N92ZW`f;E>pkBK2mg6;n0U8n[pg@P2iek$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA112T(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
YQ<PhSQ:5DT^<i0hV2HK]_3aWh_>PWXmCiL_9D?QX\i??RRKpQ6ZIgn\ZS?6b4g>
bP=pBMA28F>L=63V?EQO[foh;7YUTbQ\n@P^CU5imC=b1VMC06NTp974l7?pA`an
:N3K==KQBmjUM`i0ALg[oEn1;QA=c^qmS]M8:<7TFoQ]MP27@A?OlCP>`=R6;A2Y
SUKOL@Gp\TbhNR:im1>9E>TYBYOb?67>QWq7>D>8:7p3lDm]BqIh`0Tjfe`hR88`
RJS<CO280XqhV_kiK`>`GM]gLm[?]78e`[^FooQ6FmK6?Wk]amEciN;]fOGgBUOK
eRiOeGg?eS[YCXJb90WAj4a8C>PQ@n@:_AG<TUbe]ZLeBFaHaKK[GVCR=XlXM2[>
of5FPpA`I<J;So]WdoKe=eLMbn;YT5GS[k0fW7A>>a09Mj]W\\2?]H38;C_;UaT\
P[Mgn4O0TP>?KdRfOU_lmZF`EQXC\Wd][SJBaIP?P[J9NbKX6KQlkaH^<=^:Aj>a
paKCCN4c^GO\j<D51CET]OX3T<lZPa4kS7f>OBW;492Bg<U<SK3<n?^kE`Tif=>;
hN`jW[I>Q\UWJ76nlEQ6e19jZ6lAkV6gFbG[@V_:UK9B`amdF53H3MJ;aXVliinp
dbhcJ8_X`UjmTcnJTDEb\hM2UcJ19]]fO<;]^_iAYEB_>CJhIl[m88lSC;_8RgVj
mN6UOg9gCe9@A5]WknF2YSHSD8V^g5qd]7;n399UnWHlNkA<eiO1agGL7AYl3^Sh
Y?SGbLXekPiD9B_^V^0[l`pG1KLg>T_`hKmHW`iIVPdZk8okPa?8M<4ETfBJ1\C2
\bJ6UDRW=DT^KU=OM_O7N^\OO`OFkek94@6i@bCi4=YCAbNg0bN7Ig;W;CAf1od]
Rcm<3KdP>gFF@:<kBp`TGOUXJFo<QAVh:9Q<c?A4hH>DSFUeaKenl=b?a4TPal]6
jK_em=GVmnEghT1K]Go@Ho0;nQ@ZjZk;b80Q@;i<2V5Da33DJB\L;]?VGP_ZaZBY
iiXc\@=m8lN0>dA=qT]A=21E:38]l<N:7KdQSkS>ND7h_aAGAf_TZO;Ybb?SnAB_
jl2j]in<W`N89J]\Lce2ChJN57S=`8ocCn_U2=X?W=\mFO=Vj>\<3X;ag@L>I@Fm
NlKbQ^jA?81qWBkkGD:h=A3H@O::TBG`9QXfaBo6DU<T34\A;8`IKoEnf=[_EnNW
Ql>>NW<56OJ4_6g:MZ@oAYTo6P_jbKJLW[0d]BpD0GXi:qJcb:=P_Y=fDoff>MHE
[pM1l;cf2E]5G4<A?KOl:mh\fT[O_\235PdUb2<_XC5V53N6G=Zi=]KjcYkEGGda
@Dh5[L_H@l1ablS;KJ2\bFabg@2fCq?=34YI^^^Wc`_;\MUAY31mh=[XD`Bk8J<K
ZF]JZ`cWfoT<R:QE<F>6SA3cI[na[hQBURCLI[Z>XM0OeF5T<NWFbc3`npN^P\iE
0$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA12(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
i80d;SQ:5DT^<e4a^?`J_le1lQ9Km<;RT2>>DB@fgQb[^<hh8@nBhjo4GBjFkop4
BVZ7E3d`V;k_3SoDN;ZEWAi0PB?``4:4TNf?anXR?=n@b`^A?2Mg1EhRUY=QQPlh
:fC7HKqg<=i7iZB?=@OI<2>86hSVec28R]UbiU6:BqT24V::pd[boZ5dgc=IM]^@
PI7[dPnWH9>51mBE<gdq1X`DXH?cX5NVil>M\?fT3`fj?9hC6Rh=8^qQc^WShA0m
B?ABE_\?MNI=IL>n7q6I7nN`:qh2L]`dqoAU==O1B8ULh;<nYl9gMC>_@j^V3EVi
b0ILIFB`R=A18;6@mgOFjnFNg1lJheKM@oTXhh?iCZl[JOd?3XkZD>38>ck_46c@
VCI?oY_b1Al0CZkb`2<\hSPphTS?^1L21Jao[JWYc@ZThJLQDK]DaTUc3ib5>8S]
INE:Vo1_RX<U=gEWUTEF4UiWh^HVMj[b3JnGZ=fLahL7Vo<k`GOhAHfJ7i=mjVHH
`8GQiDS8OIj9dmp4Wn\LRcB:h30R;c]EO^TnRKim3eNnF^kP^J:;@H=n9^[32_FM
YDZkBYnO^?qU;dB:RoeJKm@lF8ch_nfS?2=X@1j`moM>R\oVB1Se`IXIHlJDe99j
aZ<Oom9g]@NUOUI_J;@FM43A6PUo]b<8k9U@N_iXhe[bRL]iFTDj]k\c;4iSLgbE
GqRHLiQn04\6I=T=mIBdhIfLoY:=W]KhD48;d8E?E2?]W\_Ilh_GEP^AoXX]c8@>
5BRVEJe2d`;ESOn]U8iJhlY3p@5`Z2YqkFcd>a[ePP]C=KjH@EQTYI\APdfD]11@
lCQ7k9=e:2gl8>UdeioB=jgK^AmkAoJQk;GkMMEBm>c62QO?d0GqmZ\IlFX7W01I
oXmMmR4m@bAkk>^bELM\][kVWEO6E7XGR<SF;3\JjIBFcY>\HG:Tm_7fMSb2CGhj
@T_Sj@=p@N;NEB:$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA12P(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
0o2^4SQ:5DT^<EmH^;4JH49K[C1H_KL3PdYL][?mJ4X4Ol6H2:^1S0KI7m3=PchS
SBITiD0E_iI>p59cgnh2HalENkZ1>8nRbOWQV=T9B62X82Kk?FoWYMAbG@i5G>3`
9G8^cD8:oYgT6KRikAG5pPIIA5kN]MRT3KXoIH?EA;W<WJX6<82k1l71doTAZHA;
e4B6;ofTY=0HfHT98P>gO04aNpA]b`Y<qSKlPQ<=XFg:jPJjk^RbR2kV7P0>2Y6f
CbmqiHmd4?DVAcm_Sa>7SZQ3TnQ>?@:k2Fo=AJp1E5h5I=^S;EdRGk]XMf=2Ng10
9pMX5[F@2qhneM?kqfARR`mY_=FmP1@B4dLGTWK6cnK<YPfZT>k9g<Zej3R5Jhc7
:Zb1J[1LUGOW_2^]NfTDSF]C?M@l0Me0gQhhU20U;\h?4OP<JOkC6FEG>2L=Z<@4
L@m4EenpBHM4f27HFR>Pf=XS00SYc4<hEaj0;?a7;ncn\1@e\P1Ygc;=KJ7P57B0
DdWVL37aBi^YEE82mQ9I_I68^3Cl_K5E^9d`eiR6knS;k]]L]=d:LG82O4MHTapf
T\1@3f>JH>;JYED0m387`NZ]UcgA46pPP;F=P57Bll?\W2PE;0Tf^84I`fCe^Wo8
<fK95l_?925VWfGmE9g9DTiI7hcIjPOPcJP64bQ2WcTSHdDVjamm5T>8]nkVd0d\
<f\Sj2RC:h8]X94jCI\C8pfLMEP1T>h52nOJ\iUSD;@Xm<MWC5`;?l`G;3CT<D2C
1F`;;^_R[_d2Q`HO3Y^Yc[fXF8Qd_dj5:Me`o5:dS[@Kp>]CGjRpn2SA92?6WW6e
jMf9ee0b8[7aiVCdZTF^BCOQ:2aVj@KD^HmpdY;^:;\HkinXMBO_cnhCNO<E;U0o
Z>Q=C[FFkVh1m^@F]Mj3`2@QK??>dV<dD]IBdFJRmhk2T3879nE\@3apOZkWn?@=
[OM@9;RJL\]PnkP3b1Mm>J;gZbbaM7>nXI`INE3?heJ4ERACi35K>G=3OgTC5i;:
AgNF9X7iTH]q4ZNF2_Q$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA12S(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
ToUR7SQV5DT^<9Xl>R\\U7daB5J25=pJnIlA4a8b]j=8KC`7GL<HN:n`jako]m8h
f3iO9fFNBd9im;egT<LBHgpBh0_c63b[H18KY:01ZXEd<]fljLZcGbIkOa5hhfhD
0M\KZT[O5TXom?oK0@c:@X?E=aXbZqSJSFI?pbOf5Vn5fe2Z>IC=MGM2M1aU:NE@
[KKeU6<qXXI7FhWE[K4X7XYBe@k\ijBIX?I8Bgo;Y^p7hnd1i^GTUm]PiQjnElLg
b1o0Zqd[S7]6:q25A97Xq?L>_WASY3^GR[@6c^K]9NEnM5MA@Ie0DAHDY:bMkOHW
32>4UCU9b\?c:NVlDVemj?4<QkdWAK25PZ42\QI;bGV0go08N@Tf\[HGgK:FeaX:
1o4@AN]D2E=qo3B]0Bo7K]fO5<=YLF5_?UNNdO6\QMWBKI<b`GHfkg=W>nb]]Wn=
I<c\50aCS?c_ok6QW8Z_HQn91?ei>J@LOEdO4M\oW`PK>I5alE9aC>Z27FIF0M7=
W1p3NR3Q9Tj?4<CJnnB@Qk\]d\l<@kKcU=1`ZF3b\ngd1R[0R_>4J_Noj^ld]GVI
EH;36T9g6eK6;PbhIM2:gPmA`mfe086\`YnGZFfVlB2BD:gJSfOl`k^GTpg>U:Lm
UHXkPX`]m[e`eG^J2;=Il7ehmA>G6h?c6Q539G?U15W1R:SdRe[V1LBDbIR0Hdm>
qVA?nTeLYDN5DIOU0O=oHoM<6A?@F8R<9Di`iJHS>7kO`_n@GgPe_2=[bD>5X\Bf
aVe6>ZJmJi5AiZfdX2?h7h6p7h=M:Ep37MK15cQ\nWZ`no@;\oG050^KlFn>6:W]
Cn5bNMdUeC`ERh2Z[I`W3=2mh`Y5>1>3lbafnQYO7l?le_]1f:pR172MK6EaXN2A
WF:E2hO;O:D\hMdoRl[[OTl`f\=fM:WcHg1ema@GEXAgm=m\F2^R=W91]PcW3<2N
>Bn?[_pZIgoAl8U[WIiE`=^khPRkgWZpl>J^d__$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA12T(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
oe[j9SQd5DT^<XkYQanmi6TaTmEWiDJf[dJKIdP5B[ZqWfa[G;k^blKoLHb[q<]d
ol_ba1ifV[49G<G>^aL8mXAY3Ciaeqo7_GXMpG6A[N7D\:HG[cc6S6Ui`MQ8GAPF
dDcYcURp]:Q9F`;^U74NOM;HH@CT3_GX5Z`3cN><aOq@lMYYAf5AOl?B]:4^X13G
7dCa^p0>YP1U8p:S3WU7q1JLfEFm\fW?PK8h9@nFJL<?j=2>PeAIlM>ZH:;3JW8G
ZN2bW]OPcHO`?4VPBVHE31Rh=JZ8S2k`n2NUM^2k8^AY<k[]bi89X5>Zj7kN`X34
4KS5O1cTC\mp\:JT;JKB33Q\gVbVcI<PS=EYc3A6H>1e?M[gC:8O@Xi3b0KODM[N
1VUAQ1RNUOkD\Qh[HAJW\l;\e@VnReO7[Rk[[6^NO@WXfMB<m9WQRUObZbA\CD8k
3[pQWhcU\h1gNK=jBUnLc_g05gQbBcb>6dniUQ@B2plb7D4=oJ@LW3MTP5Rn3d:l
WmW?[EfY7iESUiB1]B3Y]_VIjNES[:eUOc;10A\^5alT;ajF3^G[H@SRF367jQ^5
oNJ^aQ<aFkGS?\keBX24fL9oN]5BDK;`pWLBXdM9F`A?0AS3K`<Y3D`n=W@\[;>\
[dfcWLT6ihF;k4SQFehZUFl`h68oXi]APW<93cFQSCbE8]UZiBVY_XXp=7\i_mq8
\hX4Ckj\c62kXO4[NPE4jgCh:?kX9T[km^d;O\Z]YR?fP;^f8Fj3:NGkI?o:b8h5
NZiBPb`i3Sb[lCAifaN59dp76VJTHMl=J::KdKoKjoYE:Gd:9>MWihN6d2n<ZLi8
_F1cQS[@Io0Mg20oW\B1P<<7?dU<EgQ>OfAAaPkXh6qZ>T=C=:aQ?`Ua^IW;fYIU
;Vp@nT;@Xj$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA13(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
7cLB]SQ:5DT^<NKR4DiQcT>FSk<4QOL0HcT71m5noI03^MG4We<f4[F=q^SUH8dU
OJEG`<NC;]=q5VJZfToO2iLFhJDKkCZ7]iJBh^iq7PjkAPq`8J3Mk\0oHPAEZ:^5
:2MbUk9SBg\80LO?jU8mejYp[`IedO23@WnG>]cJ97cHMRae9CggXe@R<?qU@Ri3
GgYK<9HVk[JiBO07DTAi<qU[EK:n[qL2RmmdTEm\J?Hi3@k<p`dSaU@pT^XMYoH5
XI[m[91`@G6m=5T3k_cQ27MG[bjDFaTH_0g_LcJW53_m[X\o6[9<7;U^T6`M_j;g
mVih6e`NTjDQMQTVBE?29SXbDbDDY\N=55KJL3\gPWW9dG_98CMN0V?Rf00X<BpF
E8M8efA[N=JV:Ee[Eh`V7m6W?6l^T\N8]UkO96;74\]1RdhC[k>mL9cVOWkO;10F
`m`KN0MSX>Q:G8X^Qo]Ah]JFTU6]4iCh]4MLiK;]MA=4`IRU5UNJcG`Q6o03_<9Z
ZdOG`p]NRe]Mo8gJ]>9IVY[kDZ>[ZOY3_;<F\2PK8c?[U0@Rhk=\HG3jj8iXaT@B
OWOLiE6=dgOJKqTfE:_dBL`:>RdbZhO>bfCIWBiWG5?lnS8^moH`Fd8KQI@<A21P
k\^lg_gIHa_6ETT<0J4hoHRYHOETC`VD0]RQ^P9[Rb?30?1^`oiF?Fk;AAGU97gk
TJQR`9]R5\?Li:]Ji`Y8qYWLG7Q^HkdL^J[WTYdbfQ60HDmC4Ikebg1@?R_C\a1K
:HZlZ:`6YS^SjEi1ZmTJnYAIXUnlW\Mbh<PZZniWN@E8@8NG4@jcbg1eEVbb>iEf
ff0S6Dm@=fHlQC[oG\P0XUEQ8m?p;mhD8;Jilnc;W9Zm:3VMIUTSc8G8]IfRn8=2
Ll]51^eo?TQ9K=hi;RZb?^]9bPXH;nWShM=1U^V1A1HnUIG7\bkc2>MPOk:6V8ZI
E1F:AoUYkiQP\jcg:<PcAG\AK23C:K9AWWq@R]62>\5oAMJ=^:TlE3W;F1OP5V6E
jUFXlf]fbYkUokj?84f<ahW]_:D@MY_1b:@@QF11R4?]8LbK;;cf:^BEUXHJ;ASN
f53[ldJnLhUPc:nW89Cbmk_L6h5107iN4\gd8gZEnpS_[T:e`fZ@CcXTVP>?ARI7
=:m1ad_M3GAAZ_e1f?28QLQ=U>\Gc]eN<n35OR>SLcSS^fNJn<Lh@JbGSO6C;hkX
>WEQ:?SINDdACjGZWSk=`f@`>g31:P912WZ`1>MWeYRD1Nd6pd9YASN6^m^5aG3<
nf:Ji_n9VFgmHI3cePVVbFbB6ZZJ;HfI0H7oJ9_Lld^C<FT]MdEBQ^2Ooi3oNo>l
:gbmXH?q3?^UKNpQWeK^M7=JGi[N;D1pgQRbeQ4K1hMbcbdcWUnB;_aEGhb8:ohB
EISEdmnC`[gE7X=iUKZ;U7PE8IhmRh:g[]2<iBe4OFBL7lTYco`:_93p6iJTRN9L
8e]YVcAFalmQnUPMlEDDhe1;1@UKj_O@><e>WHR=k=RK?LmQ5gRjfN@P12ahGHTT
a1Sl?^8P]XA^k\?q?`44U]F^Jol:Z034?E2`E;6Yf=WIgRjCk\UEn^aem>h>dPmN
K:Cc=O:AJObNCP>P?EYLPAA1B9SaKG3ARPQp6Q:Odeh$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA13P(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
UE\G2SQH5DT^<RbM_0b<Fkj2deJ]2_b2J<Wn_;7688WR:ISS4[UjNCCd8\4<XX6E
WfNEW3epN7]9i1gE29So4SRX^:5=@Mo]jbeDi8dTj[0iRGR1lMSkNaUa0eRYl^ql
Ddki=1n_9LRf<54L?N>=h03Va\NnEdlNc;a1SlqFQTC2Tp0_45HPZXmD82TU3[i7
9ZN_I^T6R73GY5c3EiJf`]qXSb5a7LJ=8eE9?e;W2<SCMfP7EU:L[DQ2Cq5@>H:l
;^ENS>N<O:i21ZoV0VXKlXYIY42S31fSA_ZLYSQU9i0nipFSG[NXLnoCMg]TZd9o
i4RF5CHlq>B1cM>8pL=f[F<q7ajG;4>8V7[Rg:\IZ:?GJ?M6He>0VBL9[IV=`]jU
ohm@l?5:TH9g\oG1:oHcd`k<7IQ=XXH\cScbETF6LZE4Q^@\j47RJOcd;I1><SfD
clQ:ZSR_hcQ?nmm5Z9P3Tgb7Y\;nCXp?4W[Y5MY^3hJB@]>A8c<<G4kHc;2h6L>O
\_NS1]Z4fPX26Rn<6dI4gdbK1C1minE?:PCa:>6MFO6KVHn]FGU@C_\bi9nZ_P^b
\S>=d16h[\58XG4_aCQ2Y?PX@P2]W[gd78\>lqS1f6\LDb2FPjS9JEi76Gbjg[SE
U<4ZV4hWCZ2D3@JB:Go9>BOV1^nW<?Z6jC?\i3SCgCcgS]b`nH6870a4SC`ReTL6
MVQo2>XWhZXmV:b?7XL\Hf:AY<LGTOmfNn@RXKb_ZYK=qmE>m<;D9gF>9VB21k6U
SDhXmJWeDkW0^PM[eJ\[nMalei[Ve9D;F0Z\q;UIGF:n:B@IH>VN>F23GUiTWJ7h
j1nhi7ZE0HQR4<8Oma19fEYbAL2`:k7`La8YW;WNj`J>R6]_eGdG?oMNC0TOl<79
jfW1NDZP1;9W9;5SXmJ;>]h^12WP\GmJ>3@BXklE94mp0Bd`naUG2a_?am?6M^Pk
6:clFREmIG\A>O7;OM6Jed42`hkM26GXaIfn>iL\jTCn07_ce<_OlZD]RbN>7`2N
OPUO0Ri_6PZm2O7;iHc4iC_]]O8@WTCTQiiC:j:AU\_I2DDY<Bp=cP6VX8ngU=a]
A>i8k]U[[fXdV\F<o`o5jGLZmRQlQ4jV]o]P[\K37=IQe;n\[PX=iWZURXo\m?gL
XACWPdZknUQCC?1o`jldjke[b<Y6\on>dFSHVmeZ@CIjO\ID]<hUnXP[`pTZ3gXJ
<Qgi\b2Cj0jcPKeg4`52?LSmUl3lZE<e;eck:e]m\`fK]VlICe;8]5e4?3T8eOSl
D`_V7MV2E@:CKRJHc39258leN5JlfI:IO@9N7:MZlMGXGRF8SlmoFek<_Xi5o;oc
p5`:l@dgDf;IC8Li0BkAX8[nRaU^7:Sn;BB0Qi5dGV0=^Wh3L9;WWLd[27[8XCoJ
05nX=cE\?3hSCgVE[WDESf2qORe7E6pEf:Weag@A4Ah4a`F2a9?MTLP6?ehaORnS
<A5E8MTb`^QIN3HABVJ87YWhmHdKYXQ[dM0c@9]JONn@O6WQfe;dG1pOFL7ifW=Y
9YXf_=b8OnO;kgJKG[8]lmB@ZmE\NPj[GLTVMTXPP3Y4d[]]Iim]PeW:fYn;WqTb
SJ3F4\OUF<Ac52SgEBYeX_V^>49d>ckJnG2B8EBD`e@J8]d@jm22fO\`nEGof_g\
L2NnZ]bU91=;NHEYN1IMKq9_?jdZh7>TTIc[Zj>1Vj^T4EAgA_[aRYZC>WH1F;gO
dDlTHON\CNmJDHlVI^D3m7HUK^JiZ?NfK3[2304]akJf7qFTN]kHZ$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA13S(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
5=fSnSQV5DT^<C3]L^OdYYe9qjS3BDEBP@]X9Xk@lPd83O8NqQA6aF8[e;71jZL=
Oa@I:0eJZVdn\01]DF6WDChYWj=13CV5IGog2NJE`[F4qIl?AG=ql\AWokj`aLI<
QCGBF89fE<]<?hfRUNOIY2c\\i\dqZ\DIB>=hj:8h>W;l4_K9>F[[]P9E\\h5d@p
JDlUG68B7BW5P>8hK11jB^o8R<qf88VI3RqMa6n4j4IY]3Nh_?[n]o9mEJPBZqC\
>3m8p^3J[kXjWnm^YYa9bT6YMnChAeKcG;b1;\d?V];ZMcY8NUALgS67MYdC5lC[
7aCKn^XCEI64B<bHgnT43VZAk^83DOhaXS`gH2d]Z_8hGB>hHFdUR[JcVicT@gL;
9`?4DNB5]?Cq\2@eVMKd8oFhR9ET7=OhUQ^iTDcEQ;leA1]_ACFC\m<EU:h4^G1=
n0HQ:l<?eKKn\U`VHU0o6\ik>JaGBkhLWjDG3=OjjdF0N1NXdl56AMB1Vc>;`K]i
S?<>e0Wg?d\j=lmdANpMo?g92_`7?OIm9Gj[8;P7WBaHGR5l>05YXIITS6[@]hQ9
RXejLJJKfCobgiYl?HMMJ^lXPLNH<5o;O=UZ8UIGPo@mCmZ>___8X^hH0KXS:B=W
jFhhK=`L\kblk99MnN\]SN;GYql6Nb:IEQam:bM\42_G]RbPQ6=]QS48VVB:0@o7
J[8[BBTFCGh7]XDV^iSN64N>3^l?jD`P9>0lBKEa?k^71G4j>1?[E]A2N@2:\Y1I
;H@RNIY\md7mA15N;@Ia9Y<>ehZW3D;6qYNiUcZQMeC7^boNgo6QICJ3U71?WE9Y
l?ciaTV5IZ9iV^:;mB\QKb7AKd_^>h[[PYhMRBk8[b?7L?4X\WSlnfhCP9ZKCh0j
XAc@FEl2d:8ZNf@kiVQY4WagNOROKfGXhMn?K4BpARKM8l60WQcZdAai18JCS;>3
:CIq^d?g>Kk=a[oDBP]>1ZS\=6kT]XPg=39PL^J6WVcM<5GU]N9f^Nae8hTbFRfK
?RW?^;UC_8[Pg9BAa9nUYHAm>8N3PUUgEXmHX^DMFWGQQW]K=m25;:;4DfUd6F?T
ea\YB^D;`CpDA6[hB]6gGfA?PGXTZkXN<6gjJ26MZ\HT`;bmDR1KBk0fFDKjNO\`
dM`ic3WonR8D?a<`2Bc_VRogV?`mm1SQTGVT^[G9RN6G`BA4RRS:A0iO8Y=?Ia>H
D27kZ`m8;cj>bCI[_p?oFI\nWAg1b^h\=_dAoDc9TfYFI4X0mS]m>RYnVeC>EiI@
CgdBDFj[EMdA6543[M?X9Wl1DGYhVBhLAaTOA\PYpokanASp<US<dV?`28mRQ<9;
UMZB>oW<l_AmUMAmmJl`WaFbo4KM=PB6YeM_Klk9=5?emGR9Al=`Nk;4FLiZHZcF
@I@?5e;poN3]86iQ_G<h<G2`?4mdC8g85L;bZbBmfUY=_^@0g_@6Y5J>0B;`[@\l
gI<=AdjC>l0<TdAl?`2eG[6\a5jbX<Gqh?3eQKYhbKTH\h=QYPYO[B^WSI^D=Li9
HMV=mgB2BlmRd>M;j3e=[WahAc]IM5JIh3[5L`DPa_WTK\jXgYbpVNGb0lHoi>D:
dSeqP[^o2:H$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA13T(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
bcUhkSQd5DT^<LC`4n1Fgi^iMLW_NVje3F3AKPq7DKm8L;?QBH1@PJ7CbW7keA9X
LNei=TCq6KjOU<jRNK6MF6><m2f78WXoo]4ZXXW?B^KP1J1Lgb5Mn2;QP\kbZk_D
;151b\QK>:O@W298qM[PTj`q;\gfHB3?]XSed<O:F7d`J6k_0dA4ZURXe4AU^NIb
q^@6h7QNjC:51knaRS?<gb1fL;dEJFP`@>Bq01n]:<_eY;=cKHVSVa`W`?f7lYpk
:O4Zckq\SR^7XqU063?\CSBUh1UR2=3?NVXolNPNQ>m0QikXa9j?qX`=dkMR^[HD
6]oBIdO:nRi2C\0:=V2<W8>klnZcaRYC6`]IUA<7D6h1N7NTiIhb\<HV0W9J?]oU
\l3cG>bEDKBmlY2?PCHW[PS8MbZCZcoV`Hi7mm9ibo^jY=[ilejT`miWi=lJ66Xq
KQ0L[l^PNEKGMOmIK>[6:ng5Z;j\^l5\boj6eObe1`P[L2=oJ00DMBE^RH9TXFB5
laR?9bLNI0GG[XI2E438P8=]^j2?SL36Q[ZeFO_g?NRYASJe@RfTd3LhK\8HiR@H
:5e9_Yj3@BpbaQPgo^WbLkF8ViDCM04HUbB\d2O3:m\ZO>`XQKL`bN=U57;]VUcK
TF=TV0HmKTl@M6cRF3R0lWfKV@3_dADInIT7e<To115CT@ElQoZ\7?6XUj3<BaNF
eOd2c=Z6]1ZZ9=IYGA_Hgq:0IkQ\SBK?a5`Kg6?9\7gJS0HkRKWUiYo^WJT9XXna
77]W^:f8[56_b^D[1_XaW1fGN@[@obNn7DR_9E[Y5k6iceQai`X:bY0WKi;9VWZf
C@\SmH4H2b\d[P>]ceLh\abY:3D][9ZcqiY6Fib\W<_FP_n9VPdmP6?6>DV0V;bQ
8X0FfbdblOIP8EifLBRZTN1gUeMSbcNCU:mX=7GUoOb9JI7BFj:W@8i4MQA:^7E^
T2cP]kd2Y?cPZBSha]Pm@D93=9b5dUf\;8E\O^JML8CqJ1RS3QNh=d[e3R;0VS@Q
=8ol9EJ<I:DkE52YRaBZi>]=[]cE0`chkA3iUnD\:oX:>?Q<fak:804e@<nHK0>3
@K2l=i@PEU^kRWboIaQGf:fMi5hlB0VonnYW`lfl1MolSNk^9n_U\dqWoi]jfa7D
Y<:UF?Dp^7:>fVOlTk7Cf9VR@l:QTPi2oj8]V`JRNfdBKI\]]fgZW8=P9:UgGaKO
CcjK<N7A]\kRE9gNbkF4ohihk[khmnUNZS1W4QV5hS]ThIKMN^l>a]R>7Z@7VG6U
494ooo1dFIAD^=CP1GpB3DC^5^ZZRZi:dgkab\eR=A3BdFIK[bXNDgF[hYk7Kg]9
W@<S@9EKbSkb3VGI>0[4^TQdKU>=D@]TDBBPO<DDJX[3GqXa^1`WqVFl9`c]HRCd
Q`b@MJ6]B\o7263iN@YndM]a8e]7k6\O<BT\o28H<dfX>W5[?[fV30CLOWJdT=:h
MQe<;PH5b2Va`oMUqAnZNO6cP[WUP6HbRPMpUlg5CLk8SBAe2VW8h_W]M5?3>6JI
1]mV_MT29Qk:i7Y`<o[4OZQ]VJ011AGeQ=2kMPXH6YZS30>J5MTG7:ACdXnq_L69
OTQlF[`KX_Dl_WbX31b5A=]Vk>glQT1WHFcLeIg]El;Y8KYGIFhMC_7j_If6U5FK
g3W71A78DLY9W@Ng2D@pk]m[hS:$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA22(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
BEfJ>SQH5DT^<>:lTQ_O1OFD2OjCoa1nRh8<0<1oY3Bk>YV;Fh6q8DE_JcSF];IJ
40]YH^dmh]_GPHWhLDjN@i<134kURjO:qIcl36BdX_RW\c5C?:AH180\jDPL\`IN
^?68kC\gRVnnQ;@H@:^Q>@5=LpKF_BFbq=eXijL0j?>?G00I@1\<Z6amhL`^^?lK
^@0plffQ92[@gY@DcZI=CL]39nPjN9K\4S_]QWpZ0ehQCA\G]\WGgB4LWC5NGLoJ
[^[ZgQM81p7J?>>MNmaXeb`0Y7o>Gg6_ITI1p7?`3ef_p^_:ohZpHOa2ieULE<;0
h:1bif7<H1bD0PVM_?@2;i3beFH^V1MB1E^`f>DBaJ?d1Jb^6FO^HXKnonWYB5XL
c\XX>ghdM1^nPglVP05`Zij;4CM[WFiW53di>B4i`7p>2VDJBbZD:G1gM[[SEfjl
SH=b@NI=???LKiOF4bpV9<edN5D;NoR^PM[B4@7Q\aoMVQ@0c6P^9f4BDCEP9<=X
U]Ko`b_VVIbmH>R<eNBVSK[K1JInIGV]L]TJndC3`S:_:hH;0oS[9=YS[E`@[_J8
kcd2lFA[>pdOJ1KHNM]So7lg>k8JTmR055RE`39X9;e:[Q^Q^c:]l8IO9jaOSe\U
:9dhMMkLDXdZT4nl1n:^?2\Hm3gj5OcKQEL<l1^Uc5::>58JU@jdE1V\cQb4V:bI
q2H@N2I:[7MO_3FPgC@G8QNMD[R1U6dmEGeZ;X0EiifEOKgQ[JYk:k`KN9]\In=[
Q254V\?PZ?QjYF8=k35S@VNpAD54QnMoUoU[^g2@`Dj5C[2WlQP?C>U8KKP:l4be
i@dMlV0Hc8lXEUjP;JmML[2RA35:W36dZ_6TjMZRh\GfEFgjnSfH4iSXGKS\_mE@
66m]ioBS:E1K7bpY2F>UK\<LYGbNW\D_fVVm:7cFg^He9e8OSQ5?l=EcnfqhRXkC
DFiJ@RVJIS9V<SBm2oONNFVJ:kY0ROY98_e2Ia7K7e5:jm3H1oojih<^<9_h1L\Z
g7N3mC];AfV`k4YP9`U2NoAk9L3kROYdCBDlH\H<b\Q]QQodOq8_1^jAK5>KRj^i
M^1<TXGB;G4eo7d@EI34]V7O=I8iGLlNC=[<N;fI1]@FjlICaV8V0O3m>TG3\I?V
L@@o<8aTi9S^=LQbmn^40lWTTojJC6HCSBc81H[hq04W;:cJ8h>\H[PHB8bLLeSh
kbVQB?m3MOoR0]Ch[c_IlAH:[hK]TQWNH2f]54b6l0BUiEL7^>HicDK9lT0UbKPp
\b@59nNo1VAXInC>0ahjCOja^hM<Bbfca_DU5]b6dHC5oMm\qD=7AhS`8XT49Y=i
HWbY0Ck6VVYW2HCjcPoI?J]HU[Ye]a_TcEaFTd1hJJ_FT[>W\;dkHDdiVoEa7:Ek
ELd>54YQngngaL`C@>[No6]^bAAY:7B0Hf5^0DGjja>q_B^\_aHQ`_Fdf=Y>SR8@
9RCDM194=0T\]B\bkJd?2<JL@:6<?J79[\AEPZ5nbZH<B:<X;Rah?3j8:fNc>W==
JI0cRcj1LG`^Q`X=fJ8iN:4iS9FbfW:mkLhTeYqAESdB5afW4B\JADeF=ge3T7HW
\:<nYUc=^>CG7;?QI@Cd\9:P^gkl21GVKV5]0Ln\^aW7SmSMC1332lI1nSZIFj:T
HfCU]fTBok5]7;eNe6Z<f78Pnl<Z_DSmcp3oGoUG>80jS>c73T4oiEB0GQW1JI\1
VLEOX[1GXBkejiBXTEJTRXgnclFnk_]ZU<^IZY`GAGOKg>NYTQ4dAkgLb=H7qb1`
US5EY?gTUB[dif1F;pjXID_ccMbDn6NTPik@m6G2:Qe1:ZeKdZ7FW\bO`IXQUQ9@
ITPgTad`g?j6P9fgnP\N96:0Y@gB7i>=?GloEd>\6oIn0WY:7a=`A73O:S?V=jCk
k@bX4[TiJjbLp_7ke[\5kTABW;A^[fbH[;G4\AL\OYS\g]<1iTE<B=E2>KmWReaV
`5nEQa`A7k=gC35`KTMDn<\j2LiJK\\c:M>adk99lYm?PLI^bUEPhW@?A\gYN=af
ONo:YK7p6<^ADNJM>9B3PNm>DMi_b\>UZXU:KLN6^8SALRhmVI88Tlf_X<CcCmdR
DZ?;TTGinRm`TRkKTGImNZMEIo1N@E@b=RGh:e6:5N7QaR5JD2W[P6J[_mAAE6XZ
kapU\4JE@^AP<HRh[gH?\SlE4g[oMUHB5Tm4d`d<4CeJ>>>]ObGmgOCAMiU^C^bE
3f8^LY:96g]mUXmKdnL_LRX5]EIWQpKN<>nlR1C730MLCQY<@_Md:;XV^cn0WWDR
qI3k?GWqJmIgj:b$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA222(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
>[aF`SQd5DT^<N;:U@hkcC<\YNRC;YKfaBS1o2Z=b^>kY7l@QBD7VBikRbMB7QED
pDd\\P=5oLGLmG<LZ`mj6nT9Oa_a]SLL6WUG86fnp?lK@ecPd23hYL2gYDOaca:g
0aKQ>YilKPWdZ0CJf1P7bT?@X?=Y46D4J=5i`L@Pp;6d18Lq60bRhmj:NL5kJW5B
BRgIR6RNZZ]8S@nhg8p=cP6`F\R\k:29UAOYAV<lUn<8hMl]`i=aBqcY0DJNWIJ`
4i?LYUGahdhLCaiP7Hd?1J54p4=cO=d:0G?3B_gD]R3ckmEgN>PBVPfo5JOZW@gI
WqLj7aYkl3me0[M@\H`<2[=<jVSJq;`elAn0q02QiR\AQ`?EIkFN4MDS=0cXW;KL
II45dE^d1^39j2ZXnbRQcHPpkNF_]_plDNV0>LBkGhI`O?B<ha@:7Wd`8OPOJ;jS
Nl0OW0BjK^:[W^iIhCZlWIQX9[[HVIilYc^cb``X414L8SkBGgN^TWFnO:i5:Wi8
Nk_C>7QLi;ZZmY0bO;LIG_:C41G=V3FljF`Nb11XEDDL8SkMCQe\Sq72Sdb9T76@
hBm6mg;eSbiXQ?Yc^DPEi;G3NjbPZ4]I1dbhMe\NKW8?5L[[=Y6c3IV`WXi5B4N=
=KA<]a:^mVP9A;:1Nakf0:Ln22G3OH@]>G^8:cl4SO2TnFF04Ml@GLn`i=iJ_ii=
XmAPYk:^mV\>jQ>ep3AfNTOIgBE\aoc5UiCo9>:0E`NMgQdUnjd_GXGj027[?naB
2:D8C>PC1M3\9O_XX34YlX?FP2B`ZemKa21li7aRVo`NaUTT_ld01b>:?N`<W^P=
cg[c1`5agcL8_f_Xl3[?F0?Ic2]mJemKa<4?j=5q3cEXLGFAS=0I;G=AiT>>G6aP
O]LIGQZOU4jU]a<969CW8[YK\cW`mA]n@\?NA;YK3I8<O\]6W7VfR8`]KmTkb51^
baH=JTV7i4^4LNgEEclJ[>_3]m>ic?_]BcbeT;4F3VVJH\IRW4WOR8`]kl<Nbkq_
foS:KjZRQalZ<]Z@LfhV;M=^H;T@W\@66Z7H5\[<3LYEVE;KeY3b\^DNkm_n375?
hLOB1EmBj>FMKX4JCDBF5U3SMYQ33eTcm\[kM\[87QiRVn8BA81m3o2:?BE==i_G
hXWBC3^fj3RMV=RJCDB9G>7:BqWB2eMJJOC1G07=KbD21;06WSODcd;hQBl<FFUM
TQd0Xmb5M^\8P0JU]?M?\dnGj?WAVK_oXH>hMI4OK;Xj^4cHh6@NBeKaISl<2g4h
k0PWk?NMN?VefE\nJgm^K=CG0gWPbKOo66>_C34OK;1[oL;>q0Ukcl][VH0FGCEk
[@7Hk9`Cd0^_iXClS8NG4D0a>VeBVZ8<Y`]Y:>>TKGMlD`^;=0g2Ve5A39hMFUlY
\\8AeEM083N]`;PglgN=F4H6XeR@eI^9VBV<6?[f0k`OiB^m^0LAn55dE97J3UlY
\>9[Y<2q<OQF<\V>3TWg`RN]5ZHbMif7Lmmo[Fa2OB0_AV57ediOOU5CfM0IE\jV
Ta^bCgY6J>9:<0Tf<`TlFQ4ln@<KSO?:GQCoCX85Z4U9KK5YK1ec3^b8dVmakm=U
2U5?CoobV>::<[H_F`L=FCein@<KL<`AjBp3YbVd@knV>H9Z6PQMCfdSfQ<QhYm`
1m=HWlk<j2_Dla[EgYpUCj8=V@XeejLISVlHbHWFQ@?3i<UYWA2ZanD_WoJL2P=Q
DgR>hXm\FQ9<EAP2BE6USijDO@[KKi_1?iO`\7@J<Sh41^m3FIa]aQC@lm0FjFoc
Ym<551OScXfNQfcmB_`UM9@2O^MK5RT1?iO`A7BVCq6K]c_2DYkC9[D@45h3c]P4
0\M60DoToA\CkJf`1OY;H\:KMn2ZUB0UjR7<B<k1M@6Ydc]I>\h5G1lCnQ^NC`Pa
qYGNh3]_8LkD@Y2G5ADS3PJIja_j3kC6^:CL6IOH?>SV_Y8clQnVk_SKH6ofFcOe
@4nV50a5V=Lh7KAOGR@@O?db1BS;kbd@T1Oa>jO3B7Re6AOGAg;[=j;F1f3Ab1=n
EWn5g0_=NLLNKKADmR@@OOM4>RlqGA5:kJ3Ld6GF7=b`eU5eP`L\D[8V:6:lSP`c
D^W]Z4dH[n?16[H_e;\kNCF=aW0;[g8dQQdWKG?HTMYZWS[2g2Hfm7a042JLj7AZ
^^k[1janBYVD[TDd:mQ:N3C0:ACIYgHdQOm@\G]<TMaKWS[20FLP>cqOWecMenH:
jmY9dUH[DDV\onWcDogUS3=MLQWMH<R?eeca;iC5[3c\MFN8a;G;kCRmFEDHh=0k
=@QZTWeIh3V03=EADonH6C4Ecmd0Z2PThHJU<ol9?CZ]e1hVkRVc`:SO=`Heh0bk
cHLUT@XIhHF03=E=lK?RSqa`E_3]<JU6E1j=M[2g0M?oGY:V]S?Q;h;Zd6S_<>cK
7CWaAKL:[Ckcb]`GeR;=L^Vk1>@^2Y=M<M>@JF`@c]o\:UTW8Ei@RG@Q4>8_G\JX
;?VT1;P>[^E:B6i9\27GJ=>k2a@]N32M]N>@^_`@c]XXBb@BqhKJAc83894eT4m:
Do9m:HBVCc001;;e[WX2j3oIVomCFKLco0W@Y5`2oEPSfUmqPD@`Q92@:<b_:12m
3Kg_:n=hMYd6Y^U`h_OY81i3L<;?A`Eb9<hG[NiYK:J`H<Wo?T<1?ScanY668]BZ
lHoV2cYDlY[;6Z[@`\Qcl5BcOSm8=X7biYj8_dgj\NMC7^cfP6Mc<SXKn;6mK]XW
lH2V2cYDhOLinmqOdl2<;cW@BbU3HZddDCUcbl<fZVFj?ofnOc6cJ;T8<BOY=U8P
@<a=in?l3IJdGUVWJ[ia5^^M3AKZn1GTG`PQ;[>Mi2[lh95f;3[LJ\F6X207L6SV
5HOPfea6df=Yj]0kJ5oa3\fe3oVZngGTG`P;n5QfRp_6MBdXB?3fEi4^6WSOM[1l
L:;]5B2VYkajNm9ah1k_o;kifHC53JFA110D4d=F:[VIo;QTkNVmme1F0LoaZEKC
;;`]f8ON[97LW5_?T_ZfPghD50`XB8@o5Q5nGKhJG4_G3g[Ti]V1\gVFZ7oaoMKC
;;0aU0j8pU0dMTgmH?K4P]R649mF30\1Z\]1mfRUO5AN93D?a?^C0kXnC8OmQL[W
>aZEUB7dV>Th3oE7[gfBne16jUK6XZj0QJ]TXbJIf2Wg>5]jBMU6?igfgbOh<>:f
abK]P?jJAUjTI<Em^gM4Go176UK]UZj0Q4hYBG:q<akNSN6OJ`fVVZC>K<IZ46eb
GoDK>V]cV@d?ckXj;S`WcR<9FXTY:Y_L7T>9X8V<KIj=]J`H[Y9:71Nmk:aDXKMB
Iolcj[JJb2i1^P<L`V`8Ii0I]6O@e6f:@L9cmeGH<el^PJ^L[<f^C1Nkk:>dXKMB
h:cQo<pA95HF@3\@g_IT\_5b2Hl50UKS0K?oA\`9l=aTAjEH9M[aUJ5^knCR:okC
aT50RQ?e=57Y@oXQO77<dG3GXiNn6BoV4TL1PqEAGHleXk3C7[mn=O4Y;>?PWod\
XSZkn\[b^R]JeLBJh^DeF]TU]O=6CYMhYWU5G@9b>A3`_56ZEKB1A>LnPUcNGRB\
L33[I<`GdcSG3Al7h9?@SYKW`n6hT>We]oKlF\E\hl<`ma6h7<T1=:LEVUcNGR=O
lLFep=HPCKYW^\oE=if?eW2[2Y=f]S3Mmon3Jn]Xli0Gc^Y_kn@5KPi1TS8^g90R
U]3e174`S^A\jkfS?IREP495\F?`4O3UPC[4bFCR0_H;>:1:9jPmX1leoXM<AfiM
o0B=;=F[JOA65k^RhgRQ944R1F?`4^DS1`cqMZXJQgLie=cRGj7@5jGT>SR5MlWo
hFb>P8J\jJni;eWV?c:K3Tb<XCFgJ>af[3QM5FHFZn6p1?ccmk?;3I8M>LcQRXUf
_2bh60?NakWEB1mO?WDe=@A8FhPPlf?ZUj3Lfk8Gk\YhWS:=<08cd2_3dn^e>cML
G8ee`0;ejQ1M[_3b4YN3nUU3L1\c\7YFb9G^A^d8\?:61I5hd0:cde88DnbY>=B2
G8eeCEZ\?1q`J^]W;eNC2@6OiOnE@K<cHlnNE]0?FFZFdg4W[mg`?GFTJebnhI_Q
]GXTZ<_JUR1BS=9dG4a0iPZa>E1R?0oC_Wm@EFagZmLW9JCl3D@VPTI>]mag<DeZ
1O5[[_[`a:l`<g^HG?70dJNC>4OR@k?C_WmCinLITqFPhMC;3ngUGG7S4T=EEB2Z
7fn_=Po0NVgJ\iocg?k>i<8VRISmQY_B0Mhe4nL[]]7XZF?a]:c4i5f]UVYVg<0F
\4h_=P_bG^SWcP:6E>Fki@[Xf:3mOJZUoSA<A]8`MJF]<62a^fccG_i]=@YVXg0F
\45DW>[=q[=m]>;7Z[P@2YBC2=QCKdUV\AD<1cOP=JLG=V5E3X^`jC4Nj=d\6XFO
7eiVDmeUJkZYJZcRLWLf9mgDGmBH4Q^I_KD^1B8PRmmZbNShj\l<cb]E4m:392a?
5WYN\;jGi[]nflc8`WH@\SgZQmFiSQ^I_fZ41N2qV8eU@mcDCIMB:Z7=FcWV>Gdb
FA1KK9JD;;Y\b1M@fl:nAE>ZKXh4ib3VjG@X?=\U\3H;2?NUUC91@jY7jYm7l[\8
aTK[GnK4?UH[M1f:n8W]eC]_n]9E]lKZg[UiTWLM?3dB2k`O^CkS@EWJjYm742kA
n<qW9fXm<S4ONR]?Al6cc=P^9li:3DiIh[P[ki9H;RjJ9E][gN;]lS<TSjl5iI08
Re6LIRRdc573[3]EUGI[WGmiUI]_3DiQm<Nno=GGge0?`EkIWJ^>@GR2>HgNnglY
]D=W1YdPcV73ZR]gUiE[g^XiUI]BXIL<6q[YIcD;;;b8A]b;>2laYiMh7HNXmP[F
LK7\TmbFbG]9g^Z\KG>`nlaMhiX26?Fj4B`ei=:_24N=HC3aDlka:kVAcdGXd4dR
3O_5?O[daDlnG?Ymd\=D7lP:<f?OHfHbQf[O:F]_ZaNM]KmaKik9PJVAcd<Z=0C2
pUMU7c3RH6eKF1Q_EQ??CP7CMRjm>3@_;K<Ya=3RobhGiOHRCn[4iNLnfl]1K_EJ
@fGm1=<0=4<4P:I5YM?ahX09j_gcoj>qg]Uj;]4`6HB0[\ADLcJn7EIlT=3Ihd[4
A1klJJQ\:ojn9DQT[e?m59IeC6cIEf9hcUN:?c?SM>3BR4j]edX<TPT>7VEJ]6`B
bA;I5JLQ[\n<:^bO3A[Lkc:29;BSR^hIPU\:?`@U<>16R4jSedX<6ejT02qkP_bW
`P?[c73a^n:d\T?o_c?`L`>:KXDleL7HNABCZc7JCSA4Z2ObX=q\K]]7bSNQNC:6
KQlj33Ym19eRJZhW[n\``h@;cln0MQ3jV[`kLn7B4\ndYi=m?BXeX>leVfP_<>n7
YNPXcHS=m8lXJU]Xk20`of]f;8R@BQdS;Td0Qbki4bKBDaL3DJB\La]?VGP_ZaZB
YiiXc?2=m8lN0K]OHqHmSBH^:<1V[=YLMVN6kdPRmA^UTl;MMTR;IT\SfFSXCLe4
L3mm=>HkEK=>4KPT:\CC?KRTQ^e=\oV1l89ZC7iCYagUElOClJm_j=mbPE6Dk88L
<NLXDbL=<C>_7_lXe0H]Zi:T5>eH[3X1[89Z=2iCYai0QBZlqc=K8CEKFQ0?<PNK
>K5Ec3@1eC@@;dEb;D\PZ?8YF;L_g:O3AWXM5A3KKbF`[WIeP6@hM9[cTHW:>82L
aaIX78OEnghQ[H7S=7K:A<8dGI9Zd`]@IJglTjQT[5Q\\\MdF9@?:9een=W2E82S
aaIX7gBd_OWq0XC8:d>I3W88[4FFgkf4DEeqdbIPo<N`;1\3nX=\QUH1bebc_1<b
9bBWbW1WDXgVaM;\eQ[`<EW6n0Wg7VH^Z5mjVDeag[YE64ADNX`?0O422``V>1b_
JX<R9\0nici:?jhUHb@NRHmdNNBX]8N`gDGmdImcH[9<6B\_QXN20OL92``VLjBj
`DpGGJJ2ek8a9C1[8F>g\Bf>Mo3K]H>:GMg2[I4`dmbb\3I7lYeo13V`nFbAOG8B
\1lZ<L7;g=ncA0NmKlThnh;d]FF7]H>_W:o@ofYjGQ2WlTTm2ajg14RYB_QO[o5Z
PJdGh9>mgi6cfC7QK<lhnind]FF8Emm2lpUn`Pa2eY5X[V5Ti6=nWZjiM8TiAb4U
;X\:X4N8:SPjab[ldB[KId^gda^Ni5b<M[kC4H3nLc1bEd]T8:E9j[Z[Uagonj][
Vm7eR4<8KMVWC=2SJEEl>`0GlG_^XN7WkMMC7V3M4I:bEH]TGBE9j[a;_EH0qj;=
4k0ZcRL0IbgGj6:06gMaDZFS7hTC4TXD1JF2\\PMO1bm^eEL8DXYP;CHEfGm1:nX
_\]K<1nIHmelUhQB`RMGQ8F3NoeeY8IROK\hF]?b8h=7<F3Rk=DC`gA`MDD1YjC1
B`]Uc1P0:[e@bhQ:cRMGQjj:07VpchE>HQ6BSO69JWPkjjeR9<o\c06<N3KWYO7o
;hfHOb:VN[Sd;a;:@]H@mUY5dh:cClQVgZjoM7gdRd>1XeC?:TDZ<06T0?Y4hXe_
V`aP\A:>G@JA8O]i_doogi_WE350c`iU0Z<HM29a1doeXe>Z:TDZ`eVbR4q>CW8m
]I^AM]?F?`2A5^8Y\YT<MAR_nS[=OAhVZBm9dnZd:nJ]4c[F<2KidoOmZK>n=hO3
31fcMbo6conCoY=`[1ZNn=cgnq:edShR4K9biQdg6[L@cIj[QP`6kVXU>c`UXj9n
8VdeLGXdTBkllq91V33KC2Pf6COUaCeQlaFm5g0kImEHJ_`XmQO0iBFA>@bo9WeR
T\6T4d<`2o9S?`\C21[7fOm>Y3nmm:4B@fO4^dEkIA3>e7H>kTV4Xf\bFbHA;J1R
JZ4KNd1=h:GMHI9KE4M7RgmXjJ2mDY4Q3IO4^dn@JObCpl7iBCmkA@`QAXX94K?C
<W`81;?Ed:3_NZX44B1;J0ZdFmgZEmJ4eGd37dHo64AiNdacH]6eo=]M9?PO]nFN
J6`5G[?];JF^`GF=h>fM?[65TVaoA@>Y2a8^NGL60A^U:ldiNB6Q]=8Q_@PB4n7P
16`5G1G4EM:qLS[L>aBUa3=jWSm[I;<Kk2^lB@9294kJn@>bU:fG[Fl<h]ebBOkV
AQW\UD;;ZOVCYfXkG\A<m]g=CmF@PFjB_TPRg@h=TSR4>KbG555LcQiPN8Igh:WR
Z80WT>k>9ANKL7`\>\7YmU]comI?PLd0_TPRWh3URhp>jE16W`m8Uh9ZI]TZk:4h
cI1NABFa2JnjIkclZ=MW`qSE\8AGllAL7A2B_4DiTcFIW1:i0_RP\2S3CN_3ERaF
P6n`NFjg>PJC4k?ALKL94KHR9O:>Dj5fGWKRge8iG@8T65\i2fiOciAY=IiL[`\f
O``G<Tm^KNMS_2CLic35jLSk\:Z>Z35c79]R\_8nJa8T65nFjOL0qLa320nfBR9a
Q9]bB^mgmaNR<aE<kNEE9f;bZdF_W6@a;Rhmm1hd90@QU[aoHT:mL8PSgHWWaOL3
U4L^hi_VKkJV019<VIifX1P1e<FY0Hojo[^kd1SNG_XRKYl<iOCSc?P^gHRi2hLZ
44W:5i_VK\I]E41p<LN:\Mf]ja`oH:7M:0E4l61S3Y4mi\X2;nQ3B>cFo;7:nBJQ
Jm=c[OfWFQcSQ3KLk`KcTNgg>X[^AfnMnkkjiRPWTYe=UWLeC=QXk=jdF5<n@onS
4TY`a9?0:f=n<0jk<5_RmNi0>>`m>f5Vn=40iRPW9Ph\i^qZ;XQC>5jJ]IRS<2gC
9gNl;R5EO<n@:Uc7QF8GJqd[bFIFa1X]9h8GCmRceX3D=?7k9CL;dG5AP8_=3M<R
^;f\FR^M@C3P5UH[RS0B?GVbJBD@eeU_94g7WlOB8>^h7mfk90`imC_2_9And8o9
M=MHEMk>F\e`g`4IJNmceedK9JQ@H`UH90n7CKOcnY^h7mOZCG1Bq44=Y]coD1U^
alTUL:@ERkDV^BAP8X^@h99\[og7WbLGMUJFLjddj\^nBKT\:BE]@VF\EZ[E;Q6]
In6gGiB99KnHOgh@XWWLdeEdGjg7n6EZ5c`mUQO3251M8AWN0^`15_Fo1Z;[436Q
nn]<GiB99Vk0l7]q0\IRB;IBh=73PdDKQI=DmSZAOmO?1nA7N7ci=QV_l:eLNVCe
TkdD1`bHk6MmT8da2S32mQb:Em6F7S<\l=naVHW_\m=`=BOVYk7NkoYAY_eo2kHA
iDRVNh:CI0Mn5B520g>9hQLiEN7RJSYYlOB5VHW_VU^OC5qKF5F]CT<;k3842UJ4
YClpfP_08\eREfQ2`fn];ha>C^NUeJN2I5C3P70AMlJAj7Hi[VH>M]IEk>TRmH`a
>A:>M?CeoTBW^FC8je8ZL@2=Oe8;7OhZ_WpcQ3>4oD_@Ag^5<V`n[66V_M[7:9Y0
OE:1a<iLnmAT@[68mb0A0nim4ReID=5lB3o@\G[AW_AH4L[E<CkNZA^3g^dN:OYX
8]:H]j7B5f5_34?EPJ>WOafhl^hm5\TnMFGcT9[jW6fH^g^C<]]NZ^N3g^d65NOg
Dp4ff`lnIE@3h=eUfR=5J_hQVo=49J^450DTCjZVkKMR3C958<WQ54;oM[Wn?\3o
<^SENUgJ0=g[;I[k=ggeF1\C?[;4Sgjf91gHBHaliA8HX^_4Mk==bm^XZAbhXLdf
KU4FAO0JOmgkhf8k8Lge70\C?[3E3B_Cq_Oe[j>JEBn6>n63VCXC72RCT09cB[kZ
=X2=UM\`EP7^j2YV4NgOP20jL_P68Qh>9C7BB\P9TXBUoLmFBPhaUN`T1?9HAW4@
kBFNPLC0KV94Fg::XM3lA9NPhl4T2aGEX_[YfgP2AXo6S3mQEPh_cN`T1B?EUDip
gFC6:Kj[O\mOL`UgGXkJ8`WilZ2oN2`cjMjnmkFESF\n2SLY5IbK@8b[A@69dWEV
dNe?gmR9YPKOZU_Fb1`TgXJoFZd\oa^bIJ\bgYCB`SAhj7fG3??SEHCoZd=jbKPY
g444jmekY^`gOU[kb1ERgXJoP3iEQaqS5FNd9Rb@<gT6FHHgL]91Z:nE\ZQZAR70
SECf617;LVg12JB3=kajW^2VO^n^=2XGGMG<dB7SW_mcob]88:iK^10I\50d>ilI
aUo`LVPJ9V=mHQ1`IL97_L^0Y]fe8:cS_AjDdgjSfgiFoG:889gK^1097`Bg^qAZ
JJaf@i8TLI2X@?A;CH[Q:]GYF345Ed]3e<\hODbGi6]bVCCE[AS1LQiMlVO`FaR3
kQ[[LWZ@>mb\@JkUTV4D@gCYKn`m;?[Q3?2_^[UW;JhY<\HY7HUgWC19Ti`kRgAF
Z<T[gjZXL[T\nLkUS[4D@g<dLEJGq90mT=EiiKmllGK@diH4OG9mbm;na[Za\@e`
l_7BTUbBekI;=fgOUn6PDnZ7Ce0S`g[p\Q6a;Q_X<mFhVKOJ@^FS\V6Lb9RQ4GZH
2T\OmGBSTADD8bQ;_G?GSmLBg8g]?mi;cOFD8d9`@Y>ohPBCJc;=F;YCCDMg4^?l
T3TYKG`>^CP0@W_K84l29R8KUoOlF;9n=OS@8EHbWYcWhPG:Jc;=a`VQUXq;jH:^
eQDgli7VVQ8eNT85K43Om3iI[PQngNY48PkXML1<L@>O2M3`cbNFC[7SNOdG2Y>O
a9gWnaWYeZVYNJHLP73<m3KW3KH[Y_RQDcVH=Lkljb9V_P\eF7fE=V]j;YZ;PQa]
a@gWKiH@e^`YN^HLP73B]=>1ap9`bAfdF<R2[7oTNQDT2@_F7@aYY76k^091T2an
Hk2^N8_KU@@Q2Yl]UZ^alC?i`W2L=MAaMh<gP`f1Ik@Sod\6FH[YYRoU3knLof>=
G<]=R2Mm80RI_W<ZD3cFCNHcUQ9M^Bga_D<5[mP11j@SI`\6FHeEk=W=qloifFcN
<>A6XR79gIN<I@?mQQgIJogSX82Gl>\TDmd`=OWF2XXQJ7;mKD1YD8SG\Sd2gD9H
=HSYI`fNIGcK5`ceS8<9`lmqi_JYeKiSkE<oH3N2h_9>5AC0YLIm6A`C1O=Kqf`T
lKCpIGUX8\\$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA222P(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
_d^RlSQV5DT^<OZKOP4RG]B]^8PY]1:SM>l4Dli7D>F8\aTnM7Q\oC_RRTFV?A@i
iNaMN4FoB;\khF8pZS:L6oCLUdRgMFI0dAU`Mem8UT`M[WBY]YhI?dXfI]XDK<g_
fQp1<Mok?Vd7HVShDC;iB7>Wg_IG<[7@?698@q:8n[fGp0QUiQFHSJ5h]liO]dcZ
;Eb64dG>[EE_?Mmpc0`afVOGK0TTWGAa2Ufn@42^2>2:j@a5N1pg0Dff7S]W:gT?
51FfHe<:`>0EBZp0LL5?P7eC2ZKoWYdF2eC=Q7DDZF^2kSabLpkU1SWOIk9K1HL_
QF4GHY<];:Q:o\4C6E;]A?Ob:8qa3]>9^[V][8E5<L5J_?:AeA=SPp8Ghg4Z>q:b
1:G6pTEoIIXMC3?ae<iIZ;=nCgNY0?Y<VcN\]2G@Y[1Xl;iP[O:S_fIS]GM>3HGf
cbmM@i<@UOHoT;]TYO_0ROA9_QcO;B0n:dJZ:3K]IC1Xb^UCgVedB9PM_T3<:jRj
^:mFmN<A_OcATk]kWO`oZOA9_lW<bX4pd82\=3mc\\7WUAX3]h>gmRa4FEUgI\pE
XnNN>QWCBPbfJ>R9=FYJIcj?lEQOc5^4631EFdhi6Z?i4?7Njm9D7CdR19PaB[63
6VmQiHQ\fH\mFfld>fOS@jPmlE\@YW8VmSXc7oc:cZe:_S5Udmm4Y2`3nKNK?4AE
k_\7i_=\BPZFF_adDkfS@jP<SW;4=pE:F`UkWZQ9V3I8lJEcMGbWm8FGNjEgnM:J
_kOi9:QAibU]6SQhcMjgI2>JPkZhKh4>VNUU`E`WY1B6<8eH=`R^;NPG8GGMOc0o
EDBi062M3LhbUR]S3kZka\kU6Y^VT^M>R0UBR=JWJWB@GGeH=`95jIb2qnTR1HeT
C^P>X7P00PP_mTcU1hE950U;JS6cZ;>B=f_OQ3gJ@SZ^FYC0EZbVhVhjhL[BJYc_
aO7TaaCn1nbdj;1eN0La`[ADQGadQ7>7n<ZlX=:V0dGcB0M]XcXnP6<aSj[FJY5B
ej7[EaHSWnbdj\PE]:Lp]^<i[5S^5F4K=94MbUQA]WKISBAKbYgbNDo8=Fa<N]`S
Ca7n13XTkkWXJIT6U03eZ1QnbQmp1eFAV?GnH=L1:[YHg2efQ[8kb<>DTe<TX;B_
8:^R=?13W7CTeJYgL\_F2jg>KlYK@ldS5KClI6@j@lG2>A350IRA7<2KSHNc6\NI
>Q[K1E5N@\1N;1l`>650^SX0`2dI1Dc<mKK[ISLCFl9A>o[h0IRAkCdMJgp55L4M
2`o2\j>OMUL^DU[AL^6hJYB<k`L^d>2n8BeECa;hVEmU2263eL7`PKggNK`E<8dR
SU:GfH\@T9Mh5ge0RT9Ef\njVjEYA:ZA8fIA=2K?[4o[\`[V6DEM=LP\]@fm<RgR
RI3BfcF@`n6h5geBQ0a0nq=hoL2>Z:aOB99=:JAXK>dNQ^hMY]hHZY^U>4mOZ^`5
A:oPMTk`9?_i45\6F<^UXZ:K73nSe14ng^`Col3E]j?dhIV2;kYN54JTf7cO^EXF
?Jn?^R2K6@:MYQRanlT0>kJKBfnc6?SnHh`D`W3E]jEgJFI3qQ2S=K7HGJNRR;@j
^;7eA8G6^?>HdCL5<beCQ2Ca]C<RFDB:K;K\SojKJ:Ijagj7?0dOF3b7G2PNUDek
SJhVVWVf]c>ZJMd=O\hi3Sc[OBCoFQPZObR]Zh>IhXAd<0hYjQAB6:bG\2?Wa4eN
@Jln9WVf]P<QTi?q_5G@bNU3l]`D:=FAMSg?aG1Lgk_gk=?>[?0@ALiCV`UidIgY
EKDg`eJ8Q2ZUCk@eAYl`@iaK5BU0<=LZM6M^gmNcYkZmW2mVS4m`>m\fdmlH147U
=DM\cLNT2N\X0^6Y_jM3fi\651MWg=I7MV3_gmNc9Xh6S9poZe1o]HnoWj\5UCXQ
0E6VZo\okp[\UP7H9@Be5LMQMNR5NBdJ_7d`Tn3HAG<[Q]XO:mTB1\meN;^BA4[I
K::2==m<HYIK3M0jHDJfo@j>bT5TSX0LU1?^S_7Xp50]=SCZ7E\=iN4HnkoE:5Mg
OF?fH@M3KN?e<3SFiZW<l6D7<D;1=gN5_QW1H2:ohU4M5NUAF:<boO]I7@MZ=1J;
Zd5P<WCOTK=aMPSSL:3NE4_=mFYY@OU>L`0L=YBX2@4aENn0@D<D5O]G6@MZ=4ah
?jbqCa=iEgIA1a4a=P]e3joMlF29gd1?^dToI`;1Zg6G@@OYd0@PlQiIDMkmoiRd
0Vi>RZ707fSk`P0fBjB@8WaGbTeKkhQlMXi8eJa9lg]1c:008nGC`mD=eC5_DT9h
Ti?8[ZX[7V_U_Pi`Bj208WaGJINkR6q9KI:7UkfH1cb_e]^U9bA<aCQY`Y<C8biQ
>dQ39loL<e8OB;LMc[HYBXacHAj;GbNXdmak7gdJEkhJ6C>^gA9UnGgk`Z]l]CTg
i^]^H5W2in:dog<5nnj1G<\M`6lRkQX9TcVQ74]JolSi6YE^gS^UnGg^NVmn7pXZ
=UMQF97_c\Ibd8fPQIjiMTddAZPP:;53M8AZol\`d=l;Y<[<hQjJ9e_IAHD98;nA
Dleb[enRI<C5EOL7XVF_d=X<KT63f58VXeSZnomW2Y;A?1FD]:R\WUYC[H9>?\GA
hoedQCMR?OC5O^L7XV:?H?B9qo<aNhhY1c3;:0fW1]UL1c?46Of9W3aa_RcXilic
G1jCD`o0WWm4MAenBJXL@4@<Z=SSc8RdEHHKa;55ILULBkYAB:fHTO_ZWhMeZD@3
XJ^:HF57D?\2?fkm8KQkXILdUoNW3bREDHlO^?5n]LUm5kYABi;EfXaqSjn?c?U5
MPaG<g5YM?_:A@8MW]38EM;4k;Q42Z<g;n\dOKq[SgLhld^Q9FQP?23FXTFka1Y=
`<ULYdJ<D>DS?gid20HVgK@0l:98JXO=0XNhFd4Y@JR<ZIaT:VO?YLioKed3@;Zo
`KU@8KmS4OG]ZD\XR_1Hhhm07FdF9Yj\0a[Jm9_[eooEZ_PT4FCLYWfoKGB3@;Zo
l<DJ>pKN=2[2dNo<[75n`2G\i?O32[oBYmdBbIF:h`f:G\_NA:jQFmT=8\_E:JoJ
ahLRNk@eh?W2gf5mheSP`=>nG71<6k]B9@i63S73oS9R[FU=AZN@RkKOUXM:\k9l
46F1C>K]1nd2T`5@<PMPG=>n981<6kiFH[Z@pQomINFagB@eZJXT9\MOPdonfUhb
DO]Ym4L0MAB6TkKbWnB4jDV7]Q>9?MkogFEQ\EKJUEn[06CgHi2CGFHF;]ZofSh9
Y[BmV63APf]hAo48`0e>5jG4c>SDA=L1fn4fAQ829Cn8m6XeHY22UFHI<]ZofAT:
lODqlfLmj<T_DgJYCW4cBDRbY5:4M3QU2;^C[ZS7NNT`C0VC_YJJ4fKTDh]M\?lK
EME6<PiNLoUh`75;fEHb[FVba;cHP3e4d0LiXN;[U1oL@iUUOS8ABJ[8>XNNJCcA
4[^4l<9kloPL`:J[7Edc[Fcba;cHcS=OVhqc:eZGhcggQDg0kdBWGHhc>Z3:oSOa
]mNVl8l55<7;;5bXKoKmCYkMlD^QEXbXK8JU57Aon37j;Sa2L`G;d9P:bHF864]R
Dp4PJ]U_YFDbi9doMBRh:W=D?lMHglS709RQk2YJM_QAXX`<KZE?VMjo[>dJc=9X
5GMdc;M8bZk\kNWbXe0\27aaB[6H=d3S2DgbeX>fXABSX7[IMCGWI@J2_VLdV_1D
]b4Slkj8[`kWi_abgS0h`daaB[:W>@_9pW;HdAA>4Y0U3_L?daW>653oQTKn:2D5
8`[?1T]6\EEWKQ6[YD^j;@Amo47Wll3>@78Q[lgAA0[aQEd4M9EjETe_\SK>EDZ5
@_fLT@ibc]W\SP3CJHLlnAB^c]gSg^=W:WTLo]gF]0EG[cd]I91\8Te_\lh_JM>q
CdDJ<BUMM:;N>Vm2S;W2?\0koiaD71Do74oS[o3bY`m2_o;UQEl>U\3>Pi@MdF]7
RK\;[OH[qO@h2Z1H_malN[31\S]giG4c=2[m=j0UJi6`6:BbGK48Jn\h<6L2?:2K
AJWm3a?ZDG?e0PdT3bSC^OFGn[`2=cA9<e[DDD`^1fL\mkkI=WnY8`9f6;LL9hZZ
2AmmLTAE8OYEHOd:\bml_4F<k[Y:8cA9<jHmA83q042IEHm:mU133RJ5JW[gF``6
nUho1o4PBV;8]kLa>BBIhdYB3mb]_CXXmo?1_cPLN]6?3X:>5_<b=U<b\<`VDXkZ
5UUm4@f@23EoG0hlaA4CGBiAOhY^I\<UH76JS_9a0mYIXXZ]5:VEFU11\8ChDXkZ
]A_[jDpB\Tmd7UY47bD[iccLMI?hXXjg^2GSB>YWFaU6TH:h\<hYOB3[1G9]Y[0[
X7\2i:`l0X=cEMZdgGOn3olQiQ@D`]YE^2`X]>IS161m?Zf\K\HCK6Q;d?5PN\G@
7N8\D5_B?<FSEJfdibK>3n@Q6<eD`]Y6k6n8kpa@QjEK?0hIGSXY`V;[<ni0?i[O
PcNY=REC9@LGiP[KI44jm7d3dkX24j6]9oN[>nK?8k4YOlEceVWFR9bKBaFUmB2O
ljFPTm=:\hgbZ>n<_T6eIH6G\^DiUK1nlM^OdOa84mLYA7EEGVXFd6b2]PFUmBLN
i_V6pS1f6\a<X2]K=_g4K::]Ja>?gK0O`2k=IHi8?MU36e6U6;IRD?72NYTDFPYD
5QlnB1_g1m\jfXLh49O_8D<Jg9S;TfmH<gbRF@::8MUUIY7BeB=P`d0d;3YQoo0P
j6DAFE_7ImX<YOL5T9]W0D<JgFR^aM6pV4c^Ub25Si_9Z_o12VM8i6SkY1BM;_oL
V4DXO=N45CSbVV;9\WaETX@m]U044S[h]kZ]]hCcM5=NKLJ[04DmQg<?F1D>RobR
8>3I4ii4fV^Y3FLmFO;??_3k_FG7ni_:VD@k4h[VM]_gNLh\0DbYQg<?C[NXbgp6
O\<U;<2jRedAHWd:nXgQGE1ZIK\h3AcgS_8lnDIkBgXYIVf@9K:_l89?<i2^^o7o
TCHFR8h30l44G4k[LUn>WXHUI?1Pd?ldD>mg@A?U\<FOdeNG2Y5J\?<ajmP1;AN6
V8;:R[:3:NA>GMU[l7K>WXH=E2@HmpZRlh=SIZa>35g9F;QegCXDedUZDp2::mWN
9EXi>a7bm9>O:MiU4588oaNef_OlFNX@ibC[iAiPQcPC7a5QR>aLEEiMgNR=TI<V
YCDb6TPc\KEC>X`i62MJe1@jqoD<66YO<cBWXhVX]DU_2G?3Ko8I0_QRUm:T^MH3
A99e=PBhY:m@O\d2TSMA@:NNiTZX_c\K6WKfEE\`bJVnIkghQB8@o3^dPP^\Z1C7
F4Ke@lH;e19I0Q;KLA`KS_YmfoG7cK\[hWFW0o\H]JVZIkghQZ<_D9nq\@@ZYX?f
PY\QEK1mNOfgJ\_\3X5ZU5gKG[L\[9>`W;8lEmT<4_\_Rk1i07naR<\SV>=VVU8H
YXV2I?c=^OKl4?8fgXm>V0n81]HZIf6oZOJFOWUUQ]FJn<FC;3B8[gk^\=kI]UYf
YknIc?j=^OcW4?8fOmZ:o3p]V?WEB6DfFTNAIn6ecQ_3_Ta0lb_<AEmN\Sh6Sd=m
>GmZ[22>A2E>1_m6:V`\G6OCi[Zd:O_e\NL0g7EVcbRR7[ROld_]Dn6\K^X2T9==
`gHg7XMDfhKe0;gD\FF^;M0]gXcG:e1eUTRUgAEVc1LR7[RLeAf\TqE79\CVaghA
?W5Njc_hml0?ElGCi8I]aEbI@C[8N6:Vd:WKOSFH@F\MSCc1MCS0Z8V1UFPI`iko
Wdb:fCdKblZ[oH3D96jmeK0[cVX8O@cm2oiVFo?L3R1Sm2GBZn`jAnn1h6PmbRHo
5Lb:ERdKblO6OTQ5q0`L_[X<H<Y5Df67bZg6Zoni^gEfW43j\=JHXPd?Yj@9Ki6F
YZZ8eg<ZFbE\L:;A9V0SBinQT6I]5X^dmd5jM5K_HGEg<9mkOZn0kG@DWm_9C_AL
V=@gBNS9aHhM[J_3l03ao]n2:6O5YA^Ufd5aC5K_HO0?haEpE@9oJ1?0G;==M[Ia
;4Vi:e\PQG2aCgENL8oGXM:BEm7j;XbGD3kJ890G_Lb[857NceBh^Nb\JA>5d0`D
Fl_X>9]haGHaY;58?H\@_>mnk<JTm^R:j1ji\R^NOh:`g<O@EH=o]N1PJI=590Gn
Fl?l>9]hAgCk[0pfL8HfkB<c7l0M54@^@`n[G`d7BB4bN5^m6:R_Bemid1OD`Sf9
YNd`^S1IP]Q?BLgWJ6Wf4FWGiXika9g9][i`c;5>B=h`O=ec27^HB0A5:RhFZ\;B
kG??J2dL;gmjL1:mJLWfKEH5idYka^n9][i]I=TB@qK0gLSLBBT9e3\ZFG[3RU82
IQhA[;BE]]me2`80NehMAL1S95D_i5;XFgZlWol8_S@YhKcCY^lVL;Uk@Y63[I38
A?OA[ChB]nQOm]l>M4\ZA<Oa9:6_blY6LK2d4_1:bNKilO1CV^lYeGnkFI63[`38
A?d;Ug:_pG@AKLVIfl<jVl8ghK7CS?bC?7=D?9UT=WSH6jW3?ShA<p5S_QP_Zbh=
i>o<L3TJTFRSWaR>1Z:h6\NeanWIUKcVY?^F@oVGbK_DQbXQC37Z@TZdfTUnc[H?
HDG<?n<\j:gcSf3>PVA^0\@ENcHk[@lS`H8oa<5<1\\9Wdn:gfk3GL5]>emn26Hg
2>1<6]<\YMgcSf5^^CeTpT6XE9BEYT=;FaCN75a=F1Q@0jE5:6hRWCU8kcd`N<nA
Ng3Z^gl[CJUU8cBJiHfKb[2^J=D_lVG7JBH_A5:8XkF_J\]H23QqMj8FYYn0j0f>
=F6hofmgmV;SDnnfSLEaD;=JT8?HM2gS1CQEBmiBZ;BLfnR108Sg6I8Kof7:Bi\]
_NT5=k;2mnLl7nP?oH4QoI1nE:LG]=mX>?IAVeJd=NmjN1QEE24GMO@Z[fVdBAY^
[N^P=>@fmnLl[PW972qm1d`7ab9nnZZaOflf3fCZQP?RH:RQ:5Lo56:m::nc;a]i
fd\6J?PnDF:Zc=mSI]a2_TKW^7b75Bj4n_c4HBGj6K>]HYLggmdZ3?U`XY<BjC_6
o[XQJb4R?mDN>H[cJSXmLeBP^1=7MZG1nAG44m7j6K>6YFIBTqmlmPa4k[GTOc3l
TJ<m=]5:A?N;nGf@LaK==TWad[f^?I5bomT2XDWFB2EoAJpm]5midodF1SYlh^aH
=Phnlcj0BJF=MFj1B?k_VD2@EL<1df8N:S_NTM2hBj=CA;[GL=Zllh852_a48MhD
Vjnj>>?bBgWGn;1ldFaR73b>AL@aj]C]mlf2B`n6S2?GiKjmHi93lRU58B>f8GMD
[ZWj>>?GE@6B`pgQ0U1JoG85Jn7j6;oPDWSJH;C<fV4D;7MiXka]1EEkk:HkZXhT
\@gV0NLA3@EMogcSCdi5_k2mQm<`VKf@BBXGB>2<a>4M=eOVdkGocF<6Go2`\mom
6P1f\L^MlL1E=fgm:Z25D@25JX_`J]f]:bXGB>_P<`AXp3O3_H[1SWh6fIlH;U25
=87k4Rb?Re46kW4[M1F]Xk;A=3>7n7P_O`Z8@RHELFIlQ_bNXSgMamELEdBYQbl6
kTf^1YbZmHo>TEjYZhl8V=DQHQdo^=P`Zi2n>G^Ie=Ja]3V=;6gmQm<PJ=B:nbV?
eTf^1;SokYEq3PUlkBKnFB_i^VFLW?Xb_X4H6Q]MmJ3K3UJZjj4J_AZ4UVMi4CeQ
4ndK5m23K1lI8aJGD7UjeB<@AgSZcUNUo352TQTX`?68O>fPSoP`JG6BIN>c`238
gK[=ecA1RS2a3\TP17P9eF_nbgoBc4=7o352HYXlDLp^eL46C1ck29bH2Kb9jVG8
e913fHiXFAK38@\T]bbQP8SRRJmQ>oJ>lUeESAD\Cko8jXaUYElOB2UMEflS2J??
1>BHfRE?mGam9L1ahIL`;=3n^O4Xi^R^kE`WJ=OI]4g^gSWFYd=O59`1E=nSXl_?
1>BBfRc>dp:UVL\i;NWF0lMb4U:kG:m8L2kXMeW[M8T[58kCU>CNZF>0nmonCcni
aKHmJcH;cAS=IDP]P\i_RH1iD[oGb7^H5Y1fl[\cRcH21:hCNgO67NcbXb]RG`7d
FYO6:leMH^:=MAPNAA__nK1>gooGb7G_\CIep[0hQVojY0ZjWEI`NB7Gm9k>p_aC
69>QfBGHNYio7Ybd5;:a^KMV3:S?l=l=c__`R5430>E_kI]I1SFadFEBV6MZH\Qe
dE6ikXjUBkZ3DVQWTh0<W>MO>eXdO;M1nU6TIKb3Ke21BooYMee78<=X\fZ3O_L?
Mb63KX5HgQZj>VP[Sh0<WPa`gK0q\JMS;V^A<o6\5b;PO`Z8cO^Gfm^;V33`F2^C
cmf9\kofTPOXHOah[MhnXPl;Ge2n`Bjco13QLZ55^m:TQ9IBn@RP1>ei0cqXDo=n
UU>^0Ado>fI;Ph;dKlWL6Rdj>43[7V;]VGWZ9Pko7EE:8`Q[G:8IMj1dFZgOcX43
nA?SN@h[J9lSX_L]aL\36R9jAFHZc2;LW559Aibl=ai\RMUb;1bkVf<aeo]Xn1BW
nL3SXAkeJNLSXOS]aL\HLU977q1a9eGo6?5R[P2UVI07EDH`6=fBM[=gnL`CF_2P
HWe4J9nHSUcEj^>cM93;?\N0k[_S:h3YLkIG[HCAJFKHLRh;PK?B4[_3oTNINNPU
3T2nDbi?Z<\nZe;390`D_5C^j:1C6XMYgoIf[PeA3DKHiLh;PKZhea47qeX5U=DG
^NA`QXO11AgXAl1?2Lk56NUicDeM0H>@b\9=18EF][S`eK4X2fbaZYP[RTL>K;F[
XRMj;\n_LbjTLeCd`<k2\VX[khg50Vc96ALT`l0o9COlblXN5JHRbFJiFe<EOCF4
oRoBlKn9cbj]LeCd`2dhPZSqVWMl>>5Qag=?OHL2UOeZMhe[lcfWU4PnDXaoNA4j
JYhfIe279R22[4aD`4O4=IjOYLKFUF3Ac3m6g3F`]lQiMKkV4cf<bF8SB?oeSc70
Fbh59Yf5ARWhfDRB47AijSKdVJ9lJFhdcm?5832j]lPkMKkVUI@KFCq0J?@D;0ZS
kJnLMU`>iCf4edL>0le>o;XMNE@E;PA@C35FEO?SXW4Jmf9f]78Fl_Yoo0\A:Y=6
nU?AQb;Zh>BjA[6Z0Ck4Y@1e6YSf4n5`c3_85d`hDCCVT@]TUfm1Und01Zlg:H86
aJ7<Q\kZhHJjA[6l5AA[op2820<ThC4?T7UflO\nLkhoC=O3MK6:[E8nKMgXCT5K
?oN1\Nc0dmSm660SY_kZfHDR85HmOkTITCbj850YE5:mF1;3W>oWFf@>DmVI6b^i
>XNEekL:U2llKZUljjiQ3<2SZn9m7mTGTFaj`;0Y7a:mF1`FE`99qE^T@Z8oCOQK
H5JkZN4LgUECIZ;DaQN=KoXeON56>2fObJXK2bnSM9:f@9k5MH7VCjT:;06qgaiO
QHHPlBFka7TSW`ZRSao@Sn;0GcX<jFRgMh8hTN6:n>27Go:WJK8Wh<2cTWQ>ADF;
?E`RX4cRHH8]5nPJ7=BT8QdIZf^d?XK2lhco0Fd_B:me4mG8jH=`6e2IEY1WEDFa
?WRRJ41QHHi]5nPJP^jRk6qS_aaO\8Yj=4T2JQ\iJX[WLT[Td:PIXk2>DkJW2Q4a
YMi2L[hDL>AdkZ6m=6KFaYB2GWI4g\9Y9BM^hmQIm9DSDlmddjSUYNiF^H4cLe3`
;2XTlBogdb6_J_UNf01T`XTSf0\ngi]YI4l8hfaImbFSDlm]<Hb1MqbccE9K6oX:
o0WGj`>Ah?i=d>YncLdNdc4VTk8JMGiGJH;H09W<FnLjPfYT18W7B?V3TSQe=kem
oB0l;nS;O=CR7?InBD[k=Z_JBL68O?8AdhOf=foUZZiT]PFlEiXAjNb?gk3eE:ea
Gl8lCdS;5`CR7?KemN;ephnm2iC<AbL:hK1I6CRG;jnCn5lObDbT@]m]epiUKg3i
ojIc=X8KQIX<AKEenKh`gmXO1klSil@nfLZA_aB7mO@kdg>W0eCIWBoRG5lUIZQB
]0mf`j3<E:EGE908;B7R;:B^qo9:V?0q9_SYDDk$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA222S(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
W:`21SQ:5DT^<LQX47aLATJY>UlQRnFcq^<BQ2R\jbN<iG>eKd^aXRZfNQ^\5P4\
NW^:B;81V?gZ`T9YjdIDW0AFj=`OpBPNc1FSLP6^>9Z>[M2pP@T;;=q1BeJI0n@h
:jIMcGEhP3Q4_Ci[iDME\jVomq^ODBXcH=C52nQeX@W:E;F@E9aIl\E`a3X1pY8[
2<hGM9a<:jKFeg]TH=196hLZ3bbZ9n<p87mJB:1=<D38e?jYS^1`:LZ4Ze?B_HAY
>eBGL_GGpnlZ14H^FE^X73X@?hRYRSl6W;gi1_Z1HhWYI1`0WAa:K1_o<3BA_ZAF
X2I5UMhoBpYDPVJ_\_aR0Fl?kMJG<nQLVkCkp4>5TIXbq\9ZnXCpoRAH]?f\D;@i
N^:1YDn]iQTnOHZm9K5Yh4;iM@W0MCp>S7HQnCX0FZg9O?bdG=]Q[0hBG<EB[=1D
oV]KHJ7PRAk4nOCLj=ccIm2N_RWBEi`>R1\AFRPL3gJbEE0cHZ4=R<0Q]8K8:kgZ
oaC@ck[HQeT^<O3DakI6POj7C6[<E[C>Gl;VF2eLU4RbEE0]][b[_qhVWME2biGK
`;K\PD8g\LABQ7VPm]hP6X17n[1[f_l<ibgIaWLPkoP0_f\H0M3m1Oh4gMZL]1HH
eR2bU<3XZE9g;6B0kVM40_G7n8EmYNBZ[TnCPLk6]KH?C<8h`MZmkmhLW7FLAcH_
O22bU<ViVhmYq9\?G?i]ZfiQ4PG97c:=odkl;lR09`1fST8FiV?UM<hh^@E[hGIJ
^gJ2`T5LjVL1e92T7Lm5YO^AedV?d2YPjG:VAMDL4T7UEB8DK:0163f:_50l56<D
eZ_JXmU^FIL3f9GDWHm_QOOPcdV?dDoHjAYqUmg3ENTn;<5?F5VlFa:Q97mZO9O=
H0C?U?B5XD>B2T]:UG;j`n1OY[@dV5C5;Q4oUj<mjiNYkihXWhgF8DL=Z1dV\CP]
UYGWL?cKKg:I796>IEjVZ1l9YGHHFEljOQhWUn\V;i80k0KXWhgF<CnJM7qQl7J_
2IYKRSgaAnYF[<ocb4Ia>jYeLX8?FGQnk5oJaV7TNYTh<5X\UKQZdFdd17aQ[m@o
WZ3Xi\RF[0A^G=YNn]3903hQPebkF@15jI9MEgBGbiP\i5c2_13W]4HF1oBQZaI2
WLOXB_AF[0Am1[1H?pf1Mg;aK]fK8HQ:9K_LHZ8<ae4\G]\mY:Y:PE65F`SfmoIY
8lY5Ahe0CfT[D6@[]]fN2EDlCg2T`I`FS`f[f6YJ^>WcQaYWDDi:P>D]VNBm4352
9hQimbi1^YadlGZ[XOfmnZol\Z2VJ:`FS`_cIWC[paGX7_UH[E>_\e3=J]jm@UAW
]oAbXLgbgZL8XClQ^2Y>4qAlcF8KO`0_DO66FX^kkfEW5VBKoVMCReTSAG54^80<
3OLNh;LT\P`N`\dj;b:iH:ARee9SjB9N`7VZ0;I\T3DEb=cmgjQ:Dh8SESUA:AZY
F@CQiMkC2kdG:7OI:R5iHHA<@6VSEF9Z]6VZ0;a7OVEVpomVPQoRUM>oWRcVg7oM
oMc]Ub0L]Q9c`KD9IX]cJb?_lP6f;NE4QDVP0>M@k63m5oKG@i?dlQE1Q]b`H[HM
di3a]M\`Y0Jo^1DH@7^[i<QVMnJ39iOD75QbJGc2>33FaoSF66?A1QRb?]b`HY7T
F@nq\c7:=3LNOF:]d6@mPi>Z_:he\ZjU=0j90UdkPggIW;@_RnVB20N[1XV@n<3?
cj9G\[obMAZjPPBCGC`V=DPka6SV?8b79PTmUUPLmY\=9Ii@<BR05ALoVLCMSPo>
RjAO\`[c=AN@PTA7GC`VITiBJJpi3;jGCF`3RUQNfFLQ32gQL6W_a4XjPbHjWPA0
g>S^d0G;OnSB?WEp=;Ua5bbkN^Umgi^AocL:<HXcH:Tc4bd8=SW88G^c:dV[0OTR
]?o@Z]`R\XonRC65=P0QcPlQ>I1o\SkXZ>8=fUqd8:H`MHRcoifY`I_gINRieoEd
`SL5X3SS3R]QYi[Yc65g9U5T_k:hQ`<RZOenl_c1FGEVX3P75W@7@0j]G@N^TTKX
^YSXKBS1MVh8YBVJ834[V4AT;@<CT5fZ08hFXM`dFhPV^==956R7@Hi]G@NVM=]N
epWmI38Lo7g><A;i3oA=LQZL0ARb?K:23e0dEBS^CMTg2>0E7mNKB<`g434b6^B=
K?WLVWY74X[2[eeNdnaQoIQUmFJCB5TU319DUUB^C^Z0e_jn7lAWje4DEW1JAFUG
>J:LhMY>3\E2NoeNDOaQoIT?\H\Ip\lXPIV2\2L=e<:WdP0`QN5I4Oai7CG^1DT7
M0Z6ohP_?bdQFP;0Q>29\cRd;YFQk?FVOOPYl]ZcO?<_E5]HMPLCGbHjHkLWTKk6
@FZFR7X1hc6f1T<AiIgLHHV8:72\PmF98OSKV_ZW0?<T65]HMb5Xe[1qca>^:IRK
f`HUJ[aN^iW31hWcA`DBK;iY4cckfFZ]oV@\=KMVTZ<Fa\TK@gZ:9ZE>:46PSNTi
?@SA7]GK\Pl6QFjRN]GIdY;DL27@?FZPZJOJoWoJlB><NI5V^AH=K?Y1i4m4S16_
k@YH7]1R\Pl6WFhccnpA5S4Lfhe\3=>ZORm=5i@n5`aa@VRk:92`o@]:]KR@9D:k
SURLA3H<ooS0VAMh^ggM?o39:5^4BFQ]OClWlmg7L<LadoUEcOo1O\Vj]D?2L_Hm
?lfoB`OHLZD:B\Bl:5QV?4]9nl7XBg_]OXRWlmgon49jKpgkTh^]Deg76A0ff>l^
XeQJMEBW4H3Sb=aAXe2>Wbif<eEU@SLab<`l`R`6h4TYE`Djl^eSW_WeEbLHJT>U
7fU0kkNNGMf=9oLQRW[>aZHYRaiU`jGBKomT>4e<OGE6430j]?e`DGTeCVLH@m>U
7f4hl=f4pBOPbI5g=YZ83^4ggAbEnm6;]M^F^JdF>_8^Y3Snf7dQX45_ol9N>fSc
l;O1_oHQLROg\K;SB1=BfW\:7\^bhN;N<1FSa][QZNlB>FSie`Y`]5noCQcaTNY6
LbBWfUCnTDOenK68TT=O_W\S7\^bh4JP>@mqV6`_fl>aRB54c1b\Fano??MM6IjA
ieo=>NP8R>b;[gEMcfIJFG>[LhTdPZ7C_kCkJKWSNE=YESX:B;D5X4[TB9`O?Gk3
Y=@5>nhj^>180G^YjcZWdgYcT:MI4YfPQ5@FjKf<NgDgnSboB;IIX4[TH2_A6^qh
F7joBTJK3N]HQB@C6bR>OAAIn;0eZN@^KaT:nmd<=q=NRLLVBl_:TJRbWZ80NoQm
RIJIdh<<BaUERZljgUfCDFPU1>X=QCcPNioBTFQUUfBoWal?j4@<mDhO\3Z8[2Pe
=S7H\XWUea]9?^2jidc92Yk6XNnC>Gl>fj[eG:JOJbLojClCjGP<QMhO>_Z8[2Za
2eG9p1]LD]5h7>Ud<5J9KZ6KP2MEGRlQM6K8C=NK8XTe6HS=LclSkGg2K7`Pg7Ql
]Dje\PnF[feL5O3m\dI`EiE;0;LFggEp:HJ3k1S0UDhAC>R`k6ICnY9R_Z<W>N\K
`9e[holMPG[l\[ZoeL41RPN=:DkL?`mk?HKD2QddNoI65VY61`2n]`6nRkQX9T?N
Q74]JolSi6YE^gK9Ui]dO`Zhl]CTgiK[^H5W2iH:dog<5n3T1`2nGPdSW@q6BN<=
gY>C[WGBKe<;KTiNZiVi:d0D^6P>h4E1^Q8:NYgiMDjCdU7iMRIC2HfNZCkA=`WR
n^FgiDd6aBX@Nj486iA^OKk_eO\?<h?M^FA:k7nfW;8dYJA2GW3UO9m6O9i:=EGR
fMVoi:l6JlX@Nj4kSD[8?pg3ejN3_UFaIGi`oc4CGcHQ?GeTEM2PYL2SG5VUWT=X
qST7<O7@6JN9ZQg1O8Q6Tk;=W[@C3Fh@albScab]F@]GnGH^3hT>H<RQC^jd]6W5
NeGSYogWU0[KJlEFJBBHh6>d=aGQD2\7\GlDDJbd`G=fUgGRe]n2YBH:dU>h7`@F
Y9G?Wom@6O[o?lDAgBBHh4i]H\TpVLFBPC5O9FePheLfh\\4k00EjhM`?aFgooVj
b6YeLHN??\kVGb:WQYQ7KdZ7=llcHHLeMPGiWknJ>:_WH`A?3hSOcD?h>RTP?RA;
d6mlibdS^<l:4`YXllKSP=^nY=E2]Ha?McBSQkFA>Qk3H`A?;ML@_[qJ@dgcFI47
^FAK6@P60]h`O5_KXU09Mi?;37fKk`^FLgnCIk;V<j;U9oNIG:Zd_1?cXAQ0Qf2F
8TVNNg=V>c;06kE24_beZ6RJGS0Tk\:;VlagN>?<Mg[TY\?2PFQ?`:eXX2R0^D[8
882Ni<DV>c;gc1;S5pMGT?:HW8[:S3VDhDXOfAG>Z2>;heKgBPRY;OM[kRI6aVG[
05jm[QD6C>32EjoamHIBi`PN]dnNQ[^ULKmA@9VUdTM;BZX?L00APJ;Z^HMC:VP`
XW7d5Hi@8jHh2AFM2iM<`hYN2JngS=6UdAmWb^VUdTST4f71qgH6H^N5WSVG?^A6
11X7Dle@eFCP@]=moV^QifUfWOY@0f2JTf<AkI\mN5HTJq6jCY]h]H`k<V<T]QIf
7\WHTLgfkPj7T88nHgABedL271d@;S@K2[7BF;CDkg5Y\U4`0PAheAhPTFOQZmfQ
=8aBPhSWCAFd7:`mXbWBJ_=ZnE_7jQ79KU7n\SjX^Hg9>>Y`<fAJUimPZdO:nNfQ
=8>Q61O[p1066V:ZC^oEB1b25leJl0YXZGDB_SFDTZh[fQZa0nS[hn6JSHi:R1[C
^T7n^=5OM`b8gJ`:kLYd[0mhKQc6gMckaDfHdhV`[MI<aWZ0J>XQ:FX1MEf>a\3Y
OG@8f<S>ISbKiJ3Z>cY370=jaQc6gi9agKDpVAZ>R0gPSoFI^Qbi\1f<?e\YXKZF
OWOeeWQ7n^CgXm_cEI1Bm=Y=Z3MT78]EQ^k7;WblN`;I:eX6R]4MTYAdOoQDD70]
aWHDhf9]0^3Lj]DA0e9`d6]jj88MoLKP[CIRdW<]NTd;TeWQRYjSTYAdOaYi:bp?
a4eK;JhLcYMIjDYCEg?m=8al5dJ]W1DYkkJ:hHC@TW2V<X4]0g3iCTKUhWk5VXi>
B[ES2mPcZmKa6DK5<`R9R38ZBpRk=A=^7]RiB^a?K`O[AKe>MgYol7`0id^hZXgE
52>1<k4bHD2Olb__LbE?:m@1W@6G>alHnK7L;;Wm<P9[m_gdcORE\PSCmGnCJdUE
<dgK<Kd>IE5b25oUFfj8_cbgK:=GVolPkF5L[>Wme99[m_]e3AD=qC?4iQh3hfU3
\o?W;05U\mNF2<;JB5I>dck^2Fo12ChCL<>IdWFIL^Ll^S6WhHn:ULoV<]_YT1<I
1kEK]TS[cbLWjldJ3JS?k@^PJJoQdDT@]JJ`[:nV_A:d_f]R?QKeBao\5]\SZ\<G
YkEEDTS[c81\kRhq^WcLcnf]>D\YU>JN2nHb?@7IE:JRGE4;T;8d8`iJK44XH2^U
gUQl[PU3LaA94jD[^AO5=34Tb`R1?S:9nGI^T1Nn\O_WU<LPElCOS`hN1EZ;mM]a
Jj0C^lW4\oQj>Ieb<AZI=W9G^`WD?SEDnGI^?>nUh_qQGdi15SW0c\E4g0eA]06;
bE^o6>>n7;c\XcNG]gX;]:3C\>lIemIQ>o9bb@L>`\n[Rh_Y@@h^nnXBBAQCBhcA
Q6^HCYTjcXGN]Ble]OWDiknJ8V5=38DNeRRmCPJQfWI=R9^YcoONna[BBASCBhc3
64L9IqYZ5:ZiM]KLc:kEGGd6@715[\Bhg`mZIAI6ORYkH9obCRCJI<hURN1USeZ[
DOOaoRFngSg=`0\QAN5DHoc:bGj_fcRH_@158KS;DJ2kBkRMNQd>lIInHH]6\A6]
0YSkZ];nHbgY=0>Q8d5Do9c:bGZHNnFBpRhB3MiQSVgNOT;4FoCCU4Eg8WOM8d=3
J5FPEe[P[F9ClOISKhfl4M>L_MTjb\km6>;fpCYh\Q`HdeWO68eE4eW4\0Gld\CI
ai182d183J==Yj66P=WO;CXKJ2WkPIG23_D^YHk@M9jFlo[UG\5BJNen@f7kP6Co
hZB]A>\Q?lhcED\8oIn0WYNne=`A73O4F?V=jC^k:bj]PokO;>5AANeQkf7kP2ED
87lq3GS5SfD^J9eMVenY@F\N=NRfc]j[0LFgeo`ER1ZO=gH:AjQNa9IUlZ@`=6Od
@9CUDMCn\VRO]lF>JSUoP145jO:chDARHo34QcCK117D?:53_kche1DNIcODlHdd
V8ESXMH<\W:^Xlf>JS5oP145OZi3lnpE9e`K=?@noXd=\i74T4Z=e=A;8XQ5dNkV
R3:0555jMV:4>96;V`l6eN;^5O?[kT^2FNBP=bT0lC46ej;Wc14?<<`dDHl?WD2@
^hji5AMmNP21:^T^5hG_>a=6ETSom7MAFg0PM>UhljI6eoNWc142>3:Gmp?<?g1c
jGXZ`1k3UTUVTPI_WkZ<II>T`T`B`MfbH8M:OYCZGN\I5JmSK6N2V0g4N8[OkkkO
bkF5L2<hoH0K2W3Sn5N67den?b^G@f7bHC5Aj>MoS`d0bJQb[T[ond>YUMSO4<k?
^1b5[n<hB@0K2WFogfT2q:aUBLi14X7=Al[[1EAZW4]gSY\I=iFP7oHUQLWZ<Jn;
9@kNXm[EC=^?XilYPC06VUIiG;=Pca<;6FHdhZeo_Gd>dSAqW4U5Zl\9G4hLM\TF
lmFLRlm7VMg9\O8GXXG@bcqgbal@_J6<`R>^^CLc=9C6Xl57PNg]J\Z1Hlc0AHDI
o@\C6a;h3FF2a3C5c9d^OH97]PSbWm:3@91AEU1G__f9>6LNTAC19Ki[S8QeA=\Q
UePo1lQ6F7>YAZbl?4Hi@mI3]3Mb[<mh@>MA4mKG__fI>bGLnqlNWl5dJ7ob@Y2?
5>jk4cW5?X[X?l\Zb6bD9iW\on^T`<DkEg`hnkOM765[[nER9aFCdIC[IlRY7fjC
VBC]EfIbF:5=F_f;fK^85<n\>MFgF;Q\G?diP]XTCA;Dm16LLVDC93Cc\FdYlbj[
>7C]Ef=j3J4[p7617b?3WVKL4D\\@lYo0`>[C=focon:LGZ\=36DMehk8CAifmd9
M;Pk98NP1\V0?XQ6E0\VS?c82YOR<KHEg@4cEB?[lWo[Y9K=a66QRmXZU[n1DW2W
`K=YDh9Ink05VJQRE0<AAfc42Ye8dKHEg1Y0eN>q\;mo[RVm0RWBDKl:8LaG8HAM
1If@bP24ibDe]d9R9fXlV4fbk2O`05Z4X1Gg>2^FQM_[_QNdd>S]Y?^eSYMWnoK8
5ID7Z@=H2VbUDYSW5kXQT0FZ<2dYQMX`2LOHQQN<\hH2\Qfkd1W^=??;Sj\`noK8
FSHZ;Mqm?JAb<FZ`;F\YGYNe2=9l7F<`jG=ck=YIj@Z0NMFK:=?iUB\m\N[KkbWM
HA2jl4a1imi]^dBK:6;VI0Q1nVmnBn<ONjdLo;]RdTC^N8nGn1EWl^8R<7<=367Y
WJCQclVWiCI]7ffZ:ASVB3i1nVmIe1H3CqB>ai\BCnB:KVQFOQ2ANQ]K7^XVenjS
DQDCVcYI;FgT3P`gKjIPWIgnbe=6aO4Ik6`T\BjkC\REVTR3ZSKU`WaEfj5W:cZn
Vk?3;cTIOj24lQiOmk7W>6o:FX:kdPEKb0OT<[jPCPYE7;R80:KU`WI6;=blp[P[
meFKhmQm^4Jc@eWZ=BB2K>3S>VS<[lj0M\S7Xib]aM=1Y2;iM?O:b9>I:oGMP@^N
Om5RjAThg0A\dCn]4P7f^G1GEhZ`4Ucg<kSbVYG>82_I6oknM1_6`69M`Ujci9^S
gmPIMmTfF0NT;Cn]4WOX:^XpMf\=ie0NAPDBS3=7J1YQm?l8d6E\N5hNOWbV_dg[
gEH2MMQiDPXeEOg=nk]Y\X9Q>hLlS[B7dM_=``l=74>O\YO:SAIeKN93Bh@UKd[G
SfC]eDQ9:3;Z`ecWaTd[4kKMNh6gSYV]>M4P`g@W74>OlmL8C`pbOlh8[:NhiFPF
=M0V5h>dEq1n9:Dk]djdSnF0IS6i77OH7kd:6l1l2`nBf[;_jCI@fJSaBA1oHSTG
CO\H\Nd:G;dM19EP>WG6n91UHIoY[L>6Tj:lD1?RLISM\c8_1C:>=RL80@S?e^ES
OdnGO1``[\HMX0E;6IA6;?1g\AoY[LHVnjHVq^RT37?:7GolKZf?Olo^hde3FLFY
S9?cmi=4BYDil3nQ`aC\DPhD:]N<\N^Sf6090R[TKIgdGVcnC`WTEJ\>7GdLX>kp
AZP8FHkngSIRbZN18gQ9mJTM8_g>:l:MMbPoMT7i42Ng>QeS0bjhjneEhLbckO]N
?f[O;eA7F;NOo@?02kgFhK^DogaM`HHlX7f2gT^SPcDQ@kT6d4DPHA]718KZCL<4
Tf0;;[>l3;<:o@J^2kgFg]cmU=q<0dWaDjZAGN[=3ldQ6bcRok4Sdg2=5V2McnJ9
FCBOPnmi\OC_7UheNmUQi;WW3ZZWkD]pP2kR6eJmW6MaYi30;HmU_Zn7MQMZ8i3e
<SI3>;<9\`c@l3VO8C0QkDn`l\7ZAXfU8=f_4P6?mMn:>UeCEO[LH2NfBQb:`Q_=
GidMmVn\hb5;Re^;Z^N>n5Mi5dEfZS0MPSCB^PNWm2MHRUF5EObOH2NfAE134Ip7
^5?<OljV]C6[cONX3K]]Nd:LZ0E^=?f5^8OcaON2ocAoD=CF]<dNd8B=@AP9c@Fh
]`_eXgnbQEH=gnW55GSL10VUNa4D?`VGXMZja1TK\@kFbTCE5F8;bKJlAB@aKM<`
]c:eQT@;Qnf=gJl55GS1i;>=4pm;K<^I1?@CaAC3YEn_7Z4K;LTd1U[=c@0;<YB;
5_\[BJ^@6b2PA>@f?;f^8Bk=Bd2^N8=cUU5M82OIJP0>2dR>POZ;Pf<RYe6EBiR;
5:CkK<<]D?dTdI1ZNR^49?B1P]`^4B=F1SbMbaOI>`0>2dA=hlndqOUPjOdIQ1@n
>L812f>YXf7S7L_n22Do?c?p?D1E`N?dk1?9@B;dI?4YkR:Q8k=a?BhFMe1<29VF
bKImND4ZRk2\3I<LfZGLJ@K^C\nm>6ODW7=RCKF[>MDRmOJIaaEcBemTU^3Ej9V8
SPZg8NZ^DSM_f`LMQV=7=7C9<\W7>=3VO7hUCKb[>MDRHF5>8QpSbXN9S><<P=N?
3XM>^SPW[UaE:BlBD]U[a2IdeWnO:7A9j33?jo=`m`P7gMBc;_M5e8nHVYUgo=cY
KfP_lK:N5Nf;:2kRSAlCMoOmcO@KP;Re?5a0jhELXTd>RoV7d7<S^kd\VfkgB=N3
K5\_l\dN5NfS1[;?=pVO5Jc3llZoJZUdiLdS>GJjM9nC5mUI>m\L3Yj;ZeO3nlM<
[n^FOFmDBlf_cIMA\9kIKQL=LJjbfD;KZGil02b>03C_lMOZVSag4VR;RYDL=6;:
JnonM?3kIJWC^<n^=22ILkL_3H[baa;Kkgil02eO<@2XpWf5^SZ8=dj5B@8E=4Zd
H7U=Te0G;IWEcF^nL\Z5AC9WDWS3RYd_1>7WoqMGT?:245[iS?VDhD6afB2>ZL>;
<ZbgP9RY;OM[kRR6Al5m]QHc8bF[U_:>kme_DSR:]1\j2>M68K3aedYjmPdZmQnT
90;@j`QVf[j[Lm;5Zd\4obAb^WQTVFX]MmS:BTd:f<\<@?76Aa3aU@YjmPMbX@R0
q;Y0dXHiSj6`0c\VcVFUI\6:[@hbPWL`O_1ag<lVk4hlcj20k]>U2NWJ3KWUTLal
VD]JB@DLCgCIL?Q?VWCoGC=?EVhB[9:@Cb@=[TkXk=3lSC`MLP>b`^X9;2gcA=l8
;;NkTnD7<gC[VVQ67WCWlC=?EiEdGg6qCd]j4^?kki;PKW3@W>BSX=_Ya8m99`A\
[[1hGfXY?oI42VP0ckc^EMm3]06bOBIU:2f:g?fSODV:P\VV\7g[>X<DjH923^pY
aFg6:q=3]M@>d$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA222T(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
XoahNSQd5DT^<A?YAXe]9LbL71F:0GTXZilMZC\^TSGTJIp4023cY:O@lKCjRTDW
EGmROj]7BHUj;HH54bD?^=G3_ncmOmqeecZMYa0T1P;n39R<in>2CmeI[GRlVJCZ
Oo`FaXWaCm]g_m17aVei;Y7VJ0DXe^mYj9ji<5q?RUi``p`l6e[D2N9HRh5U5OFV
gcB_G>Zik0UmlJOXq7Ji=a^nanH20loE]c^E08H>\jHOJ9d4H\Cq;o]1KcA=?og<
>kY9P;AKI<1`X^j7=B8OGmpP0BVV6;cG`j^^JGPPPc1d\Vb3S=@?4Z=G6`EKSlYp
HjX;^bChHnV9P2eOfaiW[eXK79p^8DZm5Q0?NR0UF`]TUDf2ADi]T2P3XV4g6;pP
GLim]Cp^ChYI_qXSb5^3CX`me]PX6T;J0ETa99QB9Be7an[f?8lEW7Q\ScRST9c9
6g?@e1U<Pii01fgf>oc<Gd=?Z_6]bj22^9CM=PmB1U?[9P5IjLUW:X>mSbD[TRT3
6X0DU5__KlJ8S1XRQ8><Qd=oeEN]6c2J^oCM=POaQ:R[pON^QYBb10K[J0kZfn>8
b:QX4>Ee9mC@9<[Lo\j5OA295PV^VXgFc?6_d3_LNhGcW`PDjWld3U]f3Lm_X^>R
=nWEY2Eej@Y6^\R5oZF;G93G5e;K8H5iK4mT8Y:`FEAR5OeP>kl=eUM[ckmY7^KQ
:nWEYmX8_B0pG?]5d^eBVHXlS[PeRa?X8DAZZ;a3N=l;]hLSR[YG<3PMgQK\hl<_
B85kTIaVU<4B\l[DLW2VX2LQ@^cDQZk]aB[6=1Il[?NnnMh2<[Jg=OLnnB\fB\VE
jI99fj8@`LKJ=l5SLm_gf29:@aY=QZk]50<g28qX41GAlUc8QddIVKQ5\=7H10da
Wm4GK>Ok1nZ6C0YodCBS3]^325R^6D<oHFPLHZLQ@VSYKZqf5?]S69nd_]jV>H1B
\46o_m>8hXXajOLS`gR6UP=j4OL0W^H=0E`VL8I1Kkk`:XTHTAe>jUaSOBfEIU9G
8<dgEdiBhKVn5iPN32<IJO@bR2S1abTaHo9TNB9?Fk2?L6BfNb:jjYFS=]M^IG1G
\\dgEdi[:U>blqeSjN0NUV2]=\>O]kBi;_nT3h]I=i17]nLi^T`VCH<>AMKiMB[?
5TE:Ffb3A8mDYSl>ob9`CJ0@chXkRiSi8AHgZC>IO7J=66>4QLbLFFX`W31WDnlY
0o=cnUTBN?nE>GehHFd`c[0G6HMk:NSLQgHgZCGMk7]Bq7<hoD4Hb;SFgZlWoJO_
:ZYh0UeCkk]^?oeOJh@?Zn7GB`2m6oVJNSlE`Ai`3Dj_V=4EALhhHR^\_Wij1`gd
;k9`e6eBk:;lJJ3W95R0bCWGmg;^[hca]SK>^>0NHl5ZL7fJh9hnbRgFGOi86`83
Ok9`e`CX]4BqVUnlBTVQ4`?A=9o^QF;^`MZcheK[p3>IPnibVSl3j:ZEl37@SBO5
]n:8^jXN4UV46W`ABdYkl091`;WRV=<P4gBn:M1heR@eaGmU=Cf4CUW2o[=iBj]:
g=:YOafXg;PC8Q6^>[[E=Yj0TQ3ejQ8fX:@KWQgPE3;RoWmRNC^3]OW<4[76Mj]:
gRmVMQNqb^\ZS^J[]3l?=`cdEAhU]ZN<8cfNR;5T0`K2`9Za2M[J1EU:0JjVZU7;
KOdW:82_GBQ<`EFhneeM28fELE`aPDhSaclcR5BPYR>m@5n8P18fOH\1BAY]F6]P
;:`0PbWYb0`\VEE<nI>?8826LXkRPDhSUX3Zc`q000;U^0?Fj`0Io<Eo4V9EO7>Y
RlH:92B<cLc_86ad\4dIcBB5Zl^9MI5ThD9OHjdjLFVP>R76__4ajfFX4];B`6Ch
RlKMH6F<TaJ7Y9SB?kWf4fP_U]O6>G[H[cm^CDe0AkF`>mM6O7o[jGBXI2^B`6CR
9_2GQq`RlimHkbSj81EhTYJ_?M0=]1[A;6KYKGUdQ]BmEV\8RdYgj<ZMEK_lkin>
8@WTLd:[a]PN=eTNOg1?0iV_2NHB=]YSMCPBqN23c<BM9=U_5_Ii\:_hD^hbPn>g
J@ohmCcJlloAmEJ]D6]m@5WIjD?F^bdf[2lQ\1T;n6l^h;?FA8ToOE3j[HJn[W>;
>a8AOO<=0RfW:^HlEJ?;RhW^F@^=K\U44Cm^2N^UQLlD^;?_OKT7WE3:[HJn[Sb]
k9DpDH;G?_ji3O[UX11V`H_QYdAQ9?KiOak<d[GkhoXd1i7nacF;<ihEJKOY_[Z:
BVgSNFCV4T@>FVm2V47dfi1T7dSn[?9m3H=@8Nh4QVo3^X<V77]=6HC941T_P9C\
ilnIDdZB3TkCF?[d=4mVfi<F7dSnH8l<`epNmmX6PeO]?mmfUlAd`TLXM0K6Qm`k
AC3K9E@A8;KF3Q:nIA3Y=[CC6e^4B<_5c1]:ig\29LAnRLUO@BW19n5[fPefQU:W
mLWK5N9G<CY^n:OH?jZjeNOGBnD1^W2BZWNNT1eN9_TnMAd:@eD198C[fPeBSX2W
mpSaA<mm@A@MVB6<A6glg;gQ;DS^jegTO<_b71Jn3USa4Y@d[G>N[4DA_XdJiGcF
e2?U;ga0A[3Q6<XM8A7W9;[YCK@^[WadnFZB6@9Sa2dF6Gh2IK\N?H08FWgcZ4Ai
oLSRPQk0=?3mVc0M<n7W;5[YCK:In8Mmp^3CO7VfgQdcg0GM\V4A=m9Kjhbk9Qe6
_`C0i4MX5Ee`Y]loF1m]c88Jn7j6;\MDn6JH`3P=LVEAiLmCMDlmToYI[5bDA;7T
bc5U88;7\@iNQ6=NMPdU=E1E16P0jA=hG^ag`EPC1Vmb^@mK_Dl^ToYI[Z`bk7Eq
2W03k]bXdXaPQAkiZW?;4J[BgFDCY:=Z[?;jGAocpB[R@Hg0;?0mc@_UCjWDWTUf
hQ1cjMDcDO7;cNEjmQ8]1F;2Y>CUV4O\OEnR:Ri5V=>X`1W><jYc?a1P[><QeORb
R=1h_D3:Y]Vo4eQAKV93MXYgcO=o^KV5eL<fDWm_MBL;J5Wd6jimJU1Ll><9fORb
R@U4BG0qc0NAblUGH03la`XH3WL7LbF;^C7o;@YddYMS@aGg`hR53?;m2N1X^HPP
4`5IYnXaG\D@c:PK8RC9AA_;ZYk@Ci@]QCBRdG:7OI\D5iHHA<@6VSEF9Z4WV^dJ
W\ThDEb=cmjOQ:Dh8SESUA:AZYM7Ci@]Ad8\V=q]P<k^Sca>Th_fP2k<9\Mm`>@E
FLl8EHl;@Si5GdNAZOYJP^jVm0H4@kSbZeBaZFb11\X8:BSPga@a6dV_^m`INb<A
FW6?]gJ:nXgPC2nlmhHP_jLEU@OZoVb<[@Q25=5]CMkl:2[PghJl6fj_^SjINb<_
bg9?lpF_CKaM2g?@=cM3R8Difkn4\bbT8ioi=I]JMZm6E\IdZc4N6KAX9?MChA6_
4_KDjV<o_`1FGEVX3P75W@7@0j]G@N^Ta1X^YSXKBS1MVh8YBVJ834[V4AT;@<CT
B<Z08hFXM`dFhPV^==956R7@Hi]G@NVMTl4JpClS<Nn`9[MA6k2b;OP5W5bi]mlV
Ie28W_Chm9K<9eS>Ek0Yke1W];32]7`B5[MhEdAP@ed7n7]Bg6ZH2gWHIUlYkU0C
]icq715hZ4SAFTSQ^F6>nN8k?\D;APUnlhPF]lMJT@6kogOL<HVQ6]oSYcdB5_To
af?2k5Ea]kOFm=S3CR;FK=]e;0XUdPHJle0?H?3?n3\OQ;hI_lGbQEAcFAc9Hh^3
eT6E7gUf3kcbm>Sg8R_OK=`V;0XU6nnD@Rp3<7O>Y_CkR^lR=FM5?^O:8YAaGTN3
WMn^j=MiG3[bdIl1cjG=5hP4o;eXia4eoFm^d[G=l:j=W?XZC\RCIV8o3hDjG4K4
iZA@<Q[UcIJTS2``O50Ro?LBE^\]lTQIAD?393c^l[Y=5__LC1SCJeAo3hDJiX3n
<p0aQ:=@oFFKfB:62QHb`;]8PRT0[gi]FhQnjhR48\\Sk@_^hUgNWVZLd_^1_AUm
X9hf[ER6_aX;X`D@bJJn7QOH8;S009AO>2ni2NJ;a0g:0j0>`YX7^nhMR_c2c=gJ
:n0SV[36;XXOf2J@d1J7eMOH8;LUok^kqeA39S>RSdSI=@K\hXVE]:b?6cmQ:jQh
@kKJE_4d]I4Dl:G>T^3X@MRR5\AGiickb8UN?_Z[WiaQ;i<G7@M^kaoXS3ma7E?I
S[ENJ<SDK8Ma6>kdBG3BX063^6DJ^YNnbeKoi]ZI6i[\HT<bl@AiQaoXSN44`Rmq
4LkN?OEe`8gS`AG@7F9Jl5DTGjcGV?7lZ8P`Ca=g6S^OWdSm9H@nGhqOS=6C2Tj<
?N\SkMWUbZ;haD7Aj`_`U:ne535KJ4JZDS64ITNk^H_kofMCT>W^M=ijWH6bH_UI
_Xo<S@l1ENC[hX]LjOlIln_ak4ZYH@6L?_A_H<lW3PLeHCN6\C5Pn>;O;4nBHFnI
ONNAS611c2n[hX]N]li;MqmSokVV3TZ8ciP=\da8NQLdm1aNbMndGcWRfPi3N]mV
Jh@\C>bCH0n:eIW9_4IfK?AeYol0liJi2;AFB\8d^68DS1fNT1lK2kf8E[9Tn=gb
6Aa0B]RjH[DBdNJS6<^h<=mBCTG0h_Jcc9mFJM8[EY8DS1IW\0]8peWU2=6WZGe_
Kg6:YV>Yd7nJlea`>Ko?QI]KWNEi2Wcj?WifTE?_J<^XN13d4Il\Vl@B`?dgoFQi
kiJPH7AmMC^UHba<>Ih3VXjnJn>72blj0E7_6l\RMAREaFab3b`4beZg@jdQEFd_
KMJmR7[SQC^UH5HlMK9qg409FlM=OH@=J[:VBF62bb[[6JA5]Yap4M>iF4F=egZJ
CeS=MCd\_n9MKZj7X^S28=U\ZY4_I>QfTROnEen<=:`TegQ_UCjVSS0Neoe1dH5E
G<SGdPkjOAXDOZj\63BK3X26I@e@NNiE;1C\cajlMdi5T8ZE1l2g4Gn6]o3=dbZ\
X<4Gd;3^OAXDf=Mfohp9:VI:BW_`IQneo>gHc_<_BCPIoGkEk4mF]ZNWZhMFTBRQ
Yinn_jlhFiLBD=6<>@RAdgV>;i?HF?C4mO8YTY>1MBFaol_dl7eUK<=Lm9X^NT4o
FAB9k[BPY`n\@keTFlK9VCU];<DH2mKYmMFYWe?1MBFRCO1oXpT>m`JWAD>4hZ7f
Zg\6@0QE<N]Ln\3oEGD32nh1a^hIPl2=YB`0ndFLmDoTo]@k^6S]lchA[nRc^MXW
1cRXDi1PBM`^14@Rq@;hiL=RJ17iDI?4F`?WEnSVZJSFn07CHDkN=3NHTMoN]ITR
RZm;UIQdc0N39AX<b6cD`CS4oE7\3^GmfVWXMSFe<PSF[h>\?0T1NKj4TG^6B<JE
WllPDXM0>LM9_mZ=_@T00kS25E5iKRGF@VW3=SFe<9ROB<Xp1Z_b9k?\C^2a8iLU
Y\6^_[FL113[;_oldAg^aNL6PX2Q3oIooVl7ibZ9cFTUG9fZ;O3k98:LlRD9khmE
TmPbEBgb711ZQBJk1UOVVB^RH:c;oGl=Vi_J8Be^7YZ]:kO714<En8I4lh99Hh=b
Tm;>EBgb\[`=BOq]MKnEY>P0^HUgK?cc?dO6Ec8p1ZZdG^8[SNmAI=G=FSAFD7f2
Cl`_DW9ec5ToVNgaA0i4FnS?kX4lVif<?9@L<]P1R3iNVNUO@5@oQ0?9O0gEVmOd
ll=hP37hJ:ZcK`R=F[82eX8n>IbEPSjhli`hiEB91lFCbNAL@im7o0CQO0Z7VmOd
5ZEFDJq[L7dg@:4gnL^bX[9>HhcCOd[^PB6_fDd[EcDihhm@_`k\Ii>WdaRPI8:O
iV:BV[0VYD0XcQScC`E?J[LMQRRMRWNIPB6IZ>j>KHkNJCVW<`hoiAj73MAmG]Gj
Md60FfT[el1DcYFc^Z68JE2MQ?TMRWNcEiFG:poXPgNU2:NoaXfJoJT;;kENK84D
Ug>lPaWT[f]0;Uho\OMN[;kf]W6S3_]8WY9h>1Jmnd<X<8=BAec=]oloLMaRPGID
EVG?K@QnfH@59N=>:hB>MXcRNR3T>`lI@R<__dogC3RXJL=^aX0=nmlo8MaRPG`Q
eM_KqjZEl?DWm]CNSO29L3jP4ofH:47eICO;K7f;koPa<0dL:h^i>a6XM@VT=Gjm
j66?ZEPR7\aNd;2c?:P0bj4MC2]7a17GSa?kB\dn6>97e3ij5079XDSI4Ho2Jl5f
ER`V_jcTONai\;lN[bP@[j4I72]7aD^:WJZp7MIlR@L]WV071Dg2FP4[PlPFELfG
_@iEH04?E^B;F7FMU^g652iYnjFjNFFm<VH@b7QD?FVOOPYl]ZcO?<T65]HMPLCG
bHjHkLWTKk6@FZ4R7X1hc6f1T<AiIgLHHV8:72k0mF98OS04_ZW0?<_E5]HMb5jT
;5q]Y1bQmlgNM@MNIFT^=DdcKfnnCLNYHE6hh1@4gGF\KJjW1OUkaY^3FRH44]C_
bJfM<h@OLjh;oO4EUV<[^jL^hUXcCBHHKYW[SHjj<99DUOR1b4N82Yj`0EN<Kek@
\Ul]9;bXLYE;C@E;UN_[^3L^hUX]IGd>iqh=SMNB[FK2STaagQ\oI;R><T@@hXLc
8UFb<;CCBT[IUn9jkJoohfKj2HIe5;UTcLh;6pT`9oZgN38Yi_>nbgg00f<\^R@d
7lX=amRG5[7_\BI1DnQIS5I<IC`VH4i6>G]gGY1TWU0dQ<4i\40^_T^@ood\nK5d
G2F<5IoAMTelkh;ZFhco4:E<UOcc<mkfGoIO\;T;8kWdGY41cff^4e^@jYd\nKll
G;hAp`h5cUS:5IjQ88]D]9?@lRS4^e8ca^=7]A?Jgcg[ZJc]oS`jhmcbU:]lFEHS
N9Um3=T7A:?V@f[7>JBPcENj9OF]\aHjQZTpP2g5k6gX:GeAdV^e`9d_<kJDC>\H
o=RWh@4AahZW@JLobZSeP\P7oJ_SFP<RF0>hNS?KB2C;EL2g@m8j498eIdY1F>^D
UPLNjE8Xl409dPW9?nh2@QV@2T]R<3:a9NjdPFne32=GEo:INmBE4>VKIdY17nH>
UJq9[Ec[k]a6cP\F;EC:SCDEckkd1^H?EN?ILR]jkR`Wj6XHM;JIQAOmG_9<FYmI
EK`=TXMnU5\YAh>>GfMK=lC4c<@L1K_]6eUS^YV`32kLIBT8[e1Ch\[K_g1_e2jP
d`?91\3UUYYYoP9DGnMK>BC4c<@aQdRS2qDGD6HL[j2W9l[eUR1>\VO@gY_R[V=<
mA5L51ij2C`:9MD4UJIgX86BZFV08eLA67^cCQPULd=SifH]4c6eVQG\]EkR7GEO
Q<Tn40`>>DSiUYW<\U^gFk217K``oi>okADeWSFUCn=C><I]3n6?c;G\]E?lKbTB
pn@EB1^BfV4P=bb`X0S?>mDNUi\`fe@ebRS_Vh:39U:@00ehTc>A]\`3gHb=ldLG
HZjnlbN7;1[0W7FFI98:1GC<gH\`iC6\:4]O_7@5j>:Q`jD`b<>1J4PDejF<Bbm_
:n\>^VNSF18PoEFcR9P7WGC<g9ZcZWIq2YB[0?Q=ke4U1^OdEh;63kcGTWh55^XU
]Ib=k8U79Y2VS:jj89mP<8HYVdgN5EY32Ui8QVTFQ;>ePmH=Y4>]@G?9KW1Xo[@S
9GhKZoUC?42]m]Pa0mo<:jR2ncaTW]_`2<4k<V6FQh7Vhm40YAm^@G?9XO8mLHp6
7WXKNj1b::F_3fAB2R_baZN`ol_573AgKQ^QkK:Di5fmXjo8Ib_7?;ko?_5Vn1]b
9[VH8h`IKb:m>;@Fjb0M8DoHo^;6oUn<O_;3FlEoI5l6HmEN58k`bJeAhVDlE6I6
cS1f8j>IG:7]>B6FW0GM8Do?4ZW91pK;5mWmLW9S4lf6P4cSFY5Kb0eb32YI>T@9
^V3^0o1ZnfS:d[ckjfE4=a8Bdh@;[>eND`6TR<lX@g^hAKSS@difgihb32XPM8k2
i1kdh\f6JGQT>VSFL==>9EN[Sj?@X6Kc`VMTi;lg4o?h9KSnDgifgi7Z>jC]qN5o
VKcg7XeN6gjjI^=dMMPIL2Xdd4::\IW33]Q:CVaSQLk_GmFJe2Yhq42@PBDL;2OV
iGG1YJAnW6b]YdZJ:EYF^aUPa_IjKOG1W_;AR1LaomL6IDkZ^AlJ66A6]=c5OMJ`
_KR]QgOS:LV[8UQ[P572mc]>gWIQ]=2WKeEPJV6INZG0nALIK\hA^lA5I=DS5dJ2
nKCYZgOS:ckU3UBpWBkkG<0B=U3W@O::WcGYaQXaaB2Q4UAL34\A;8lN>o8LVU2e
<:dU81SjL:L>M:Gb8Ua9:nX^gLiimljeINcD5M:bKB?YnPH0L_iKnfjPbfCURdaV
en`W>8F_TNRP?\?8WS2:6n2:gi3NclgeI_LL5M:bok7Qe`plY6j2UR0d=XSW5[?[
kV^fCL8?W]Rigg\Y1AQ4EmZSo]fYWmTG]<Hi\SmeJc9D>6TNa<c\D]mF;>3cRN;?
\Wi`7Z?PJD0;8qe>cI2ODoWY@=keT]?;UfK<F^1RM8^6Na>AK0:O?GJ9;1`Z3JqU
8ID0[=@OaPd]GS<956<5oCgWPi5Nf9oQ28_l97a;lLEeaC]ZNK5<J0Y<g@I0QHQe
DHXGI<WnnQm[`V1i6F320dJJP?hTiaEaDK\@3RXKnAf:@VG0Jo83da<?NCUPZbTU
Sg2UIUdnWPeU`75i6J^20dJL<8nV1qDWhiAIa<UD^lCgQ\kjHlaPn5kWl`;hfRQ9
_7e>hLi:cjC>3L_;l9NJdgAmo4=1on31DXHmm1b6<GZNF4gCo0>?gnLWRMa4E@Jk
S9>>AP3P_4_5K<W9?6k>Cd3fcn5k]gD9XAcm89bL^?1NB?gCk1>?gnY@g`6MqAaI
TJb^[nN=NfiRX0MfG[0gclflH3@33MY7ZHd=0Q@_3HMnQHS`k5W=ETY]BgnEF=Lk
4lh719fY2Blc37:TmV]f3WflgGnl3J@29nWaaKlK\JC=1<SMWjOBRhjg6[6bZA^V
DUh:f9SDUHlfh7:g7V]f3>K]U6?p]Y>Xl[b_FcRZmUCieRP1o88H^7cU>Lc9Y5Ig
I7>ALkLNiO;UPbg;8dolaZA]J_0UN8^62_kl6AJ^F[PRLX\Ym9edS7OMOJaNnkkA
M97iH>2S^G2SF2E`\m><:XYRWT:j]=^Z0_eG6m[G5[XhLX]<m9ed4SN\8<q8Sa57
ZjkjPfaALdm5j\O`e1ncHe=_lPi_\K;39eCeL09bSV;QXWOnc0[lojV?C>IfcNOh
feZoZ^YiT2PFjiMF4^nSHa`Rea@e7bI0l9^S`?F?;U@hNg@mk7L_C_aS87T8PEN\
fS<o1fmMT8nFjV\F4^n8D57edq>9>AB7OE[m:@W\8?TZ=nnof[_5d20[<BX[`del
_U<RB30M@;3QB]GW7YDLPF9m:>>R490HKm;=51:TobNM_Q>cebd5Kb[lL4hmZUN_
9<KJ_ndWIETMNU:mD3YGE<G2\Q>cim]H_c;F:b6TMANMV^>cebRW4^ieq99hFSYE
S30BYdXPD@\cRRK?AMmT:MHAX^@g]lDdefCZ9U<EFCg6Z6\cXaIZ]iJOR<RefHdO
D0O:R_gd2BT2[b=>gIm7XALX5GF7K@Cd6>FK0WQFf]\]7QaFch_OAL_dJ99IdGd2
D0<BRIgjjBTV=b=>g<iL9lWpl3?SQm`aYSG]_:[F?EN_FGZUgI<\7MTib>>dGZmb
GYTe^PmT::jKE4U`Afl[LKK7Cmh@j5]Z21Y:6FoUW@]6CgBS4ISioWPKgddc61OJ
:l_<5bG89OcVeGHjC;0M;njel>AUR5QF2bGIcF4QW@KYCgBS\nO\67q>6M3dUEKh
@`9_3bZRGB\XIkcEMU?Dh1^V`m6aP]<i9;lNFoN@eQEC1\gYW`TX8nQO1f:KJK1W
V5:ki:j73MAm:n\6Md60FfT[eg1DcYFc^Z68JE2MQRRM3CnfPB6IZ>j>KRFNJCVW
<eSoiAj73TGm:n\T;5efWpT;1U3NLFAl[1O\NZHjZUgE;J9X@ND>PUa:F7VG;qOd
876iIM<J^Z`o>HT[D\g1\4EDIdXc`bf[G8fZcY>IF=3GABX:>5M=<SMVU:QfZJX5
bH6kL;lMRgG[DYMSgC8DBW`d=4=cq?41ILBqaZBFhLK$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA22P(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
b[h[ASQV5DT^<E2:EI;9a=1ghWIWReYf<M;V7IViRk=@iIBc<mf;CZJ9no=p:Hn:
RR=hG=hQMB04K`RNOP=LPgSJkFN\VWSYH?>0T5hXS]45\9ki8TR`<6fR>8ap@`?^
b3ShP@eR\]AG?O8`]G46885Z;`@c3iYkjDMLpdZ:Ib?p\Y]FgR]QE<C4b>jbAG=A
XckSC>>56_odA=q5`BX]TUdkemf<Wo<mLOTVQFdaM\bPidE\Yq4E0nE:n8kAAN\6
SN>CV;B;VY;GR6^S3J:1p\4KFJQOF6=QYYbH]E5efU:9JdgqO4MXn65qTI9Zd^q_
AbY>HaQVgRf^@]^H2F66VbqI[8i3n3G\WB7;WCkac>YOMi0?H[o_JDkJKPiH@IJl
o]c\@1b=OfMFBZ;m>b9YNckINkY7\j?^h[aWB@0_D?8;IYkdHkJ3lk9TK[b6]=Qo
QkfEB]0QoG>4Up2AIi>;E6Rhlm3C9D0:n=TM6o@a1RfN\Ok1Gh>8?3DePio<@WDe
BI5X>0^XDN6FCW21lmJ>AB=0a05ND[SC]X@FjJigb_okic?1_Oj>RX5OQmVJ4T82
;eD9qC=BgTX^N4@HGUJ4B@QR3ma5J<7oVCMjaM2BPODWWOQ?J>7X_KB=bBcH^1lX
n=ge^C@I[0Z;Ug:NiF@6nX9<`O`Z07WLWFGNmi2@P0<^^A>;GUFfhjhmI1RqHQYm
g?=H;KERbdQ5]`;`K`X3hD7^iCK_5R<85B51TCDMUJCc>J=o]L=DY?]4aBM3H7gf
4k13NaY[716^E?k28Rqb9\89RXoOGaOLB__cG6VZL0cmf]H^XDlK4BY33ZBZh4V5
WC@CZBEZ^LHPOJRhLjgb0m7l@j1^Y`WY90BXSV>?[U<YT<^T<<?P4;P\nbe^KEAc
FIPi\@2`LpGcV@L_LoX5`:Rno_4JMa6Q8kP43B55K[KKAoDn>hdV`DTIHT61UQIE
`XGcCDRG=kG73PUF03342;T`fl0h=Gj5b=NQg>T>8oIK]Vabj_Q8bgZN]V`fcXTB
qWejBlC<Ri4`JN^n^YW;9TW0\71nKK8=D<6eaCo`phY:JgA]Vadg4eD\=oXg?6gP
RS=XLBC<:mK@8d6SCc8:CiF5X99o26<1F77UG]aYdh6KVb:QC?R9GgA`U74=Xo\:
68NTKio2D<K^8m;J>:^3n:WCGhf26Rkq^:PY:FjWlo1gh]1nC\dYdkB8glZQKC`E
S^i469EGL3fmgCe\902\J:20lQ`VilT;^W32[;:HRnXU;4O`<iZcR4q2:V:@`gK4
130_NJ7T0nhaMfGM3<>^V^jAAWGhC3FY7=RZ^APJH=6[cL]>E7G4cZJmQHWoW2Qi
BN5H27<6X92dEMljlgVj=GE246dMCG]Kb\g?YW`:YK7hR<jZ[pLVH[`An;HA\N[h
ES4bU_FcGhFTB5K<\m7TW@8=mm2HbP_FcNdj>D]>Me<fK`glf^LUhS^aJm[283NO
Q>=^;DU\2UbfG7EaAMn9YPF==5g;HMlXoHLkbLG1CDe6pLeH^kQd\PlnDmFK;0U:
^0GC\`hcXBkqZILEgNOa0mLBALB^F1dgd]Bc;R:eT^^Lda;cblBJJ7NSK1K\A=La
WM5]JDg3\Sj@@ed0e?ZA_6_97S1O_b:WBK[GFP83omBfX>_6TlU=lfEKmCcbRCiV
RkD>gOq3MI`kiZ[9MU8C;HQMH_DG\SnKdbWn[fgK^J;=IhCZ47SFK6gXHIH<=QJH
@5\LDLi[ag`1ZkXn=2`WNR:GIbM=C;B0Qpok5I:6a8lc\NnoN0bR0_m0TlVAm\Id
`7K\V@]E7]K>mdN<a5l4;ZA[\]K0eOMKPM1U?TE=MCJ16kQ?Hg`Xmc2^lR9eA=_[
Z?LG6n4E<K<WO=>DHY4AA6f9iXjDq@kCaE[5OAhdKDK2>Yc7\4Z>PD2IG>^AC<[1
?AKq<oNYCD@VJ1_mMN22=f2K4<BQSjELFYm?n\hd\>j@MVE6J]cF;<glX^WeIdfl
Ja20HOVRgR2;JMX?Cl8JkLi[MIK\KSLE=@<ZTHfo3>d7k4?So7Dk>^n6eldWb9p`
W;<kaIgib3BXjd;g0QnE;6??_Tm61FG9[<_SnAIUPdCN]g42CLOUZjXo:2k73\>2
Q9QFU4n8I0DHSmT68;]5c==GS2dElk`5@K?8nLSCc\H>\E]]7Re;D<29Cq;LcH:>
T<Y^[8J5KjoSQY3AUgDLa87aH[jhnNn4l`_5CX2TCbfG0VLBnUjYUm\\^l2bMHkE
8Aef7jU9NGIWPdc=7@i<p`7mgnJpE7@[X5m$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA22S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
X3eD8SQ:5DT^<2DR?8c83R^KRI5Z0iEKAj`;NC5gi?=82[mW8C_`QTGD8I=\@cW9
LJhAJeSnBgp6IK_La<nVe_2nZYXFTlGR\0ERiiEAJ^AnWIlA9Af8^iY<fE[`W24o
F`5o4O`lf\=D6I1;dp]GTJ_nR;X=PnW<6a`RF1VGiUhlod9mUOJjcmXoVQHcDab1
9^q96@IdlqZ`CETPfW_Q=Xk_SfVehS_6o;8a:OdO;U43q2d9]1Y?4FPN`@UoV=j8
\LKdQ1WS>8>FmJjq0T9=BOhBm>O;VFFN7bNeQ`d^El9M`kpB?QJE;PGiDg?0[=5M
7WOgl99cYL0NV<[Vcpe?5f9mhFN:;?Pd6GfL9kA?<1\cp1>iH;9QpO=WPZJqf6L6
jmW=@S6TFB6=PJh3lY8[fAgc\C`RdT0H4FoC2V=kN\S<0SHVe9\TM`eXL[Kjf=\e
;^I0__=Noa9a2R`O?YZ>UAFLmc5BLTVf\;6R@Q@D6IbC8bSFDlqo2Qf==V1cf27G
CFHHTeJVLG^6jI3cV]]oK8ZDM:^dP?9X=RiT8N_<LlcX6X;ehmkoX[e5Y[HA0RPT
^NH1n`i`Y9jKM?nVOC@HK]k<DflecD@@4D>9N6K@VpR8S@0dNQP1BbKZ]GqD>T=W
NP[2=Z_7T93TZk<h:[TS;d5=DVda>PF<V6K8NinY?DB6GMjHf\CBCn2DhUNDiGok
5M<4Z3Qo6[>cIIS=c<;QYWF]H7=X>@PG[ROFQ\94:1[dIAG3gpM1l;cJK8]o24FX
<j<UZ^93@Me>5L2@:GD6Fbh6o^OT6;=Bn\8014SUV2h_;>8[;6MQnIaHd;15m8Sn
O_ZF0Ok8p4f_F7W:@[0A3<iFRZa8jPkg2W]4YG0i=GmObDkcAQKO0U7ek`eJ`X=b
3E\[P8lXe4mk_Eb2HmX50O5InZ[i=\13e?\oGdco8mmHM<?h;LXdZm`AVjUYd]1q
KKO0FCSQbNVK?UdRicCe[?pD=2lMP[^oblRXOFNkk`NfJOT3o6R\CdD?i5E=];2_
AdVje_k:FhCdW@WccE>EcoeD\ITnl=D^DAaN@5Dej2MQ9FTBK194cI_niZCRT;bT
j04JNnimULQ9mp6J\2??\:6YVF783miAL?OfBlW]ORPUf>Od`TcDWgD99i@O:WOj
o@ABEhlk@>QWTN6JcD\Wd:^fOdL\\hFCAGg[_SBah_7>kfCdZH`[9OUf;h@FbX;O
11eIpH49OH>_A]`eX^BM]c_lCWm[SJRWG7[]eP]j;7WQQ3JA\JQ=>ELne5c=a3IA
R9@:3Hf8VBfa]_ddI\63::oVL=Iq3aRN4GkL3977fNJjfGQY1o\YXHa2iZPCMB3b
[Fk?5af_C;4`_TOa:?a:^<J93RdNhB`jD^N1MJ_RY70S4RL_=J^9W6k6Ah;f1QHS
CFO7gH]Ql_[<Rn?Z9K[l62q=_?7MHe<jcbVb9UZ3JkYo;EBZ6`_I\iPh4^ZEjCM;
k3^3FdGi?YkgMZg22ORmNTj1;Znjg8CMAnRm2fC35GWA5FRhW?ZJ]c;5eM7Dj6M5
]^cX0Jjj4\fgnch1Kp`[HeBki[n\^TSmJD>^d;SPoUhMZNb<]>fCRK44<Y[C2XGh
2o>laj\RI2AWK?VRKhhAkH@XeCc51cb^SlYV:<4M>lmlBL?kb=Z7i9C4PYPX6YmX
HJg`X`nj;BmPpF2_nLSSK@^170e@Mm=NDk4`N8?BSW2LUebVoUFbo\H<KW=2UJ[A
dmYgjXNdN5R=6]Hm^5\bA3D1chkc^bKnO]\cV<`pSB;KXGDWZfU?KJm8ilPGJOQ<
8hSAlF=GC5V\7Rf7jR82_eXGJ9E`mBd9AX;9bhd0X9]5C\B]679jcRSXPQCMcai[
<;f\SdPAbdMW0R[f^T\VHQMU<;mo5K7AC6p2aSeBhb^OnUJ@4d:Iho^9Ph4Bo:@Z
0M4IaSjh7YJ:HV:0SXWk^o<?aC4<_Wo4N8Ri\G1am66nP>Rfd;=E3hG\;eboeO2b
]:QcAmMd7d;[B0n;MboIQY7?8ERo1q3kjGF2kha[73h7lqAg5K5;PNOCkhYJAQF3
cV3T<8dD\3k^O5J9GBB9Pomloe=@\:EmH6>?2m3H;M5JEEMl_<F<K@j8X@9e0:X=
SUSlT?]JM5MBmnM2Aac9WONEUDl5C3@kKgi=10OhqC@A_lY=kR=NA7:8EIe\n:>m
P1n>VJ3kJK`4RbIYLOi34WG2@\>?R4Vi2E8;22h0@7ia8TQ\3Z[WX]XK0KR_g`F0
ihmq50bAk9p3JlYV7W$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OA22T(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
XZVNBSQV5DT^<NVXj93YglT:\9<q\=Sg3l>dSiLJ5VgRWB<@0KZaN@_iWHobc8=M
m=fS@HW<_IkMeG\kkEhhc04K>O:GEFA8@kBqoLb`N^b4c=oe@@^2P@BA9=bm45I<
Y7NgS5jEI;mnL2XMVc^P2i39D:VD6Y:;C1Fiq=bLh[GqFIV]F=2CfJdR2hSb=k6`
0YGZ@2GhVV8P1mp>24dOM@_X\@DVmMh4bVRb:H>lCUQ]h<Vf3pJNL0`5=VWNge`Q
XWiZL;6JUIV]Ao<1`mCmq2\BZ>Zf_7_ha\lSn1A`I]MAPADpgHLo7E^Igee6O>>C
3CWQ3XSWSJqo]VE0aCpBhbRaVq^3=S`]=<EmcXNULZhD6]>?^:A=K<IJa6P@WKCR
c4:d`TNV7f\LRKPfi@@3k]CN4U^MoUa=H61Xb0CRO[XdVLW8diajS`=IXh?RC:WR
iHYekh2hAii341:cenShpE]h5``]HAQ=QbUOUIgn^Wk<XD^CgFO[Mn1XZKTQSO0[
9IZ`j56dgH\C<[FT5F@md;dOEHk5e5P40M48gAKX=@S55\THUI2GkeT0kmTWgWE^
OknbANnmP`;MSS>q4jmSA0JmPXVYC9Cm?@ELggAZ@FY0Y@9M`EE\QHM`LlHjWV`M
7BEXEEcG0hFeR:4=k9Z5Y3eWLI`eU[fUm28RADL?TlElJT_a0\o1XHAA`5_oTl^@
<CZlaPXXYVpfJAn?\mJS4Fk26kdQdS:fcRC>F6ji:KhI74MRWYHXbVF0gnGGnU:G
VZ65m`GQ;cX[7TMKeSB@bE5NWL9<`[Xm9CLa2q]gOc@4Fla=TihZD?c79GBkO_e=
4dH7J9ZJY6OUe7b9<7VJAdiIhmAD6aVE:MV9_51eMJ]DSd?\[j2C_[ao639aDKRJ
goLhVP7ebgAUg<RCXUJVoMF]L16SAGJNpJFPZnEGJo^?2\0AWOa6CG\Sgm6eYEYW
M;X1nj>f[0>k5le\`OTDTVQQMo]A[K]f<W8N5iJ[2RH<?P5TTg4DbaOiH]B=KVGo
SR1Go6>RWEdOih2d\@fZ>2`8<MBq]?D]RhG0cIT=\[Zo2k4SHah[o?kRb9R>dfRk
4iYG@8h]C>R`JfIN;Tl=PGBCKHm7k7gdJEkhJ6C>^gA9UnGgk`_kl]CTgik0^H5W
2iH:dog<5nY61`2nGP<7^hqm\nKN7;JR3CDPc_[Y858PebEM6jplh9@g]gbD_mV]
\]9\TjP0`h9kBNVTZR56ljVcQGG60F;d6G01i?^UOF9K^1^C^B;eYUfZP\DoIh]F
fiSgR<AmUKI9PpIMCZ@Xd_M;YQ\8`P:3HAoENQb2;SSJ7AYXj;lQOK1cH[hFAkH0
Sd33<2`WkCe0JoG;HV@1Z@?cllbaKMlB69c`GOK2K^^AcO\bETfQd\QjNiInRS]g
QSQI8eM>q[TM0\j1AcJ4EIdMfg64E\iYjm09Z^9;_mmk8Za5EKbb`4kZfC2IZd]j
Jl7ml23Jb\TK7j1\:lKYmG];l7QTB3L8CFDkkJ>6g<baSLaM4ZFIA1jmeK0j<kFH
[F@qMY@bH2XN6d_IECS44MHW_NZNX<A^53nk4:JYMgO05O=KfVRDki^mfEHjFocn
e65jSIGRlg^4M>8S8A=khIC?6O2db<o>D_1Wkj32MhZ9]l3`Wdgoc82O_3AK[klg
VlpXC>BF`B6K;kW4oUBW5T[g[3XNooZ^>?[Po>9Wf58^::Bo`:F8Hjdhf=eEl7c^
Lo7NlIUSGfPS;Ulhe=HoBYQP:AN7\l><lpcbSQXo>Q@b\JT1Gb[bl>>ci02hikHc
:<O]YI?]VZ_C`A7O<J]:gDa_I_OPj44OViWVAEPSFP[RA][7;Z02eAd<`aRma9E]
ZRY6k[S]4n@44R5c3kOi;SfNlmZ7qY02EC`nnEZbAn_IIQCbn;3b\F@0aM:AX8`f
U19Fj_5eNj93M6RoIkdT8^AcaRo_3WL60=?I[dX64X70jK9g?>fEciOnLYSV>RNN
=l9kDKOn6l@QAkeMZFelC=[q8@<iC2^gML6T[Io@E>CXZ8XLZU2OCMJNFH[?ekCl
2jPK9oHeaNK<L1TBGYYe5ITQSFN@ZaY@6cJXcOim`BFP7cV`d75`0PWFJOV>Bkk]
d?;mI\ei<85Fg:1Y4ipTSZM`L7m;j\>U6NGdn`:2mSgN`[0[72MQ5OPPolT54l:5
7UTmDCFCUT]c98WPcK:3849K30H]9:>fa^HF_;22SoSfoqc9D@:?KbK:C_FAUOH^
q?e[J]ApCIX5D^T$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI112H(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
KdlLlSQd5DT^<2CRk?VfF`bSf;_lBF0[mOHnf_Qeq@70;aag0`4KXMefg[GnjfH1
0DN=Hjo@;ZEW5LRH@=F2Ze2gXn\RHVLVFID\`g2p^BJRdaVC]@>Qh:LjH5V3gX5]
hTK^o>EK4heJ_79K=IO\RPbh6O@NpMgadKMp6Mf9PY2kXR7iE=^nY0`FbfU5@nk_
F[HiYdqOL:D5A2e=YSbY3]6K>GhEC@8NWoE[Ncil1><a5<q1TN1W[eqOdVZ>=qVd
o794Rbe:YCDl7PTmINeW<D<WI\LDGQiJIh5ffU>W1D]K6b9JGL3mO[cCV:ICGIVF
jl7Wg>5:2a[MlN?5II?e^hD88PV2RTkJTMbSCTS;VL;Z2QIca>a_phK[ii?=C41@
>im@8BPhWD]6YQ^^dNQJCBBBIKiBfbTUiQ0l@PYmKaXqY;_RF[b=ooH4EoSRE5BV
M=O`i0j=_gN0diJY4CKiObmhSI?JAjc<=^HbFnR5G=6nY6<:IP<dPoVjYKUPU49F
Ca[:6c]:nAf2FiTiEDT02aG\`KTSeZgAidp0T\2aLP_ALZQIUC_MO=oD?n6M^kC7
;[GoaobJT;jWhBjM7K1m8oJEj<XVfOMZ^<<0TDd<ZTU^QhVaF=`^QU=TomC[2jR6
W?EEamGkj<D6jcFMZa]FBDA5mpN:g3T`ic4nmRRRLTFJ5V_@j=Hn=N`?]0dM?8[G
Y7YAiPMG86jC>@NZKU?eTbK`YcNGc<d]RL6K[\V>6b:^bH9=qfRiTXKPKo>GZ;ZT
\Xna3Q0iAoNNEfTDLV7@B0]c>JliX\`>hO9SgYYnO8Wgh1c?]f`T3k@[FU2goIn8
5_Ni<OmMZ_5YcS5iG<7BFPMUol@I=FgaLc_@Oj1p1__^0X<65WTa5JQf0ghlNULZ
E=6hf3MM9=l??JkSOSa<o^MogaPL^h4m^glNJcQ<1FA7<:7\^X^bA2>HWmc[jTX5
P=8?DbjhX=F^ZkSE;Gc^N>5=Ve<QJmq9@YXf^`n0kMJ^5b2Bk;ALQkETOGgYJUB3
`X<I[9HiADd?nV593elkjFXD5b<9A\^922ZXl0U8BW4OV^iV5FQ1diK3O3?J0E@2
`kcR9:5MK7I@e2:b25aY`qV:2HB@LADmfohbHToil2JUF2\8M@D^;XhgO8_lf[E3
hA0PDdN6b0YMd`GZI@OVoOVKB<0O9?R4GLo1n@G:UiJ;paSa\aE<EJ@lf4iW4Zap
hAZAEcqkPXn96CW4\IXUJ;n>NF:c;QU`Y36dR_8Hf:;QYf1bIlT]Wk6Ck0BS@^MB
N78]dNKk;WC?<[0Um:XF3d4S;GpTeE3]dbe=[=N6]UNQ]LSc?_IKF5a6`SS=iTRM
c;`dhCP:d5BO1Bh3o:@ae@9[ckDTg`kH90bLjg=0h:=GP`pR6F^UUD$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI112HP(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
T_gYmSQH5DT^<h7`9AGGmCHmgCOLEUWg\9baOMMOn1XR8K8`o;g1e6qINn8YN<VD
TaMnLJ_bmX?pm]X[6lLhiRD[FP2hlE0DDGi@I9bdG<7\6@k@iDZB;[IQXB\CGNg@
qXKaZP2q4jRWKSZ\N8idNZmM=ddZ4mmj88g7_[g:4OqnN_o2@8VPAI>`BoRQh;ID
2A2jRDCgGha_UNoo]TqjnMWMKhq3UdZ\MpD]7;RmZTm90\0H[M>Jd5b]TW;^6`O8
PnZ?E`YgU>FVF9HFBA8@V25jjdOSLaI>]oDRmLV0HP>9nRRaoZcHdmgddI771:g]
5RJ?WH1?a?JCJ4<lKe:Xf\AmqSXR1kf^e2KH@ibnAY^CQ;2D=MI90A]:0Q]mf3HH
jOURQL;18qgkTh^UZZgRHQ8=8:258P5F6;n^eB37CA1D`WMOk4_fcG0RX664glZ[
CDGgXJCUf_gZOh5R_X]RY:?Li:RneFohi=R>LEE34>kD0IRQ^P9DlW?8nNDBN5@c
p[5`kb1Ph67iUUQ5WM0Y@57`Mal<>?>QFkUfEOCYEUTBSG94TMKaLO7UZDfjjYW@
Z[c<mW;;QS361c56WJQT5GOgee8O1`b<PoU>Wi[RC;i[Ca?H:akc<3jq:b=DZj4o
JD^TQ0iml6BReLYS\`3Ad@O^hYC]fG:aTWDm9]=bb7HjVQhV3TKbd`IQ:0V?A:IM
DP7iDCXDGTnGO0p8JE:8j<kSE^f9<MhVL@5fL?GVV3clPN=Oje2dmKW;PQd]E?fV
D_Lq?1J7?gU:_lUBHCFbEe2W18mC2CY153oVhI]_idg[0FnY1jl`7IFF<@4Acf_^
Dh<b?;0k8RA?077P`L5VIJleO]kcg`\KZo9aHIO_81EcY4Dgo^8gLiDGJXpWT15a
7_2bXO:==l_dQdQiPTXK?fJN1`V6[W1=gXI_HU>oH`YKm]m6C`8nB<;h>bnWe;8f
\b7`FL>4i\E5BN2FPeE>D_d\fg>[[KcSG6Eg_WXNUA;8dGjglpO1@PSgBBWfJTn5
=B6BD0LR]Ri7gfBZcSj7]:NMgITE:\jg^dCJgZ>fkESaGn\k3EO=gAjXn[NKj^19
n8GoHWcK_>DO\3J4<jC7`c9PLROQFD;@6ik@]a4aq^[b5>aCbNim3Lbi6L7odUfY
2Jo]QXK`]TIAT\VSl58;]mkZMEkPl>eGe:Ya=UTfQ^IH2Fm10R0AOfnkK>o;@>Dp
XPKR:QnE;]8R^ILb>SU0iPaMIPmo\`\`hV8a_[a4[aR7Bo34FN;K1SjF>f1CWg@D
`5MJ]SV_pFR31EhpWW24>Zc9GXA]oOc6N6IWk^Xhm]SP9@C47?L8\leG1Z\e`QSN
C1<LgT3;Q]Aogm^QWi8jf>_]1SMIG^1gaf6q6I=EMSGj^^naDmX`C71RbmI=G>>0
OfOecad_a^QOdlUJM_H]LUVjdHEj9Ef_EXUj6D<B6kJJdVT6VcgVfQDq7CajLX[q
RN5ASXh<XkA8@Ye4X`HnQ8S:>CiO2YRclbF$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI112HS(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
_\g4iSQV5DT^<E^i[giYFR:CiK?P:oC3Y3[;kPOJC[8LJficlAZidR[[VlO_JKWG
C3>q?OQYH5P3\LiSFkNUiWehVEH@0<9C05GZDcYkil=PbcOkgGGqem1Gd:3l62Te
Q`13lBRm<:Fh72VoO8Ekb6K`CULmA_;36e3^c__1LBqG;0j[Gq6P8l9>n\:]c0a]
=6Q@V?Q7j>i]\f=WolYmq;EYI=ZYT2FAjA1L=YWj>`c@:146jE[b;RJdN3]JqJBU
oei6pdPn9iBpIFEB5BV?kDKFnd8@K;WP^9N8`RNU^=gJ<jU<OElnL3eHRfCjZ2nj
Oa[?a>Cj3>HhIYcaF;A>9QNL`nch_DI9Rg]RH@Bb1@N5FjUhmgoaPo36oj2UOb_0
Y^pf:TET6K=[bCkdXj2aCq>jGBL<Xh]aJ?69HP7E\NFl<hndUCJVKT<7aAea6[EQ
IVDKG0?CN`A[GF076k0n00>_MB2laQ2NgM0gSgN=ZQTVK7]dXAHS=kc7gg_jK6oF
0gMcNI]XUjBgp9^SBii]M28<OYejZQ_0nX6>NZncZcRBY=kFKQI0203eR``cQWH]
l7Gc<O<2l>;=E9ZAAWI^H7eOI1J78UQX3D:HJ`nI;YiT2akFK5\\nP@CF@ZUnM7E
JaGp[LWA9VFnCUT?1kC291YR7]UZ^ck^gb_^h7?TPHKEm]SFQNIZcoNCGAmOO`X?
lB]Y[Jf96II;1_fMg^\JAa4\X6qkkUR6D8>j:U4Y[Um=gXI_HU><H`lKmC\K8^J5
>^WO29BJ\i`PVK:8XIGACOkQaa>kS]TcfhBOZRcWBM7W9J\ObC3OInPmdmUY8`0i
;DZYk>^NW8XH\W920qjefg:_k\[b0?AFU0EjKf;QTE2Y;53dj3G99AmT_:baNck1
<L`5EfK57DBAQG0JT0jkA^LP^3d:oY`h5a]>DnglLlc4RT:?M4?9CC^lS<KhhTN=
5MRPX7]dp3@[gPR1IH]H_``=Xkmf:H:U7P3YA]^mWYRf\5XRh3ca:;:=J\5]k0j>
9H_9kE=0l3hAn\PP`3QARe`>9I:ElaO[Dn87VDack1RQRB^gB^Cfb_>HKFZeI\cp
Q_;OFQMTaH[;;4P=gOI1?a<nT[Mahd>O\CKn13g99F04SB8H;BbQJal6CT=\n>6X
QjU2ZidaHlk7\TDQ@?U`39qbQj6LIpVVQKI]=CcFF9BX_S^G_o\ejS0RPYXO787Z
o=p]^nJ\]7955Um@0ImAfAPc[:ldZoX4@o:2MHIE<d4\T5UK;^GZEH;2Vjel];Fh
FVl]\8WNlcVFYFoc\19E6mqSdQ4jU7jZ8Q_:HOao44\=e]9l\IX`4\<37jKY4HH>
F6^SM2mGb3[>GjEReCRVDcHSc;LM^<l::9kNbaYkRBqMm\4RLT$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI112HT(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;

//Function Block
`protected
;Nk9USQH5DT^<h=`7mA6inq;4^]:ijllAST\8K;N2]\Lbo@VF8^c_G7C<KR<F>K^
h2F@H@CAeKZg`U?gbR2\DU2ELJ;p]1f[1]koR;6jhN>SUUM2in3=6dCX;bnqV]fe
i2qCgo5Sm>5H1MJZmDE2e5Ra`0Kk^L_\=[KGlpdY;^LVB^T>9P`IEIh`i;D05C<_
h`RI92Z1mA1UJp=bGaQ:IZJ64>aWg8L0c8C?o6;^i3SWm0h[GML;Xpi?gCX>epid
anY<qeX5U=Ci:Nb]2Ack;VM`PN>:9Ro[<NI\5d[VQ7jB6_0nD@P=FYLOCF:f7g7o
]<J;\ejTHCFf@RbC?\J6`l[``4g9DQMDmkX:\h[J0Qc;[A2WPK[;[;QL::hp99hF
S=c[32=Yl<=]\O[gSH]CiNT4PSNh85:J\aL=97mZUoOjk0jeTHF@EE9:Z_XG9nVk
Gdcj02lK_h?2bY_M\m;`55C=XL4[G5:g6C@7>[ioiE3cfY<191q=>e4k:^6O\nP=
o]@k6P0U==EJ?0?5[>W@9DiLEGjFl<h<AUN`V:U^NFBb[Ub4`]:=Xg<MX7\_0U4E
YW]HCo3dkM5Q79iRTS7U9@TBoCoebO2[mTRKSBF66pW\H;2]A^Lej8Z7@K_ZIY4Q
=bE9U6X1D\=YX==0neE[PfVeSc>E8HG<H3Yf\\:Xc>WQ\=XcISDLkOeS]O^8;jf2
qFhB91GG2J2B_7MVKnYBJi[`NY;7kd=JKh7P89H1F48<VXX3kbZ5cg5:5?DealgR
@F4@>\2JKHO:f^AaINeKn=MmDHEn@l92Y`7LYTJQ_=g@XL3TWm_O5BQq<m;``7>o
<h?;\5[;hEPHSTplkA14:3ZL3^4D5TgQTb]?O9S8AUga6UO:k_1Nk@D[iTOW[bAh
H;QTLc4n?U6Do29lCAkgHoeG\L::7I6B5L>ejV2Bc6jKM<aek_gY?]@M<d@[NRbT
MLF9Yp01`cbXiSMDV=R30?T^j_9XKYI\WV=dfG3CY^ViX6fMDi9b45YmhDPXcehn
L>OVe709V_hEB:oljHSj62n^e4HW`FKC3WTYMfoCKVAVb`nIA;V7616jI[=IqJ2n
T:`C4SX9YfG8?C:4T3d1fYabPZVWhmf1i0=PX;6<XhE?5FBZV8\lLlkE6Q<EfJ==
TTe4h^F74H7BM>LAS3Aq>6cL?cpYM0[fCQMdW3=aWfT[S5gj[MS_ZII:X6Sl7[;D
RnJH8VOc12>_c[3U0akY\@^@3AbYgPlIADY_g<P[=BcHl2pmOU>SY;F7n99gmG=Z
[2kFQcSFdK:CH_IB`AjB@a7H:7MekE4L1\jc4@]9UVN3o>Zmd:\QCePhdQ2keL@o
=2pC5WKaCO$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI12H(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
e2aETSQ:5DT^<<>YaAgXH4H73HgXAh0^11hp^NoDnFaB=IBAX`:U=G3nn6hOp5DR
PTOSL[m4\\FJHSQqZGRnjDq;hH0eiZhg\[gJKQ^5aa`MITE28IR0D0P<IqkPhDeI
O7j0QFZgXiBGm6AEj;AE;QO7i3pWjjDd3nC^MePP4MDfjR_?0HI6`7CEQM9^ZJ@a
<qW209U^cp\\\>CHpQ8E[DMEm^65fbXgKGeR06eRGY`6gi;3Bi3\bJ>nd>ET>MMV
HK17YFSnRY_UY`7YaQKGgRaR776FC;f=ho3Dg]];\P19538MP33@=_=[804V>hRB
==<]jV<p2nm]igT6kKA8QKSa<jL5]K:>YjO72\[Lk7\P^:nV@4=0N<0RegOb9j?Z
LhZAHoRn2KH5O2:nQfLIhDKSNO8D6VdEZZV65;D@77HOAVXdo]LG:ALCE2jLHWq6
fRTGm=<ZhQR2okNVQdod7:T_djhieDjQ2?fUVJWMoi`46U7^RZ3j16Egd=AVn8j6
F]TngQNTh<5mTKL@[dGB^g8>dmlWMXAm20DCIg3GhOdT;3NcQhZonq139H<3]Mhe
_Iag5V5dcOO\<R3GL`IQK<6[4K>=j5_BBL8c5Ll`cFAYT7gNmJ^3FO1:ZN5PIDIe
6SAA`?VG?H>ipG8KXmNqnUmXhN3X3dlC8D2MT\T1qoK@2R`P:La2?GaO8e6jIb]:
<P@=[7E7NUI3XKd1k`6_FE]QcQgG2=D2`eP7fjhU:oZT2DbMejaM<[4g9G@BpN3[
l1i<?=kBAC\Eaknm>HfDVCHR7acK9g^bGi3QjmOmnO5H?J`@K[oVNOK<J4Db=NIE
SRAANNM4@L;KE3e;q7lS?`YS$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI12HP(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
Z2FE\SQV5DT^<\fh09h^?Mj2WkM8Wil8hLJQ;9W1X\i??E4Wpn:nVonWjZHDdBg<
cW85Uh@Hj_`GW<]ChJ]ZIn2TZXA47Q<EElNq@iR8h4;Q8nK;^iLGm2q0KB>g2qGZ
YM=NDlG]OIVS^HHUUcPo5h?2FWL0O?aOp7OTN1^5N6oh:_`fi<`@:_kiJ;ON6LL_
hqUUFJGgTq_`=T2^qBB;jEDl_XbDeL]kcAD5:FI@babP998b<BFFf9KMAoEJPa<P
^^L;7EYdfhMT2b@:JBKBoLoNA\bd\FQQf=YciiJ>ebb@T`:8_JFFBkUP68Y_Njh^
Gja^Q^Vpd`[CGT10]?:<^O?1A2E7=GeGKaF6H4?JlQJGdQ8[?_35@GKXhlJ:fGb8
4Dmk8GHKdQeEb9kAm?^]IDof\aEe;\mGI4EY[82WFQNWL]Ne19Z\I`Zh<5SO;XqT
f[eH9m3TY`5P`NRhJ4`2Ube8>b=]_Gb_ijR[Ra@6fVI6YDbEe@Pf<o2nR8_HmOkT
ITCbj850Y7a:mF1;34>oWFf@>DmVI6b^i>XNEekL:U2l>oUSVAPV>pnm=B>h7KS@
VZ7j>J;4S>_A\9U4QTQAM_>J6j\YBlNg_D1DVf<J5I6;f[pYLAFNoU2YJ9l68Iib
WKKn;5lSFBDX99`UfP;A2=[@P@G\SZO4;jMEQB@8?Mb_G4[Y6l7>n[G^J`nkFGGU
6U_j=qhHZYX3p9PQ1fo^AfHUa2UPhQ<CS6V\FnH9\Ued67WAMjRdVHb=lj[GR15N
D14BHVBGkMFm59;oCG\_>VHGLaE2EQ8Aq]XE5R\OF[7QJXm7=EnJF1CMX>fT561g
K7PJ;XG1lJM[o\m6T\2AP^hW8KFB]cL1o]URaFN_GC75<8WjRl98q^HM;]E>$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI12HS(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
686C8SQH5DT^<U_HmM=Tf3RaghbX>L6o@CS>:BCfjf?KT<E60f>6Ejo4GBSbSoqS
^GmWnn6INe7VE;Z2>J>j6UPpUdEA7NE_Vb<F[MR0lgA0kaUbSWC:]3XYDH\peT=i
?6p4MYd[<Q8\8cald\Aa505dN\`=oQbHY@X0^qDUKIYh\3[[PT8aC`Zng[;@n<h2
WQfd=OqVLI:^aiq03K1N1q:RX3EaACB[aWFTR<2jV8ZVFHW:oLC3`j;ME8Tk:kS6
TOQDoJ`]b@?iZ[0MQTn\gH:0mi>bKhc[Hf5I2a]Q5ID^CG^joOHB1LoM;5E@bgZV
I;_?h_98A3`kqn9oYga`GE:Pkoa6j4;?1mN@IW=NAdG1Zp6BN<=57:Cjb73`U=Kl
0dWI@e61jfmhHKZ4aYjGTL:2m5<W[kc7Xj<3WIHF7kTKIA6O]^1gd0HFnGe3Ff@l
6nASJQ;;3jc_5oD4aSab@2_5@:gTMNdYK;CnpQGdi1<@S0bfY_;4hcYifU=2GY1l
Yen6WJ[^lR>C]Sjmo48?cdM>0W4R^SH^4EXm\QNDU4Jc83bAlM@9FfaiYT6``UnY
kR;IiR[mH\hGO6]OCVO6Rm3W<U4p7f`X7\OE0G7XBQ^:YKL9ARe;4fh_I<?W@Ulo
dOHohem@Gc?eS6\L9RW8Geol\\[o7NambLYe?G=Y;F]`4k2N<Cq`@EjfoqYR=HL_
ZVkFEfd@[Di=j[Q=jEL>oQ6]EFlI3pKn\<714]Dde0XIXZ^iR^=kVE3l[dFK;8kV
S3FAKO@iA79oe\;VX?AC6G3@]b0PRhKgg9Tc@5hdGRmm18Z8Ep\:JT;<n\3EQ_gV
=n:IFHS=EY54A60>1b?MTgC:9O@Xi3=0KQmM[f1bU6Q[R1UOkD\Qh[HAJW\lW:e@
VnC[Pq03JZhCT$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI12HT(O, A1, B1, B2);
   output O;
   input A1, B1, B2;

//Function Block
`protected
98_nRSQH5DT^<2i]=D@MN?UF[j^l1QJh6I?]j6C\KJl>\e8]RNh\SaHZjdanPSDH
O4>CiD0E_39>pc[IMhY5man4CYJQ440X`TD43YfLAPo_VoMZ28VkTW]?D:<83^ob
c@V6W37Eb3HY^N9\QNS;@panEUbMilK@6X25GQP]DmEQC60>@qh1\>^XqM^A8`gK
>>K<>MkbJ`HGIEbi1]]X;^6fcKBpeS8`TM8h\6Sk?ORM6bKjo8U39P:fUf>Pq3?Q
ORmGq[DHN[=qlG]FfcA4_8U\;WQZ2kW^I:5:0_5CZaY5ghaTR_H]1KF5?[L:68ig
No`T[i3PolGo^;?=]Vop838eMo0bi@T;l2e0CHb]\A@K?ck<n<BT<[dIh9QOfDbj
1:Xhc[3GM`jj]EPcPLJ98a@:oAO5c@8<KQo>me`>2NVAdAHX0X7CP[1:h]HD38<5
RP2?gDLFD[p;?NA_iHnE\fP[OLEh3?N^]RKl[HP5hKGJf@oY;=ia^;KgNWLnE;Wo
CmSe9`i2\Sm;Z@F^Fk`W\XAlM@]g`?glI=kRWS7f8gRYfc>N>:NijbYGVc`l[9nU
9p6M<T^WQHHPkS0TSjF6EA>^KI=mmbIAhU[PmAg]?0WBa4LEk6Io:G6nm^BAA;Jc
Yc6_iX5S`SlP>`S@U;>>E]P[E]MmhhfjjWRPU8:j:27T2;_>YFN;Z5XTqQbP4_V0
aRVRI5MT]kKQZK2RVjIbZPLdFD]K=hcm5ZFj]ZIOm0LT=W<UJ[@4[S0VSQ<:`<T0
jIVn?ZQX8WBO\n6q5lW3:6p?a8TUC=eEianG0eb4K1>;R\b0^3Q>3E2[hiVXVC:D
AhDbNU3SZ<o;^F\R[oG7l1V?UbgZ7J9Ci1`TJ=lh=9qbJZWcJ2k>@I8kCLB@3EW@
m3W>bNJIaNccVg;bcS1CMma=D55YZWZl^1d60g?VQNJbH<[=KMWn@98n0\V[cjp]
`:SoD=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI13H(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
heT1TSQH5DT^<9ERFAXY`7dIB5S15=qY2>`Z_]2m8Pf_HW<AL8COA7KL]FGGB??c
oEi2:4dbL2dV^j]h7IC6V0q^P?I^8[cc9i2JGC^q44je60pDo6G\O[>56WSUo6D1
afeW1;V\b9B9G:ecoYkn@4Lp>?m>DZ0a;>OlD\D7[noE9faeBlbdb_::p\iQB[@Z
qa?om@>qJ6[Zb8C4l:7iPF;DXRdlpcdNKagL>==UF];lE<4cb9<Qm8:8E9LS2`BZ
:c9J?l[m^?lK34\E^LAG=8j?nUjgccE]`Y[CVH=[5R[:UK>c_<a:=4A0Yj`kMeBi
]N:>O>J^CG10<L4of`=i;m=[0nhXO8AkjdmpkGY_`<2IK6:510mB5mXDEJ:HBDMm
oChn9Kj9LS@SNKj86<7=Q;1P8GU=]GHClLmVkK7fk9`<TGcU[e2\KICR60?:K7Z`
PONG1KH@Z_ok[MkXXf8O]TlF57I?DERkN15TLdE0QXqlako9PgF7oo8J>;5OF>g9
Gh7o5kkB70>l4d]@LZDRBf655^T<:ADYS4<9Waj65L=lnlLIbRHmPXnJQ`JXM=<n
jVnSVaEWeodQ4U<\]fW=KXl>9LAbfWkgK\\jXXFnDNBj`<K_[q8;chA6k8OB9?30
c9C<b97dZDW3Yl5K]Qe@h3KQ?ni=^O5BLg?:e16Pn`J[e:=4^C8A]J4UOG6BR\W4
o7hBSWlK1:C=JGM@AJW@hLd7c9cW``oF3TN=1CnSFC7:k?g6A?P=6NZSqQRDYZW`
Ma^jaDnH0@^:989KSMN[6U>EfXFCNi0OM[>RU[dPO:bJGQogiN528lnaGQj`I_UO
2n^9N>kc\:=:=Mm80Rh_n<ZD3cFDNHcUQ9M^;ga_D<5[7P11j@Sf`\6FHeEX=aDp
kZNS6Whihf\ig^KV03FPU8Ik;0=dU=<<HIAjKX]KH<P=hnMWo5^S[a<K5?>eL_IP
kRP]PoPFcfc1?IBMK4F]`4I<Kn095dMWJI;[CUW3M00;HODbBDdlnG2a4L19Dk70
\cl`HSq^N`lM:2;:T1@Q0[`DWWkBkH0Ngdi3V8[:7i1>n7iU6p0AnCg]1o_MkfJN
oLm[dJb]ecIKL9?2mf41dT@?M_fiCNDFf3d=[09b>62ML9RTH?0f?\mP3EhM`Y]5
RG6CdUWAGOjEj7Mk5;]1;lB]E@0f<oEA9<_UJHMVW:KmV\Ve7OHQigQkpEf:Wea6
SAbSl:h46>Uddc^TEDa03\>dCl04GJ`GOK2\T1Xd5of[7\FC6V4YPIEhPE`XJnBC
a:bL\N_=SSN`d?aq]QPFcTpoSf;n9EP:PSQZ6UiK3C[VB>CBX?AM`Y?>b2R:1iFE
l7cbioZa]]nF60hK?lOLe<IoGUGP;C1YP6:FI>fl96qbC7fB\iQ_9<FVn:j\1Ne\
P1YKc;=eJbjmUkUVn8A=W]=`=kaEjgg[W3I`3P^:Ae9bKGb06keRo:a:A>d:Z6q=
g3SeR[G8JeTO1oSOX=nROS36K6\h;XTo=c<<:D]7o8jhf9LSO5A0Rfo?E8eK<_W=
5_AGUWi``Jl9DjYiQHpUhDW`2M$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI13HP(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
4:oGFSQd5DT^<KGX_dnj650[Y6E][lE6a[JcIdP5SfJqCd[DgnUWd=DUM:i>RH[@
ic3eH0gBm\bJC56PfL1XUB;<a9EJq8>TI=4i]5l[e\>aM^cOqPHPYCPpeomBPjR=
H]faCQZ@6NM>O9d1M<@<hm@CSN_A4AjCqCDL;QLTEL@F2MQTBd1LOA82H2mX\0@D
LqQhE9PB3p_2SCcGp;gOZ=ea2V6EloA1S]UBcV]fRcGaKN5SBIVGal:n`cB=iZUJ
W_F=ICJmJ]\l@;LnO;_IFPH[UK6b:mQngEn]7bA=^=cPBXd62EVefgkMFU@FmJon
ln;A6KdiA?KeWCABNGAmd3_p?TQ][aG<3Ue0eCYYmDoFGV]\iXZYLTVB5@apI?<W
goI]1D]Q6F\JHKLmFA82>SC5Xh;`IA7jLJ1dO29_XEGgkSS\Ve>\3HaHj@k`IlOn
Vn7D@b\PaSGjd1l[mATXc@E16?IASA_:GVJa9;XXh\kLDUlGCRiY06Wm@SUDGR:X
7=qNVNi0Rljl7eARhl>VZK^i3e_OU`18R33AF[nBP[9Dg12Yi?3`WVP2\fE<O]=1
T8GN2Wk]\oZQGWP3lH_?7fAQaOcBURK<[BGaF[cdfJdfE6TBR_ZclNLck_S2O;_A
@W`@e??XIplD?L]dOgonHbTAIh>SIJjZaeCU1`I<]M0V;L_^S1=P]e^mo0VcY=JO
R?IXhm1JkUlg@4E:>W8nOC`EYJSC55DT9hTW?4[ZX[7V_U_Pi`B\208WTBcTeKkh
QlMhA?eN;MA:Fn6Aq9bMedCec1SZSJ9D8aXM4K=9hXPL=0Y;jCQEQnnFWemCDa92
NLF@Gg[b_AeiIlY6S9^cH;ffhWS@QKQeT_PM@oIgJ1>J6`80^gQ7[kOa@_2FT9n[
GVPc3`gG=66X5_hTg=FdI53p?8Y;9=GQj1oR<127_36ZUYU1\?PV2I13l7em^Fa^
5mg@h28`QTdI_oAAIbDVE7=Z?3@;\bCWW1\E38][kk6H=DUImYdiV@T?67amUM@U
Z^@=>S;MX\DCC@5f6fm6N[JV8hn<C8qBBTllEaQE4X30f8PT6K@14HEnm=[?P]:H
@kJQM=ng<8j6L4^b=iLEQJC>hSF7T:>BIdYIk<EA4]aXTnUo=KPioCA1YMBEl[dc
@nT\1IoeWV9\FeHGWdPDCO=WWH^fCFR^AR_5OqohFi:1K[g@@5[GUNO15LigK_K3
bIDi=RWB\5LBn[8mOU5mTA<Pl8e>IBek?m5h;9o3XiRN9YR@edFTM`JDO@aPqMD8
6bDq2L=6A?_Tb47BXiEZ]n^m;KT8\GDk=Mje19eU<JgqCM15a_HgSlIS@W7>;PV0
YEMk3]h@keIA1gS5\ge[i`C9J4[>`WOO;ohCTiC^_><lC:B4kWdD_lh[VY6ISNUp
b6iUTM82A;6<O:gV<\4Oh8GE^J:LR96Je]`ONQn=UiNXV7BWgkHTCj9W`fY0EhgZ
b3cP\_8AV8@Fc]oTULQpF3UUd?a_:aXHCa5hHE5ioo:kIN4Y2J3F54\?PkQP:OkD
Z<fmHLZ517;=cFoCagG3F[\]oVg5=W`dSS7PgN7p?USGlhJ$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI13HS(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
<RZ0bSQ:5DT^<QRHFgZ]jT@IB^Nj=gnaHZW7_e557?<_XHl4We<f4eMHp<gnZU:J
>]mXb_[le5oGbBi2MC_WC`ac>FOFmlMjE?Y`eR>JP]WNAZUm9EZXSbQ>Oq6S]81X
gC5dO=1;Z?6Z5d[O2<j<A2^^Jf;YF0?A0[GiAg=9Ank]ODW>?i<Ak:[;^ge6Q<q=
XfQ^Xq[[_baXBVlZ:6J^EbT6A]fI^l>@7UnYdifi>[6MK4q77jjR@a\5ZOGgb5MY
h7`[JO8BGE;Ah]WqYfl1HZGpeI]CYffDh[Og:F]>e<N_lUT2lK^ep?MN_o1qND7n
?:8V9\>oZX`:KLIcB;HLAc_Y08?eaAC7obCkLQc\eAQ:JNVD<86H3AS@nGQ0N?C[
I0S7Q\`jWjQlQAN6\NFHa]@F122OPA8[HodnJ3BE:e=H`n[77RJ9Ta[OTPmS^5?c
ohp^lLle5;8FVnHn_k>PJUjF_2c;Jo3]UJ=CYJ]Wf_Ih6b[Y>5`O\AmWXGIOW7Mj
9oX^QblcE[4Mi`2^R4d@<`ZGf1A_[3NPS1\bYjn_k]Qnmh566?ngTMON40DK?>Rd
eX4_N045jp\JMS;9PQ<A9ZF=P^g87Cf;<9:19fBC3HV]m9M<]SXdInWRB3H=Ae8A
g3WKOQBN`k\eaU^12NL>g5^D?GT>lBeGVB=_Ij2N[>a]58KTZao>U_c_eKP9J6L]
`Dc=Oh3_[I8=_4JRqQ27D[D?T:XXBcfU6blmLME1295cHD_l7_dH2LSFg6nW_f<?
od6FlFO9H\ZPNAJE]Q^1MD]WlnXP`]O;naG:?eJ6MYY;VF=5KUdiFZ<XleVIfUdj
lkm_aIPDEj0?>JRjXCV03LIp5V;YJ:I_gdbZO<SQLQG44NDnl]M[JC[IBGI[Z:OT
4F5DjKNBM6gYj[J:82<ogVYB5`?E6F2;GdZX0UVPR@G4=N]4>@T9SlN=OGbjUjNT
@eAgHEllZP7N2k1Mgbo3YiLeNnIR2Ypa8h270=gO@1hVO<5o2kJadk^I`Xi]d]:=
HllRgQE3Hq2EJ]P8oS=?2[IjTAkUimDhfH5YMa]Q01CQ@?DUTo7^gj87D[[C[LlA
6W5d><;GY_2iAAB6BX]O7ELXE=:Eof>d?:f[CVVA:11Qn?mZ?=JNT49Q^HCdLB<n
hL:B=H?PkjjNA[ThqAnL3AofGSIO0Za3je1F:<PBAW;M6a_kQ5]?IOo>2cYLM5bb
?Zh8aS`@>^:MS8c6EA==8UY:^JID0dMmm_?FdF]UjQWFce]E2X]WX2ao2I8HYiK=
M=Yk91;c0:]e[X=A<;gE^\_pICe^2K7Qk9JZdijbPFETV1MBa\^;g>HWOT?WnET4
Sce6f?[hn7^d7H89Abd[WhX0If12LO;aT9lZP]4`bCd:FBqnfY5:np1KK5[ZPT;=
>m_KnQSk1N<PDI_h3Bk_O:Ra>7BHC^A95hd2R8^CW@XE8ISmSg^ZVo1GLn8VeVCm
QAaUEAEddpU>QdhG4YOc9ilL<8_J\h0@b^2?F40[Gdi43^gLRl1>?Nl6HW1cBVm=
9`ie:`8``gpIK<?3?GeV\HjK<OlH?SlL1?F<OlA;[^?;32FG\TGBeeF4<>d0cWkW
_FWNjafX9iWIofQA7IknM7E=LKKUAcp]V7Pl<i5o7K5Dl3XoXcG`XR7EaB=jZU\V
6[\e8BU09nd=Io59^8U1l9BlW1=kQT_][9ZQ]8m[k3KDT0>BZjq@YcClIG$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI13HT(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;

//Function Block
`protected
=0@aXSQV5DT^<O3`UObUMDHOD_[QXUKA;BBk4kM:CS5fVVSE7Ni^ImC=Ue=:0361
WfNE33TqJCOQaF8i5Vi`XM9Tj\lUa[FHb?n^TC]>RgGqLJFoS@V3GY:61ojmB2O\
[IOacYpIOHjEnqPJahdST7CA@WlXS6^oj_U;2l>eTVUZ[=jeFgZ:aJpd?`I^X97[
X?oXbm@[C7QZQXk6h@oTlbLqhfN62KGpQN@58Gq[UXKgH6`Z89_I2gTdT1:;TTHj
RLD;lpVKT0CfgMCYXE5^j[m`HNlIgMEh1Sd;KBjQb7QZfRRn8c2bIVIVa5HV36Gj
9IP0UTV7:4ehoSJY@ZHfS[BP0a5jc0cDkX?]Af8Q1YL0?F=iRR^_AYN9Mo\KlYJV
h<OdQhf`Vl59pG]Z_f`Cl9I`MQU:mjWf[_9nZM7;ST0<iQ1nQ`?FdF9VJ`D7U2;e
S=G=F?dbj6YjfG;B3aHZP\L\;f=4=EeG85ZH_F[iP?]fSE1?i:oAU^9`=[o^N^oY
L>;V=k?oi559VCS`FH1pbM5naT5;b<C]kZGmIIEh]jc?YI^mGJ24oSN0_fG@feWN
oJ=[oQbVLfMVclneXo55bIS=AD3hFY7jISmUYPn]0KN2G`cFPFnKTS@RoOgJK^eo
ONSnlmiS>LAYDjmjiaXXFkiLM7pMMEgl]XJLYZWIObB?=fNXFUmmi:__c^DU8H9C
6KS^6nPgK1QEkO`eX8eBWZ_h=i8MY5CX0TfJYYE051^24m@oJgR[36e>`<R]87U_
7Al;eNLbI2C=MY7mNBkhVj6;;gK5i\L]0pbQO;3^No5i2CdGNXpeV<092c7n5@O<
iNLjjdmBBe5MA8W53M8AZEZ\`Hbl;Y<k<h_]J9e_<ARD>8TnADleb[enRI<C5EOL
7XVF_d=X<KT6PXX8VXeSZnomW2Y;Em@FD]:R\WUYC[H9T?QGa@1<=M0RBp8JE_\4
1:YA9c`3ef?CjVPLBb[S95AnPckJmDabKgPfK<R>\hhTU[A5NAd1AoWVQC8YO;:H
UN7A9o]l9kb=j]aA0l1M2F<mE0[JR=GI_OgW@4`mBoXJlF>DJ@SJ\Uj8l56C:Uj`
q]45NVZWhG^P4OCl]=]?4>o_]@67HQ0iLL8LVj8\Pb[7N8M>F<]U;l@@Vg]@?eMW
=]19CZ<Uh0^J;jon?8_?4c3L2ih@nKS;Z<8LWXlUKP9HOog1KL:Q_ZiG]?f3Gn]h
XLM4PhCqUD2>NH2E:SE<Vl[`;Tho=jQea^W<N3@BcI]@af=AOjB2bW=G2D:OcC1f
JLhdb?31UMF>1VU_OS=1XQe:Znhd^VqdQWddApCGh]K7W^8QaW?DX\XLS`5>NB93
a]9:4AWG@_SeKn:=Ej:]Sa397>k7oCN58VKD^bCk\B16Lf]QIW^nP[o?MqBO^Ign
m3dfA]WKpFI]mPF8W1_XN`0[iU36JB4V0_aA1U@=Q9Z37]l_Y>gj<nH4mUCUKc8\
XF@e[Lhj1FUSfVfbF^aVHEojHgAjq6AI\oY>9jB4N4I1@YJX2f1:>Oe[7=FTc?KI
0QF;jin[ERPM`4LJO=<b36T];a<Li6`458^72f0CSFK36<?=qA<CLUH7$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI222H(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
5Nj;cSQ:5DT^<eNML^OdYXSDqkm`X6RH>[IC<YRqKQGZb6fOYHOR9AQY:g7LaY?P
SmnfoLX45j4TqTgjZLKqdRdc=kh@?<JFkf81QN^CaACB5\QE:5k=IKq_4]GA:5nn
2JFFL49JH?RK>E0DPkY;lANomqO[;S_SG6i4f9Z[Sq5[>;LNJjdKU2MmZdVH@ZZ5
5VHVL1C^aDlQqXAX676XoZc\81>_l`8Q9DYOH]ACH_m:TSOfh=]@pBH1ai3RpWXA
3mP<k@OBC7m;1Ekd<I5>>4hNL`Xb]HSI<O_;gi0h`B]m7S;2c4aI?g2kTD^q@lnU
KYpTo5<a^a4e<6cm1?do1<ih\k1[;mnY[7nem@e=aM>2gfMC1E>WF:hl0XO>TQSM
V4`TN:iEO\F\<UjH45jRG`^68DhamA^;RG`[miM0@HLfPbI\9^@R31ejcT0kZ1I9
V@0Te1H>O`D\dQcH45j_HYF8`q\hF?SSUfPocKN@_EGH?UN@M;`X;ec^cQQa^@a4
`:m8@IP99TOZM0Q7A2e??E1B5I\Jl4CU6`YoSAcTFXo][l6GYanR5`:>L7iaaW@V
33B0D9I0Q=FW3JQ4aa16GV`BNB\nh56UHIYmckcTFXSjgG6Nq[DnXJMhfH^WlnRj
^7eMPNblB]a;W9X3BnE4AglaF[oh0h4PA@k]NNYDXFR@cclAJ[CIhP:V[I]Hml=I
E;MMFic\eR`o2;k57eE\@jTH4Gf^<SN=\S?\M63[lOlOc?l2`[K>Xg:nZI^UCl=I
EmO>9N]qIPbKQXRDj:Pc^3dMfXheTMLAL>\Uh>XRZ>X@AJV>To:OI]WUSC;5DedM
1VK2VVheI95iVhj9M:dCPJ>VB<eMf4laEd1591gi4>XV@V?SJPbIN6<`X\[D4Ye0
;=N>1VPZI08Leh?[MCX>PJ>V<<d6`6qfXlM6mPgV_m6G?OWCY_9hQXW;dnZd?^dS
Bn7F]`BKnAC^k0:gQ=2liWl7OSk:dd[fRF^3?I<U_a[Q1lbaJi@AB_CPmjbONk?I
BT4S4g`Ej9\G1NlXnU\21LD@7n@[d>KfW;58?Q=U^VEQ1lbmmTF5`p>SJN9?INle
850gNKH9=e?3XMRXSSkINZQ:2o^DcEkd9@0Jo^;Xb7dO4dEgJUQXR7>^jjUdiDS^
kd\D>GUB=?3K5\_[KoNc[UA:2SRSAlCn5hmcO@KP;Re?5a0fhELXTd>RX27d7<Se
TU\D>GCNk<@9qN\O=hC\C7Oci<Ui;oH?=d8;X?boO=W;OR\<B_j4P^T_3N[ET09D
mEoEdUUO6@dOVlUAhoP?Kp]`S;;>7X=I\4>6<Lm:SnF@m@gag]@PLnjZZ=\maT^Q
]\NdH9TD8EAFHYl?He9f^0]DmaBWn?[I>TWi]\^A07oAX4;27hUO?;eZ8;?bAUo_
gLB[af;hSTd0KjUDISKf49]3Ug0WTZ[n14Wi]\D@Djb]pCXb9lbeIaB5]0TA\1e^
[4LkQD@Kd89=@Ye15FKm48[78l_POkTLaEVn2K_e;]0mUCcbINgNf?9VX:0dNd@R
bC;OLDAdY;:cLbeYGOI6TOb<C@?OPHo1_RZZYThYWh0>JC<[OZgI@?M<i:0dNX7X
K4kqR>ALiT9Xi0oYgZ\HgD;ZB?Hh:cl5PT:h8PiWG76@oelKm]MdkRna_Ud1?b=4
a]7PR:_jIToFd00FK]A6SVKB7?ZH:QY^ie[abPhLF4DY_V:nGUe5a>1:hbImLdAe
9]g4R^DQ1TBQd_BLK]A6kc[cS7pXVIdGojAQdD;K6jf]cW0XEZIKOJ9;RDa3Rb?J
T::ZmOJZ]WSnF[AdhoL[fGm26gjX6kJCOd_odPYICZRlbGiZ<p:VK_BlmGAE00FJ
?N2IFbSKcjT<:j9BF?Nl6XCEkY_A6;Xadd7B^Gj2bQK>EJSH@9:MVlM4=KOVU[QQ
PB1H73fI\hN<kjV^\^Sl@eL[fW3a?G[GbD5m>aQi_2ebEU]HWg:Jam^4`EOV?[QQ
PBknVY5`pM[IIN6YkU\IADkoSp^d?g>hk=a9o>BP321ZW;=6kTZXPCF390L^H6WV
dD<5GUbN9f2Naa8nTbF?f8?RW?^;UC_8[Pg9BAa9nUYHAm>8N3P4NMEXmHX^DMFW
GQQJ0C=m25;:;4DfUd6a??eR>_^HU3n8E8g9V8a9nUJ6o:m9pcQZAO]<JPLNb8Vl
1k0PM_8l3XeFAH]i4cR:bdmOE>a]23>DR<jcHfj8mcdVegDS?cW9]D2=I4;?J9k0
T^\Si[BBmf<<<]C5H;RjFKB>bVSTScJZYg?8kO7E;7e9R^D<ncf?S22S14;`J9k0
TA[2n2=pG2bh?LN]NeZUkNN8aEMZZT0hWXW]Q1SNfVU\91mWCGH32YgVU7gkKVO9
<<1GZKK=G1P4o?YGgd7Zg?fm`=S[5?N<ZiR\kXY0\Vf_cWnJ4Ub57`2M0VRiPTJg
=09QCKeIGbQG9?P4gdSZg?fmK;MOZ3pQiZjI4>7KmAIWKef`6HUDURE7>TTLZL6o
GUTai9TRN\4L<<Pbl\FX?BC3oDR4oGAQA=?>?`[NUD1H_c5a:f24^9T7IJMdnZc4
G[aa=X]m^k1JgUQZoOAYX0PB86cSof[Q8fkc?^5NU;SH_c5F1hL94qO8^Ncm<2XQ
WoeICCM:U]J_]Nh1XL43VOm\g[XnFNfiI<WJXcI[Vi_W6>c6b\CP04OOg>1S4m[X
U87kP_R4TlPh:M4dVa36fNP\>X5dlcXSmo2BA]bj:k0Ho81Ke48P@OO1a9LSU4[X
D87kP_ZZ23EnqPdQWjYI=ajaiN5iHl;3GDCVlI0:E_EHPE2bTM;kcC:>NNF0BI7^
gJ0eePYGDFGYiPNM?L?0R^^\n5N9;bIWag]07QeVJa=eT72RRRf3XbGg8n^2OL`T
AVMnU^J??7G>kPnJHj?2X^^Y[5N9;d>cM@gqc6kIGi7dYalIWYTdR<b]:DIXXgiN
lGD@2IHDoL@XhDkS4P?EcY[VCZd74KIa[PF\c0d[3^;]13cPaL>KB<^=NQVFRgfX
_7\eOIf^<b\2XFTH_L2N5J<]4^^@a<LPnP[Ccjj@J^fn131RaL>K\I6[6?pVU8Ve
NUjhNa]3@MT5F=JWjWb3[XfdFb>9TRUZ5DfV_lS?JPR7BlKajMTT2\O_km]V1U5i
?cHPDOVE2DeeXWg2k4GiK=0\>ImET<<[oXL2\=91`L`:\F5AVnc3`>fMk``V8Q[l
?9ePD3GE2De7>_<@^qb3HYcjZJJk17@gLc<GAF5UUMl>:kXh6_5hh44R9FIWY4Sm
9kp3Ae_b]??>5QB3\Y^JDI6QoF0[ZdXUS_N^U2JD=hB9c:gKWB?V[iEc3l]>C7on
X0P3BW?fQXEd@=B7?LDia0RdTp_A<WMoA2kW_ShF?Vlmo\ldDEGk^k`P2`20F\;B
IDP4JkIdI76ncj9KRceGYXGAU>_>48[eChD81PVLGTmJTdbSCTS6V3;ncok09nN3
h?3CXkbCMeVQhi?W[?5W2a[A63_5IK?e^hD[b0VLGT^KeJMXqPA6m9naXH3gb\OB
JB8J2D[IX4DJU4[h3mkGcC9HdGk:B^=`lGhHRGgef;L3nXZDOP`QmX;H327XFDO>
VYY3Pel[3mWZbABOcZkH?93?e9<H:UiMSXBgk5h68`G?<MZj4Pi0fC;^`2hd:DO>
V^:]FoJp7@i^5nGTmc`>:3O6R33;27P=9O1<@<Q<W>2o908W6VIE]K\FfZciY1P1
DGflI7;M7AOc?^20MW3T[>fVU56R8>\_A4m2a1S?`>Jo^nZ7PUFSPGhj5[mOlO`:
BU46F7NT7Z<LT^QYMjlO[>fVo68\`6qS^;hn?9DFPBUPSRflhYdYKETo@UE@_HW[
LBMS8e<Q5e2Tj7[KaYLRSGDTDWY?RjRS:;N@k57fLnn@5m<WT:D\MI[2EXX\F8GD
L@3g`hU8YOWABeTbM?boXf=3NlTLR[^SiW@_kX]f?Fj@5m<g20iX`q=j[`ncR_Zm
_l5`<POBc4dnQT`o48\a8TFV9d]_69kUH?QBAiCQ1E2J6TbM52G=3M=>6gd0BoiY
;P[EAe0iKmNkDccZ@4TVe]4V959F_=nb:GPXdAa2M`;R<MeZl2O=Ih=>3GO0MWij
^L[EAeL_m1o8pVZlYiAb:?iTNZPT5UKemhR8@TbIEe\kU4;IISYV_mRB[eXNnYUh
fd_[V]82XKN_jVXY<OBfIo`b4;[YN<_nPiK`^4=[V=OJTL;@G4ACLkX[gMKA;4k<
_:bgnZl9IhNM6V>X[FB>EoSV:;[YNlXBD6lqZ0]M^BUmmRRM>Hg8J3fhPRaPj93`
[[coU`b;<D3W6@Wlh1[2B01VRk23<ZGQGaAbZdg?2883WR\[In`Boo;lhn0<I4^_
]bB3D`STl>QIogWH2E3fWVibZ=T_R8C`5aPHZnFCO8T^Wb;6In`BdMePW7p\aTGb
UUAZO^P@h4S]Gon6ho[O;93?XfQ<1l5MGi3;f321LY=S^A07J;^A?a`3lKp?_nhX
`l3ka^KW=I]SelN\IS3jdbl7F<SP1QlJZ<NJ[aNB3W3FL2IJQ_Tg?hmo28W?3<4F
JXWo4LNlRO<<I5I^AH=K?^0i4m4S16_k@YH7]LK\IISgF?NN]GIdY`=L27@?FL5Z
JOJoWaZlRO<4K7D]Qph5D[4oVV4n]iK\6K5INO[15<a@HbNldW_BngC3dQfdWdM]
nk>Bf<Pj]]KXhd7SOQhM:A6ZSoK[<@31c`E=ZZLA=c6SXNnU[j`BnXSKn5A11j6H
_M6ll5Le`dk7k;MS[Mh<nR0ZIaKlRT31c`Q1Hcc<q>lg@OEWT=?U`8B\KUe?j9R;
4=7j0na_58`AY_<:B9077gBTjjh:^?mY<<DDmkZ\N>K?M<1fV<\]3`1]3<Pn[@hp
I?1dl1DLbTK7[[5d7ZVH8lLT5m]lRbjh0W>RMf4kfn4@TRBk8IknIBi0kG6`0oh6
IU`W_>HI<=N_h5THGe0c_5<36WKUTjLZ_W>iV=0;igVS6UKaPY?;4Afb5NB_MoDk
Il`H6>a1<=j\h5TH_oQSTnqVfIXj6mMne[];mNAOL8C=:b0ga6c^=In_P8L1RUa7
i?43??iW;SA_c;MleUi5?1:VKBX=Nk[NYaFk>DE8D1i_f27Bo^]_Na5=P2_CSITo
M]QZHR4o9_]S:79]gQ]_?hNVF1aXNmiNY16k>DEoj^\V3pP23\khnSHjCDhnTF[G
TmA5YYQ:>im3199E?;?=]U]a8Seikoa<3_LANiWWgfS6_DPYD@3_6KRjG<7g3fdO
>1DPUBA;41h5_BDER:8IkV;;YZa<YdF8\G4nO6=^4n>6n5PY;C^_O]Rj2[7g3fi3
Ik@Bq[biG8IoEoQ<17bHRDPP`6EWB:SjolSU0hMZccDEFOJRWG9YSK:SZjZF_d54
UaVIe[A^nPZ]?EV5<K:AcXFX[D]:e@?ILH`k4VM1?e8acJTSZP1jGfjENoA4KHmo
[fVIA[H3?`Z3`EV^WK:Aco=5i^WpC[1_k\\EFP;XkOT_egR1jjH:lN^j;DjEg:Rc
]Wpj?aM?1@5[0L22YcDP?KaB5Ok]\lZSMXIfo50K7Lm?ZnjT^TOb868ZQNAn2Ibo
^FXjh8a\RkYO:Y;FLofoFn3YNLHJX<5d0<@Fo<<W<S@2JAVF;1V?>PMT>>lkYXG^
^BKj>]MjRXjO:IlFLofXei@?kq8]^]\c:NTUQ\kECkcn4dM7S?:hJo49Tka0[D@D
3lkcD:CeSL6]4Ab[?:oa457Eh<8Zid@j]@gU_1jm`K]nPMW0C2D[[19H?QC0hS1T
XmY@GiUnM;\X1eUjnG=?603EV<85?TRjLogUOZjm`KWO=]e9qe]9PPLdGU?6EGJo
hgei4N8G4VP]:?A5G4aR9jiR_U0BGJLCA9b1V0j@SL6[?9m^MehHd`d7P4cFKo=N
1<aNWG?8oG;1Y2H7ZCajBBDJPi=\N?4jHie_jZFfmXoB25m]We4XDadXE4cMKo=N
1:0Z;dKqEkL88RNmLTCW=JARe9ZH>`bX:>6DIP>D_=]Y\PJ:SII7lhAKQ8UEW0oL
LUj^T4YVEb;IG1iWX9U4PiH::ib9ZdCBfUZH3?caU=jeT9akU>XeOBB]P9jkeNd^
I^5aI4D1EDgjc1mWX9TGPiH:9lC;7YqR=1Gl6O0U1F3;JeaJXTm7m;[906aKT>WB
W6h[GPglkh_io\@defoJngg]]Pa8;HCRO2mlhJ36]OCVO6RK6>j?k4d3HCE7X\]Q
W;3]J`O3bN9MJ:aFaiWT6``UnE@R;IiR[^l\hGO6]P5VO6Rm3f<CCqVj_PcalgOX
P<b2WcZD9d8=Cj4oCRX\J;FX3effZKI<:C^l8aOik7V=UCIbT0dSH\VbU`kU=Ld^
Ko_HH][8g5ICpFH2mS8Q8N<e292G3Bmn1oc9X^An@Q<gU:?iBU9N9?85XhmX8Ie^
W2:Sgd0X5=;W]Fimm2:_mCVFgEMkj4LJ2W9bh=Y2BoO]0>?\hXWBPW5fcfcS`KWa
XZjBM_P5PS;`KF\>5Q:^mC]5gEMkjMZI>\1qVkJI1lJ@M=42VncH>me7oUmWIP[F
[0G3]9]V4SDj>^Ce77>W]B^DA;NfI@]n8i^MpcRh5FGfS@_aMO3T:@D`:dE4gDL]
0IkH02gZQGiXWdZn]j;K@:BIfo`I4C;5j7=:ac2936bCeI9=Kb@NiIME:MC3b1U`
AefFiRgL\aTKQ2kWgo]6c3@U]=CNifW:e3=9Ocm`D5b3NI4NGb@NilM8516pCo^o
4]igD8niLG=hR153?P>^:E\Uhf33GIA_P=6]?GPDM779[161Ji:O3Gn<0AYDCL<4
HYiV6jP;khd4n@NR_\bL8a5YamA9`I4Zn20e8>:i3A<EdZidD^BQc1NCbAFoCV?d
?Yac6Lnkkhd4J4\WlYpQ?_090^TG12K^L30jE`oS:X[8d8RQ\FTFec]X1[1`O;il
04cCe>`VH26^F\FPWdGQS2m?LGJOEDc<dIHaWTJUG=\A>C6:HiPTeS]eNW1H5S<i
a`KF3g\iER=1U0F]WWHQ7_>QLe>OE`d<dIHSc8ZlmqMjYI7T773JDMU6YaoYi<FJ
a27jLgY`DUGS[i6^PcMiLcbVbhd8aHP4K:MhLM>fIDM5@D6a>b>L9f4dlUP:m\2D
f]d8igQ]TfMSUZBKTM^6b1B=8kadcH^<k>gaNSEf>JMcbJ[ajk>DQ34dlU0Ma4^_
qjR63l3O_^;EhS4Bo1GR=7`h^;n`=8?hT=GTB:aReq_CIgK2aJmH5=QfNk4lQb;;
^?E@d:Oa]CgnZWeS^\AYEjKW0XY9Cc5JT:o_l<kgiN_FNII:QnW2]NR[lcVkIZAP
HoG<?P:Y4^WnX]V;cJX3c;_gPc7_Yj:@ch3^Om\gMK_Wgc5:@2WZaJR[lc^GIfe^
pnOfmE3Fj]8`N4?Y6HUYRob8aSc<^Co]3FjcZKWWB9[<fKgGGU2o7ol=c9]8KE09
en9M0>c5e9Kb>9J9nWiH?G=;NLL0Pf_TCkj7UdL2G2N]T8J1T@?;8ZC8k^@Mej0e
Vn]mZVc2\9<k]9J9nn447GepaHRLZ3YR?MeOE5acB4]PTP1m0]A63b>J0YKgj8hJ
;oWa>[fCd>WT7EIRAkJVaTZJaa0>J0?TbJI\1UF3]XFWF@79ZfQBn^XWDYSYbL[Z
KZlO;U415f_;T2lRYEXOjTY:aHm[^09bb:J21UF3m:^ld=pY;_RFiReoWHkEo>A]
5X@M=O`8cjkdgN0diMM1ClhObmhJi?Unjc<=425FERSG=6nY6<:IP<dPe5_YKUPU
4BWCa[:6c_@nAf2FiTiEDT02a?M`;:OP@3>WFIeOkgb1=@;Y3<;2Pe@PoVjYKUPj
DkMGCq^F8C[bdS?\<LfeUS>Eh`O[HFVbhSmKXS5\<X=DK\U?D1ATbT<R^p^Ul?O4
2cKUMPE]Z1@YnTZ;oIG2?Bm<gP6AnY[[<^cb4Ia;jheLd884@5>DNmAiB[^jP_9c
h_XVocE^36R1\0ICq_2?i\YXHTZI2U9:YK9^iaKmRSXG>QE9P^?ZT_5SiGe]kD>d
m5MQ;IP`5716P09H?V?RQJ_NL<XQ9QlkaH^<=]F9aj>K?DYcLV0;W>kShIf4Q_ll
HFd[Y7Cl_d][SJBAfP?P[J9NbKX6KQlm\H^<=^:gimap12`bLG=4=]8j]7K=o?^Z
XY`V15<b;5mYBOE@CYOmVSgL567Nlg>RJPd`4RAYPi1W19ANFOn1a?SnLa1WfEGR
XFd6bKBaF:g:mOl3FPTm=A7;gbZ>n<^[6eIH6llRDiUK1nB[^OdOa?4fLa1WNQQ=
IIpb55APRFh@E5NR;220ac2;CJH2OR`XCa[QDZ9e[MaPlloK3AgN4i3TDaRSOkVi
gn6bfc1C]3odcKmkIQdAT\DnEO5\Ka[G__3^DaBQ6CaQZhO>miB;[PZgb;JGDSk>
g>Ibh]FM]iFdcDekIQdPi]OW6pIT_i>3ahBnn>1n>>JOc1:07nkkN9X5`426g3qO
N^QYM;70Mo>LZB40TBN5lV@6k4BIM<NG@6JNL:bO@^_`i>>0RMoMX<Ae\9DLAfJO
deDklN0US<PL]lXfNJ9oFAB95C>PY`n\@keTFlK9dGV];<DH2Q3YmMFYTe?1AYkO
oeKdl7eUSjUL]lXgh3SEkq1PWl>=2PcRRNV4<EFDQW?`07Z_b@90:WM_NYg@\T27
h>5=3Tm:8khgPZH?HAhZ::1mWIMjaAkg;=YknMan8a=T3]d[<;^26Ji_WNEJJDGC
:XZ=MEhhB1eiNoc5gjGZ5V1G:aDj3Hkg3=YknMTP<MX_p08D_Bn4oBDJ;C5_b?Dh
1[P2K3g5FkdElP[W3o`cn`<3AfK4J:RJJQ9YR>H@=TF>H0;HUoYPZ6NfE5kBoS;I
S0Z`CG0M7=f>Z>[Q35;ZjD\]`7blQ\B?S0RoSl28D2F7[0^=C5YKX6N`_5kBo;E4
mR>pQIe\:W;6WZ68[LBdCRQ1h[gH?YSlC4JDjMUHA5TP4d[;1R^AOPE:]ObGLGO<
EYaY;;YN:=GH:LJg9NbKma8>AZS;LaP6hAPYb:gC?]`LF>5i=O]2E\FG8HYJ@oHE
<dF]`;T2:;2CJLgM9NP]ma8>QeTJg6q]MfRT_Dd898Q6LoPJ3_[A58Qj97MHFKH2
@cO`KB9R^Ci`]dcdgZ@fBPb@nUH0lO>]<W<f^>1@]68SA7?96L5M]2DPdWhc[\4E
@V7]@Wlj<g=GD38<oT3UBB1^>odKlNP]]oGa^a_@]YESA7?1ToL?;qFNAZ]:[c;4
G54de8`7B>anCS8\SaHH@F=ImIN_fDF^KbkoeG4Qk4gn8@5aXLniW7FVYn@I0MDE
7[jbSkV41me_Y2[S\UenLIUI^nognhW2mY>;5EaKXNHjN9fV<S^iiPFkn9[IM[DE
C?jbSk85D5:=q==HP4fG9l>hhK\[dIePQm_U2DW;UIfIe=Fg<ik_=0GVH<SSLRJ2
?V0m\=fWYV[ag=cfTZ`6`7iYWB7n6ZAlgZiqmVke=7O]`ck7QbW<Rb:^BnoF5<[q
AWS]g6qD[P3h?c$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI222HP(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
8FFaXSQH5DT^<`HaGX<aKiTDKkMcDVj@3Fh1VPpfJ;P^ABe:7AGGUkI;n_J^k@qR
khH;ZFKAcV1gP::2?hK_7A@ooU]hK8iaaKJ>18_<Umpf]0Go2qMbmPl92loDSN5P
09AN^6WHIhlN<31Od7e^q<kdMIHeB8cDGn<S113eUanBY9o[F<=ATD0pNK9nAcXd
Q]LEf01N^LLoZcRdiY^T2]\F1mqU`9@K@f0\>j?D4o;iW@2AL]^^OnJW<2U4FC6I
:hpDWH^U?hp5F\Am8q25RPKEiG?UMNeY45cGke46cU_j@8WK7AV64G]`;Q`CE>Sn
?k_W@G\@Mm4WnMCR4Q^SpPK\_=Y7bUCmEd0VShY_=ZM50<QBRB=oKRiRXH=lH\8_
HmfE7OF\[2mlfo2gWoJECPM1nR[\:FCjB_j_X<14XjPmX1?eIXM<AfiMo0B=;=4C
eOA65k^EHgRQ9495\FJ^QP34mC[4bFUQ@_j_XgBdTECp06AB8YiinYOXD=WkemX8
6kBW\P1:S^5h]]P;\J3YcklakGg5ffnOTj?aeb4U]];80L7Fd6>4jYjj1^Xa>R8`
NWAcN2Qn:ea6R]6;B6mI\eV1g72Na<m=Tf:c0W@:Q]?h0DN`56==j^Z>1^Xa8jfQ
^epKUSH43ibU_<L\66gWZ;m[=>aKE0P]6eHeQGN<_FPY\Q1B0C[ZSJ>2oS9;XUkG
md0K5m?0VXgRX_64Y<R[@;cIIQTGeb8g?WC2QdB:VgKBFACAUboPPSibY8WggmNe
mNMKFG?<VCMR_Sa4Y<Rk1[mA0pAHAGeC<dQe9:;gZiP_MZkJN13A[SWbAZXHFJ<I
JFDV1lQ7?P<fiEPDeAVd=_3fjCA1=O8gMTLSG=gDPR^2MLkKi9Kmk8dGD@PHO09U
?Z:ZiEYULhE;:K:>ZHJoWT2fLCAemJbg8bLeI[gDPREh^el]qUmnlLMD\Vj46G`Y
pL1L1:o`YbYa7RPdG3fEb9:]UNPUd^d@FFIceUY@3PUcmiH1FH6d@\Y2WMB=T\L<
1L\E``fd]=Y671oM37bXWTh1KLR0<<0L_GI7_=;9UISO45:gl\ZW04O4Q72]F:L?
MLh\n7fH9=b^Z1oM35LC;DGqLWTMQbD=?\o8L>bQPF^HioE^gdhJH`CMe\bPkl_R
E2Kf2kf>0>:CU=3BGU=KI]4kL^?HbGbD[PcbN8\h\e^n0d8CLi1kmaFaX\iYXW3E
;GI7hfZM\;KXXHY`\D_8I]I[L3LiaG__[\6aN8\hf^PQKPqT6CXeIh[DV1OI<Xji
F8c]E>Sk[^N^laFOBR\0>l2WDRlXC?fmP_OL2lo4`bYCXM`TjMJ_:\WfVG:BPl3E
ST@h]L1E?N=dZ<H[B\C]Zh06aDa1:3N349>D6;R`31<?XdhTf1ZB:[Uf_JjBPl3m
:;R7VqS_[T:_`YZlC3XTAE>?kRI7=:h1a4EM3iAADJG1f128QLXkUA\Gc]e:Nd35
OR>SLcSS^fNJn<Lh@obGSO6CKokX>WEO2YSINDdACjGZWSkgYY@`>g31:P912WZ5
1?MShmS5ig=JLNLhYHbGSO`SJ?]NqS;K5B:3Ielo6R;E<6jE3a]?^HoAXYAkTi7>
J[TWTh:XbaNcoNDZni0bImRBIDYScS@aHF]aPPlij[CQ5JMK>=_o@IagNO=N557A
YO_@Rd8RXjk;G;5`c<SIY82fmdYYdSGM=D]UCPa<G[CQ5KL;06gpF52?he^^FdFe
\gf0dgHSC7oC]51V=jeAAIQ>9>[:`HK[:7ep]iU:KGVA>bbH?5U^F=h\EH?XINYE
kn`G[ioC77o1^?I4JA3mkIKaMQ;mNGWOPUM2]4^D<LU44bP19?CeIc?097pB:1dd
_@OHEbOOao_YFL]0<mlVKPo;5WIL2oSBDQQYkI@\RB1gM5HOP@>h[E;U4=^B9KJ`
^VB=cPX5Gl^[UQ4Ro6S3VTio;U2<2\SnEF@RiK8ik7C<2go=TVE1FMeS4^=B7`1K
^8B=c4G5Gl^DILb8Cq>fR=f9kgkHVf?60cTD^U>@NP?W5hZ9BX`IeVV0j:oc:?VN
@QL1:na<19a@m<C4>@>L18\NBUSVNMYlh<S<m6WjKm=N];o\`2kIo\08cKH4Yhco
KV9oTM_NM_S_7oR4VO>lO1`N86SV6fYlh<UTI0BoplT<6VOMm]MZ\gIREdMj\]L?
D5Q4:GFD8Ml9?V1mT`^NN0kj?BM;\ji[H3SA8\5PMl_9<j5`PoG^aD8m>5@c^DiG
DO7Q2fMW8dl9ol[@1^\S7Y>j6EO016@mf<OiaJ5gglRT\85nIoG@4D8m>cW<cTSp
mo:D]4]d[CnkLjWf^@d;Yfc0XlV1=BNK^IOK91DgA[Ie@:V<U1E]BRXMaiF36Gg>
mhL>0ZR=^Mc0E@WU_P>S^5?;a2lZW41`iI5QYolD_OeM55bZ_nhM>8eniAZO]GOl
m;KAbZ2F^MnUE@WUB07XCWp7RVKHbcjMDNO_G9JJOC_DTPcDa6fPh=I7m;<PULgI
=`7De`8ic:I_@c2=FCEE>iQ7E_i7bHL7=Qb2I20fIZ;c60`TGFIWMnU3md]]Ce=g
TTi;8oKG4=Q_CH@o=bgK>LQ7l7ULbQT7=H22I20W9WcFGqh=0@F3_D[bb?C1`STg
hNRgN_g7f32Od<>L6Bgl9cf;CKij=lH@^@B]dZ1Db`T]_Bhn[?h@F96<U\bdDE54
\UAliUB7^4km6HHLaEI@l=Pc4<00FVSRUE`Rlj9I1YZ]AWh]M[J@[j6<<\bdDEiC
IQ`PpZ>RKB[PI:1:AG2oRc6O]]@9V4fa`KMN3bWZV<N01]nN>7<Tq954`nWQ3i`m
[4RjNO9[lTM29QKGVCcdA[G6<OgahPDBEL73S>eW1b`6`XTILeJ<H9Ti=VaOffdn
4RT7an0Nm<FThoGXF?AgYaGGTnO3lBRhIEnFi4Q5<Z4BR2IdISJ\692E2ca@6fd1
0RT7aPomXElqR[_:HY0NNjcW^UN:0S9l<\jXlF=9;YGkKcjRRScCJE@QUKnPJ;M4
?NK2HF1d^8lPR91ohR`IR1`\Tmgl_jK`]fm<;I7B^J1^BcOWaY8jGLZL=EVe<oJ<
aBXNQi1=a8?]R0lACRE0R1OETmglWN6lXMqo213P>@:L_ZiK=T]7SC72c0Sdn3@[
Ua81HjG8D@>LNih7AC6PDI8e<ORadIP]cUUod<AhMGT9oAV?i^LcV4Ciak7H^`07
hW0oHFSk\L=gNb@Z8nT22]YKg3_S7RgccPnoHQ3eM?59o[V?i^LQLU0[mpaNd@AK
?`^JcM<VH>`ghCWV8jF[_o\k<4clWod6fe><B;0Fcl<=j^W[BMGCLcT8==aH3aT5
SXYNkB3;DXc03[]GpjB7WoLN2CHBa_I>42:1UK]dLo:0i;]e9[94h>YN8^kmB>Y6
1<mid=8`g>AhY4lY4jh6><JC4hPYFHFUXZ1N5>9@0b:SC4>fhb9[IoMJ_LXK<9LI
Hdafkl@d^_`_Wcl<=jcFV]JRahW?gHFUXPc_]Hhq?P0^Z6^M8;Q0[aE>3chnJD\U
F4HfCO`Y[cOOE1L?i]3<^mK=Tn<C=Y3e1kTi_Xk7?oQcEZ:JW^gkMOb=ejQ2b3Ah
]IWdiTkUZcB33IM84;ZKZMTS8<:i;aV@A48BHX7<??k?HZDNWP:YMOb=311RQmpU
JWCh<Ck^bAcY0S7:JSWZAYG1hGE;Y2>38=?>]1PWUhaQhBJKSo1O4EkUFUKl3\ZY
7OLp2I:6A>?\Z5f?U9S3a^GSF_==Ylc=YL89<FGLic?[>NB___@41imC5YkE;A5>
RL2A2F6cM=i1SC2b9d=o_LjcJDa^mlfVTi>4oFgWPSa3oi[fSMacNP`L0ORQQA6R
_Lac22ZgB=W>S4i=9d=o>:C1fDp21;Yko7dOY[fI5ji0`eSZ?CNQOTY?U2X10IkZ
A=\;mnciOol@7Ii`A38<aRcoYCP2Gl=JNP@iVP91D02\RkWIU>U1aj08_\dS0\\_
C1OVUCUQL_Zle@f=R5om3AZ]YYN2jlNLNeJiiL91D02>S_]GBpZfHEFI50k2<0Ra
TC@<AfjQ6TJPl02gkXEEA<T80E76jf8aBZZ5XjcJ4\XWWBg@OFZPd_Te\T<Q9Xni
>BhhXDCdYkBRSiCZja[E5Hb0F[dNTV6EKH4doY4DR09U2a>@GFZHWfnegT<I1Gni
>B;L>QhcqV5WCGW>EU_ZMO[<BPaVXRVHLhjnFUV=h6a=DUecV0h2LQ^o=\eR>OR]
4d36T8?bAVnG\5Ri4gUZf^^1GUNP:^mKW6U1lT?IcWaSFG<meRQYoW4=j=7@M\8b
SKKkN4?B0VlKYiRcUgmRZ^^1G]Rnn9eqiDN7E>deUem7ZLLRUKXL@^TZ0303j3KE
;0:bgIRJlZXY]UW4\SD=PS^]m>UT5^S4iB4UFQYLWe4HJMh3iW927Lbi41lhn?kD
W0Sc^;A@k8`_^Z22TUEA7^;SElP8G^=_ijcABQLfW=>fJMh3<V>_S6qT5FKhgNV_
mmg7FdMf`EfiPG0C?;<N_7P9CgjW0<RD]:A`^lfkOCAI`;fW=aAf^b>TJ[N`3j]G
0@b8ZKPooOlPBA^i:85\NgCjCgRXKk\I:XJI3e>ok`9NA[?MLW4S^o6T8[iV3EMG
0NG8ZKPaGk4J4q40YjWHZDBf=I@9b?R=MF?XMm3UND\8hYHWj3^][O@DOe9oB9VF
6dZOUi_hV@>H;N4eMj8YfCeki5lWC\2YT;oUEA^[KMI^b:SW6eX9V>:Qda<\NdRj
bWe9^AF;W[bHNm4MDTEYIIenZ4lWC\iXG;C@qTBZINTZNU=D:j@I`E\UfKYEnU\m
d^8jY<SiS\IJn<]R6L74qTkOEm`S30ebW=R;G2i\0nJZ00A<GkF_QhVk7BUPiEZ4
OEllo^KCDk:hjFa6=5Dd`T`lL@k1k8;FQ1;9kL`iDM8qMfIBRMdHhK;`Z@R`JK9c
`VJGh?nIO4\n;8lNooC\f=[_@CNVSl>>NA>d6BJ2_6g:MZ@oAYTo6P_jbKJL9\8Z
Tk3FlOGL1[_DM8<Y17]>>c9G]=nK?HS6N0ZKG:@b065eMQd1:Y3Y6PAcbKJLF[2K
YPq2d9]K8k2W>mcSG7U04=E6kTlfmdKjao3JJYI2M@k\hb0CGNNfnfgT0D0>h61^
oQ]2E:oW2KXF3V1[Lo@TLmY9A[m_bCNa>A^1JE;j8FA^9iA@_WQjH4FN^@90gReh
oSX2LPOl2kKF3V;[Lo@P2Y;i1qio849WcG_m8@20kI]=klJeG\QlcM2j2HU<]F[R
VRLK>5;@\9ULjjHj4KK4G<_W>VidDg@Qj98eN]YXh1_F`MN>0YEee[A9Uj7<0hNk
[W@0^9=MBF>IJ[k\7GX[C=IWfViJhg_Qij8ee:YXh106baj2q]2AHLhdoTj;V_Oe
i3FTPf8<Oc`\gi]533[a;\T0K9i@aKJ>]ikfZBWbUn^X\51B6]_h0HIHANfMif8l
F[e?HN[Oga8;30_D^Q[lC;OAaH_3ZfHgK0FG4l4I\lVhT116e]8mfJIMZNfK=f8l
FLJ9TBmqJn2HB@`>\DbL9lhiQJV\Xaf`4Ui5C>1<QQSdm?nA1[K@nLkc_@6oe[I:
5U[3gl7>p54JlhEi9^f;Ml^;o]]KI^=i@fKFmHO_^^@`9C`UUK;RMd\Mj9Ii_W3;
HPkkRU;1d5=^A:IUh;@\kDfea6C7J`20Nb0EJ3EN=C@`RZBi_[9Y>abQ5;Fc<[6@
>;IlnP;ZD5i:3FIOR;@0UDfeaVJRl99qH`=UhBc@ZLP[A?[Ua:F1NHS0YlM7449[
>R7M1HCTh:f_PP0YNU[k^E1A5hMS:b3fHl;\n\AJ\Gb3UDb^SP\GQgboLh^?6:NW
IRBCJ=VI85:gPJo_>OWaeHAQT?do=bfKHZ;39\dO\GU?UDb^j]H1;;pBX^a8@1j0
M`e1=ULo8i1;UnnkR1K3G6V4kjP9g;oCZHbcMIT:9Yi]bNG?DL^`mHYB=eaYCE<k
ZL5I]7[R6^N]mfUhN6SILd1Hkfal_N8B1N;7gFHBdV`\4a4G5a:nm[6BZK=8CB2k
ZC8I]7[VF2:X1pLO8\@8mZ_?cZ4cKPaBnhkEj_E=dmS>Umn[bL:_U8OSDcJgmhbh
W6WY5ID5Pj?PLdLO1Po5h^jb:_2@4b_ETlADGTalTKfNN>d[:6FTM^lPS>k0g`0N
Z`R^cigc0QhP:_LAf885MCjbeU2@4bhKBfQ2qEZTZ1SJYfd]lPij5<PaIYI3<jn1
6=^h:L:8KUAXG=81TQ\D@p>4n<YW_H`gVN\o=JiE@AKQ4<=8Voo[f7A2fTXRgPi?
:^^aESiG`RB]EN9S?YH]Z:>5jSI=f=_j8k_VQXYZf91YK^JG_mjLbN62AIQ>k:Qb
iVhfGjFnLVYTMK_YJL?]e:>c55N=Le_jMk_VQXTbQSS=qEm;WbY_dRoO[8fN]_M1
[^KlFIhhU9=1@Ik4li4G;A>]a<SDY9nhM3W5F]^mHTI\3E0SGGdcUjMVhd^=Fb5l
>b8p@1_YbclGNb`h4=_`9TT?]1T1K2Cc27RRI6HmG]289H;11mJ7SiKL_B?9jO8=
4WPL@5RLVIQ]^GcmMLf`QC9HhlMZUiJm@QI<26O6:meVT;nFbj8;06AcNJl3bX5<
cWjV@14mmIPX^Fd6MLf`FdB1M_q5CiO@=_3R028IS7AbTPH6NQ6e8oomfElW;n:V
N5=GL5c_Dfh>PAFTO2]UT]G4QbJ5fP0nBnZnF]9ln1I_ZU\B60FMnO^4VXL[;L16
@d@>bPi648m@M4?2FFb5Re1oQ=o52ZP\BdBn8BUln1I1><57cqhB75o2d97[D26k
jX[MnMA@cCd]JK9K^fgWYmm0[cdV[?3KESdn]6jRdfEklhgLC3hOk:5Af;_PaoR^
kTdKTaa72b;CX`oAT_KWRIm]>gg3kdWDbQ@jPYLPJMglGImLfOhU1>gAWV_f^_R^
kT5L`KPWpYM[k5M_j\@?3h6>@gF_@_aT1UW8]DdP[MAN176>@Kn]e5D2:TD>JM@S
KLFP?=hCbYUH3=H3WPPcQk`f74Rf0R`[3OW\<ARHN`A?ce[1?aZY3>GQhgECmU\P
0^FNHUhERY619]HeLPHe4k`f7UUgf8?pEn=dLei]9Tgg_2Wf3?MP_?9PbIK;QKaX
EaVb:o@QAoFQ;dZ12d:U0gdD8m4Do^VHEQXJR=k]_PJc=BRSg]<N6gcO[a6efloU
AaYbX=6\mmKo6I@VM;T=C=:Dd<[bb^d`Efj?[=:]_1EF=BRSSfX9RHpeXhXnYnc9
4O?^014T?lIZF;BncSU3OU\M]Ij4P05D6niY9=P@Pe`a;>3L;f[1iQGeAaXP@FZB
iZ2jBL4oK;cGJ^^>T_dYH_IF]L\NfC]Eg[ZBQL\0c><jHe7SZ1b4i17eR6NJ@NZB
6Q2jBL4fh_:9CpDBDP;89LCC8NgE]bkVTaF5cEPJjP^TZdLod@5VBlKQQ=Ve8Hg@
BGP:I0Gj[iKSP^DfIm:c[N>mDlcT59[Wn`h06`;iM:\f^=foQ\6mHC5Cmm;1@OIR
`8[F?gCAEj3SAQDZjPUc3N>loJcT59NKlf8Vq12NWlghH0]5o>?E`a]bmJMoJiRS
e[`c`ODJLUjaWp=SW:n1IE9H=_RjD@\>[37dJ6HngGFk:1Y=cW0=U7BQ\OJHLL;d
i<`FQKg44UGRBE=Om67AM;791im2OFkaH`Yk;]2<_WHoEE6=dEOUIl]lZXkdMAnC
OM>\ZK\^bWbRTZ=KA6TA6@76g_m2OFVf>kRJp:UVL\i:NWFhX@Pj>K:2h3jOnniK
:^?YJL<TK:HUSI`81aXRQocb`SS3_RmoHL7JA:82hY;2EomG?5j<NDZEih_hRjC0
H;ok<4<Q]CaoM@YiI^6fgU=5kmH<cYDjYJ7b1:]ZFD;@6oDZK5j<NHMBG8lqc>L3
jInDQ<:Hmkh:Z[8?THNJ[V9k87HJ`h62VlTRR^S>DFhXJae^mFN;=@CR74?lcP5_
;H_JifaEE6imCDZj_4qd1LK:Chh8`lfF:FTb_Y?03LG9X80n<YHE:7\EOC6QI3G@
QT@ZH5b[>TI;[>A469?d6YE\BZZ[?Ra6OOn2a@IT6DO4GUVg9?;E:_0YHaQ\No9;
ZQO1IaAIVOLCX?Ga6GJd:DDPBj`[?X56OOnUO5La9pIUF`=?@0@9CUZ=;jUACJMP
I9`kURZ>4^RO\1ngE6oPbb``AWoXInC>@<P\[gh1Q;IlG=`HSnVN3TX9ehKW:QXl
f>JLUnP`9]7Od[hDARHZNoQcCK111l?:53_[h;e1DNIcODlHddVNE;X9ehiEen=^
qjSe<^XAR^nUCM3TP1OXWi5c]5IVHNZ6Gl_HF1TT4>MYl6CAd3L>Ajo5XMF]jlKE
kj:nTJ4i9G7JTo[=cFSlV1;Hh7ZSERJ>H5_OmD`[B1;NSPcjF@Eb=\0ZF06I2AKf
^j=MOO4H9G7Cno[=cNEk20=pDe396DCTGYKUR?UYaBHoaN1LmoXcTUNcf2CI6`7c
0?9F07TBG6FmZVoh@DIlE4E9DGSi0P\UWRE:4^DbnU7:O:c=N3JI21a7R22IWfd3
j4BH7=6FXKcnCk80c6YE34UKDem5PPheWR[J4^DbADi5oVpS;G408Fm0mETfhTcL
m;^6]eg?d>LX\Y50e;IbcqTEOB[K^2:5HNHR?Y;lYk>G_k?ViTOI9\W0Ne@lHM\J
Ef_POmfDhf;<=c_;k:7>Y]T;iBVIW`5mP:IkQdee2DDJd0SGEb2V@FV0UMV1ZQnM
il3WoSKi\aF2gRe2jN4>EAT9>`cIcM5mlHIkQd[]5KD7pQB6V<3ROaUI8\\9B5oQ
NFZj`B=DZKnHZd<RSjLYm=S:Vb0[YibFj=6EFfbXWK8EGQ1gPJTc6cLH2]iMIL0I
Dk`7P?oVGYB3oK<_6_DL>XaMF=5c<2O9VLP5C9QDQM8iAQM^:gTWncL`0]iMIQEW
2k[pJecn<APJF0aOAH:P4SC]:4dDVh^e_S`jEC2[n6^GFh2X;6D?B7__EZRjmVT9
4]lVA7G:dZ51U:7a3YNL[TVcoB96NJSN7WnhNYQa3eOJ?U1=HB;2Pn_`JCQG3Cm@
K`XGh7WidL:Ak:GL3Y?d[TVcNKO6iUpC@Lgg:75HQ?AhBi2bI9Bhd=2;nC9526oF
nhQE0_EK^NZoYkUZMbCncC3g@:SGjN7CVelQ4AWo>W=JN6Fa\bZoUNk39]2nYToL
n_SY:[JN6a>Ioh\N?mH6>I]dT7[1j^7CXl2M4`@o>8WJN6F6co>3:qMaOeH47X?e
94W>JVcTo\?il0DO;kLYkHIf6kKBm_BKe<hPTm_DWkNF9EkTJPj<OjMMeA_kE0fW
;8d\T\NGW>UO9m6Oa8:=EGRfMVoi:l6JBX@7W==6U1^OKk_eBE?<h?M^;X:k7nfW
]8d\T\i5L453ql0i0oN7l8KEgIj5CZ`7D6iP0>`@088bfh1F`V6DBV4FSYEZ9g?j
2LUUJRCZ2IM=3lCIA[R?TTlPUeZEiRWBe26qJJa<[GqJP8Y6:8$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI222HT(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
i@F65SQH5DT^<4F1]>E>jY8[hPb1W?B;I^8Z0Sdi81Bf>YV;ChMp3Ll0DT=DM2^=
Yj9j>Wmqk\<b@DJDGZ0J`DZ0>8YqP6nk5Qq1W=551STSnCaiMDIK5I1IBT6eOJ0:
MFoMHpD`681QFAX>W`^2ANOk64S1_4oaMT6;P7@lphXoiWP2\F2E7KYT5AD:^I:J
kHii2<NCkgdqC>m6=Q;X>YS\7^P`m]a3hj?RHco31YcmBjE>`KRqT3B2EM3pYHkP
L?qC1J;oC]_1NNkFTN>3G?1I[?0aSWXFT<2A5ajSBb4fdU3;MUQSjn>8jGm=^[Nn
bKkC\XVb^ldBNn9]VJIINO;\;7DKon1801L356C7Ui<A;:GXO<E^ffkYm0F3mf>R
bEhC4;;D^OHBUR^]VJIT7eBC4qe14WIeQWLENa?L:>CTCh=]ARL4cd6jjOQKDA90
SJq8:7je[dk2BPCGeF:gP:Mf3X]aU5i`hmane<fXH=XfhQ3oI7LZMiOmDH5?R7N:
\ZJ87RQnYSY>B[OS>4WgCiOT4Rk9<OJ:19R[eaLgZeJ6EB_>Qa8khF;S;@a6SM;c
\c68Y8>5Yh6>l]?S>4WoC9TQhqEhcfMo1USNM:D9hLRY@iZKC:`CHUoP8<7Em50E
n[g<[ROKCU\nP;5c4K^`35UR:MEH3TbmJFXaWQ\WGSmL@onB\>2^YXTM]9eE\M;I
6EZ@l^M34H6d4=3kbgZhld2RR;Ee<>fmE?XNX?\WGS[_6c;5q[k]ajjgbcF>=eTM
S<>KFT8FQLmYSGYJi>iWm6bTJiWUQlY=<JA4M<lb>gSEL9@<0[nD:]aaInMlBbd1
>I>KQO6nAejXgfDoZhi7R;:l`Yca@a?GP`8XQ3``\;nL[j@AO[ITLGaUHnFL=bd1
>jUY;XmpS6^d_\Ooi\E_aC2DUL]0XYHn\ee]b;PLi0\8aR9``ALj6nShOAQdo]@2
=b_0j\iPSM[<OJUKJ\f<81S=KJ[J4T6oY3gblL7bG0iMOnAihHgcDY^=dQN^JU1n
XN<OU\heSO3h_JH7J`kj81S=n_5=[hq5`:l@EbDfhIC8Lgm2kaC8[nRY^^<XSnfB
B;<15f5V0=^`Y3FC;W1LkCM7_8XCoJ05nX=cE\?33SCgVE[o0adk5R]PB8J:4f@X
BZPRhnhBBA6=a\ZJS[:0V4KZYdhho095N:ECEJB3hg?gVE[9DjRKjqlT_hl=OH34
KmV:mlH8=aeFRmkCH4g`JL;3nOi\imN;WVPZckHOMJi?TWRkJITTkIl6XCgogXQ4
530SoebFdlhnjijmhDAIFQJ3GOU^7AW>Q@GK\3I^]kVdE;E;KeXT23lT0i_oh5QE
i80SoeL3Xo=WqH8E7b[?23eIj@@Y6d2CShG[Cg[FHhiEAX]BS_XU_3O=KK>aFFg7
hdkUT8j[19mmaH<>eh@WJP=A<0VU@lRU^`Rlj9I8?Z]AWh]M[J@[j6<nAbIg7d4\
;AliUB7i4km6HHLaEI@l=PcJ<0VU@[I?X37pJNfQ<6@oj=LLKnTh9lhC:6C5c[V6
F`L0VVE\k6^7WYZ_MJRK3<9<A8o^`9\jmELoJVP4G>jYl=RSX[h]`=Aj^cU;?J5J
g=EabVQDhGTW4<?GH\mS_Z0Bc@Hl2]:1?E`HJQ30g>5Gl4HLX[h]:970@aqDLmF]
G?c37XmW[i]CAA4J?N>10::J:d6ladX?5k@=f]]LkNIjn0n5GNbNEW;f:`GI4oLK
H8]qjMUNCCLjYSL;WX29@gY1?^eba;Egg8M3C]M0CnommTk31LD^4o9Ee?Ga67;b
Sd;XjBggbAH8WSMWFg3k8mH9nhqI=NKV310Gj=caLi[f]Wl70@bSA9US5ci8\HD<
eJ3kc8E2No@P^V5Q@3l;_Xgl>P@IXH2>OPnm=e]a<b748SD2`oA9d7]`ehMD\H=e
3V2_92PYeV]EWPQ<cXbM1]]U>X2IdAd6OnGm=\]a<b7no3C8=q0dF[dD=>`\46;1
mlog:OJ?lDf>RcJo=FMlj[`[O?3=YZ]8=iG^C`BDnn=ebo4jIK0S]=1=<dF:5]Me
GC`RI>cGeXJnbeM]lG^la<QMCYM[kP5Y1@8T4BQWlV;B@BFjkG0EenU=:hF:B?Me
GC?6GUd7q\8Qg9b\4V3Yj]K>PG[MH6if4@b9LaU:kI:SY;F=ORIfg5di^QE[20SO
ObiFBF:WH\<oV9F]6L:E0H7KCf`FB5^Gaca0JF9KEF:jkK2X=\Zn04IAl7a_h5H0
:2KnT6:B\\o8<NFAfL:\4H7KC;WBk7=q5M9?gimcfe<CokmEC9[mGk:BeM`;DhFY
km^jXIDL5m[WkLeSM^L^[emdKcg4>:8D5E\OEH0hVJ=SN9_aa;^A\bi=CGg8ca]B
Dm:F`niS\UG9XUV71]5JD=37Q5XiI:8T5DN?3H;OVJXSN9_a:3:3?VqeM1UC[BQH
G1l;]gNd`EXaai:gQ?9HoL_U[l;S2`UFh8[ZR?5KYUMdS6eK8iVEFCLeJCA@h?eD
=g@k=k8[37mm;DF6KaGec0SQ[XAhHLJXT]4S[nHF`I_feYOm@o^cF3Me:D\Ih9MD
=l;k=k8biRU7Vq267QL^_eU@QNH<j3BlJ3VOB5nm<2YNAD?TIlklW9X:gq8^N=Q\
@AQHHV_3aWGKd_lJ:TSbT89m6_1kKBEJ_a`;BiQGh`2GJGacYQ:m:Me_ik8I\<lC
;E]8B2^WJKE9Y^_=L35ma1c8YnGk:g81QO9KVM;IGKI]RC38@H\e8?k_7X83ibYC
ih]888^WJK2ZK>f0qR>Y\0Hg@aMBheiL[;`S?3`E9hOG2C22=Y5?h=QXF<DZIRbn
=c<6`RimlhB:EgT7fRb9Noc=SlYfTo\JSPS8c\Cc[jQU>6UCN75cD9Zeke`[2FTP
=_I;4dhB9L<K[?TH8R2[]dcNRlYZTo\JSHR3?e<pmBmgNd<M?3P6oFNjUcbPPl]=
>?En?ERjbh7e3[K6bUOU]Sn^Z?gSNb?Zf]M=:Tn9m<bjkEofknAiNnmPa`hO3e]c
7VXZbd`\HhMaaPS_Mkf_Abd=;S55\THUI2GkeT0kmTFgWE^OknbANnmP`;JcAepE
Ji<h855D7<Lc\A_aiknZinEY]X2PWcfi?G`KVFbG=:Pma1NMPk5HNancGePJ>>QE
oF;o9nX7Aj=B;T71h^gaMRN>QZVT\eLX?GOoWaFiLRM3Q:B8iY4iX@TVO@\6>[3E
UkD[93n7AYhB;T7dV6WCJqWc3jVl8OVHc]<K\3OXgdYX_1\2[bDNKk22A@X5O6I;
GUNdfTL<G]gQ>\h0iJ@J`5WG28]\OEdKZZUGc9nn_c;hqAeM\?LA;_U:W:=<2Wib
go:oR<V2ic<Ri0Of8ZdeN_3n1KgD1RW=;MomfV?b51<:SAbI\55O>86Z=J>aKHW9
>[b;B\V@N<`K2MO53LI75jca:dnDmN>DkdMah5cZE;<iJAFeFK5]c8mQZJ>aK>ki
AAiqS3BA=O8U1iNo\BSeE[AfgL7cPDjWN99f`QhERFVUOWbeQP^YNPjJ\SUD]2L]
2JW_SDYYZi8VOAe[O<i[<0hB[P7Q?0Y4PAlMBQKIbDGKVnENWASDn^]WXJe14EM[
`JIUSPA?RiLoOUfkO<i[[V<ck7pAc2nDGC^Xb9PSDpegQK\i`TUL\L0BnlJW2Mdd
UF7l9FjV55O1X6J7kWgmUPcmA`EGhn2@XR7\@I72CaeWlJV6DoZW>SITUgFY<>`A
LI=jmbMJG_K1b2=oZGEbUZbQnA5YE;T]:?WXJY623ee^KcI68NZ1BHITUgR5?MK1
pW]:2k38@;]>V@:?P6cHL;Dh_lkOYP3kOSO7?0DR2baQe`=3eiX:acV[7ADJ;f;V
hWI?@<eL[J?[=Pfj`oi@Jl;<8Ok_]0U9ATOi8c]4WjemhN[njYb:[2SJfeYXPF;Y
8WSAfneNNJN?XPfj`ETnJK[qAnHRC@Eg=NXHIgOKKYW`hVX]FP_[GghUb8?UBQlU
Hk>e]aa7ZGNGSNcilMlDW;fCASodYYFcoGVUK?Kh3F2co\H]JVAVkLZ]Y8@m3^dP
P_\V1C7F4K\3lH;e1mJTQ;KLA`KS_YmfoZ73K?Khk3j`Dlp;>3fQ74a=aQj@HAJT
doB>NAX6_`4MU^45>WA6SkWo=Q<]>70X<o\R6EEJTJ=BEcN;LicbUX;JR`2Be0IZ
AmkBI1fcco05]cm0><>eF1WKDE<M_BF4;QL\ZhlbHOc5Em^;cghnU_;J_^MBe0Il
5bTl[qd^WYI<jJ`8bgUe712BH0Nhla7FkSdE@C90YDDdCkAUDd^ZSn`80NljI2Xb
CKGUj\d7RnPo2[683N<X?:4oH7L]VmCfFmZIAP80YlWjmSCR2CTbAj><0n>[7:bi
X7IUVSd0SY5o6g6@XK<X?:Z=bdXXqIS0RlEBQB1PUFMi6`Zm=k2b;3k5GeSYNClA
LS2=B:LW2mPoaLeI3cYJVTL68aQZFI[<E:nFKC?O5jDlGGKAc9ZH7g`T<UkH\Rlf
I5Yg\XjZg4L_elICDaSQ8^n^@ZQS\I0M]HnJ?CA6ljDlGD9=dnSq8P3E525gnKbT
TgYAT4HPM_:jngn?iXOe0X]C@5]gY3`4B=n2;mS7N[A861kAW5178j2kJ8mZXXc?
FV33PJG[CL_^\J52][ibDXoR7TC<SlHYR5KW:a^CMh`ROfV_M5Z78hkVM8jYXe@f
FV33eVb:E?p1`W\db]7lbk0_Kb_:]V>0@K4Hco=cAG?kN9InS2X\WV1n>VQ3;:eP
MKDOlSoYd`71IO0eX3b5AfMF`f\mG^4clq>IAoSJ?>cL\jOYmGEGMik03GQ^mBIM
[WcP=?hDbB<nZ83DG;QY:BOmH>FD<8oWKf>;cmTOEASOOWS`f5I8cLGe@OUaRHGh
OTcPhKoRah>3lFG6HVKWa6eXmEcjkYSW:f>jbZZOY^SOOAS`f56^SELdq0:OO_N<
h_ToCLP=P]LN;LgmERoJ0JIQJ?i?0_]`0c93dOM^FnED<OjQRq2SZ<5:libA=oN:
TC=<aH=DjKcKkDGJj8[3hXGNG`a5XgTQZE^cg1>Me0mk1P0aX`2\6=>S??QUiOSQ
5mNOWlFMV>fL:8\01G:3:?aE>k<A5h4BTbLW><7nKC_;FC>aQR2>lI<SLGQUliSQ
5mL8OGVapAT?VH<fL_U2ee8_iIln]DgO4K;MHSe?4Rbgg1LFSW3=@8oCFf_>ZJFV
<:dOV]cC:AP]8j3?FfC11DJH>`e5i>ieX>=?gg=L38bgSN_\ZML9ITQc6?^]FeL@
;HRREGcVJA=SSR3B3fCeIDJH>ah>Wn3pN3Wk\32E=`U6OD[W]7\F;dUh]ldPa2?0
A?j1gWB]o1;NGgS1C_ImJK`0H`WYedHINHEKjcN6R@a:;A3MDE\;jTH4G3^0SN=\
S?\M63[lOE38?l2`[K>Xg:nZI]Hmld5gNMMbic\eR@1j;A3MoBEg1CqTinL5>Z]`
E1V<<ffTP<ZHK]Q[8B>NCYE[`QjXLiPcbcT2N?AQZLTmIYck2eZZ=7GT3X40lZSn
^[^7QQ6nHAf;Q:eE1SbY=[Zj`F@acmbbQQ>?lYb0SDS0oVlHl732=@3T?oXOl6?n
^7S7QQ6;ZhT47p6BbI[M:g;=mM<hgUI:6GjTkSa2o^ao8D8NK<[koH;Lf^pkEHX=
eXA5XUIM6@fC<_4CQ<o3hZ1DS@6QDLi_XDkQTA1\eJaVNdfhbSJ?;Q>D3Y>kI>Mj
PakGPQ3LeXo8:m<0F>d<7bbB^]EPD7_i@Po]SIV`bJV0@9K@jY]BfLRd3G\kjlZO
PB>GPf@LeXob0<bFcpDD3^^_<n47E@V43Jec8_`fi<^O7kLC^\MN\OgbSLFj943O
7oSd=JSIK2?Smi563KD>aS[4]n3dHma??[dnX4^m3OBhloUE?GCNcRYUkCa@]fEA
J1mRW@_[o\=f>?]6GUDhjS34N13d`Ua??[VPd[fSpFSTa;R5hgOKQWN]giH]G;V8
7eHBgega@?7Nf:CMBP;5OWD0FM=@2Bo>KC6X736=4FC`B[h3Ahi[<7:`EBomo3=Y
KG0=KKiVH:7_D6PH:\CgGOGHD1XeORVVH8?=9B6i2F5XmOhHAhiJl7:`EgAH8H^p
fD?EgZBSibgjZn1;_KPFBI6h`OUO@5do`D2Scf:Y6[AnSTU2IWXiM3aD]DT`:ZBF
fea[:ik]ThEiZkAILcmlRXlXCIm9kj6L=D2M?N5jbfm6=KkaJJ2M?08;C>YC[Z`C
fgkY`i_oTh<iZkAI`4JB7:plP7;I<SJH<4lgA7_`];FCm=B8[mW8RQ3M=a75dA^8
[fLeG6UZk7bolS?i`4XBJSfl]OnXM[>LL5IBkU6RaSfnJqf_`Q=b`g>gKVX?8O6@
9SiZi^8^i:WVfZf^nXHa<h`iF7Ue6K9:afEIec:_oM@NHBf2G_@kgcmM_i9LZWX`
e>T_;iUgP_Tl^D[^>6`=m428\h\?>2?C4NZ[1JSfSN;N7Af=CMYkWPm[RW9LZWj`
7i24pmO?;`66BT<E`[k[7Z`g93d]eWS]L6C7eX0kk[G16XAFdak\[MHMI<DUO^RI
HQB]0mf`j3<E:E6E<08;Bd`DhTeCVLE@B>Jc6U0S=NNGMfGmDLQRW[>keHYRai7V
:GBKomT=4e<OGEGk908;BLRN4KYqOh=_kUTd<dc1M1N1LEd8NW_e3DKUFnbAA8l@
PBMOFDqT<DHUAK@?L0Z>CIH^^mQLMU`?7ClnT[f]0>UmoV:3EmeD[0Z5HM9KSonl
XHZNTLmTSN2fUSY01Flgg]0Pa4V<Q\kZQ:]j?56<0@a4Y@1eFYSf4n5`c3_85d`h
m?FVT@]TUH^1Und0oZagg]0E2c<T<qml4L>UoZc6gOS29NCZ_illYC88TJD@;0?H
GYT7a2M2@>;eCc]M^l1JbJ?<0W^CO;m_9JF_V:DBOX2`;Ze;8kFYReC8kE]f5B9H
GZg@A5VfM1PPPM_;TTYUeeG5d0aCgBmadGZ_BdD\OO2`;ZDh6a<`pG1_VS:JXhM4
mWcVYQb=^iV`:e?65=32nh1f^BID9P<m4PVDDEfhgP5SAZkUFSblTGadm`\lQf;B
7X54c7kcW9^SA`=VU0^VGo1Kh9cAlbIPGLKl[kemDS?ok\h7mab4BG^8_o\1HfBL
7X54cGmSAFDpo1Ai\UggJbj5b[kOX6MnNbBXQg8Q1OkGNO?K8bnm^k\?Q^IPmak>
j1:`21aZUXEJoJeKWRejmgoSFa[_S\03_okA?XM=l^f<fOf>4\IaL`Rj@iS_GcYb
PHf:J=_NHXKJo2RDlRCom@eAFa[_ElUH\WpTFdQKfSHM4mk;=kfKe;cc1?:^<gKM
F0VnanhWH[m4agGT46mLmAZSmfjoEVP4>j5TQJ1P_IZ=QRRJlKEPcTOTJlWf@_Vg
JjE?aZc_QV<^FN^E`UZmT=7>D10lNhbc>0ZTiWYT_mM=BfMJlKE_goeRKqHh1iB3
\81TS4U8o2<\4dXT\SjLddYV10H[CdZnCA\hVc_^\3ZH@RMA<L7mEZ:onPHm79fH
QG<TaJ7dHdA?kMf4fP_nFC6>G[H[cm^CDe0LkF`>mM6O`0[jGBX4];BoLAHRlKMH
6F<;Eh7dHdGNj<74pm]O^XE9G@kK4eP35lb:mNC`JRW7V_cblPWHQ50`i744ffgc
`NV[Rf^fQZfOnAYXimH9W9>bNhSmEkkFDZm4<SMQC7k843X>anW2^WE7YSbOZ8XC
J;GCV9dogo594\YZTm3TFB>nehgGgkkFDGoI[<JqM3KB7IFC5BERLH8SM81nM3cl
nVCT5`@98P7V1:8NX5N=fSmBc8N4Gc=A0V7RRO`dMg<W>?LfD\NJ?LG`]094e_qA
Cgd[>_1]R4FXJidQOWT=[Ck`FKXj[>p@HPd;cN;]OgInn?RgVLSH:Fadhgd7CoTf
GXXUI[FNjRM8nELf12B4_B<NT;JgV:=@N?XYK@j:YFAKJCAh<75b7j=^84J5VZg;
GYNSWf93Sa<_ll<n\M?Ue4OYSKP;VVC@jianKFd:Y3aKJCAA`]UBjq]0]nmLWc@P
?1Ya_@X<_N[njT_=lB>1`>Xmdge<D46FeVk@6iSXNT>\oHnCg?E>E3]9LQa?boBH
UlTNU[FVVJH\IRW7WORm9DUmnmb51^b9>5JTV7i4A?LNgEEV6a[>_3]m3Qc?_]BH
aHTNU[og:f2Sq`RXU^LYTGDVOdl0SlRGe<IZ5Y^S56@iEeI>^?BLPMVc?;[SOTSD
@SUO3S6IO6H>H`ni^7_I^07oI;4j4k>1kHdLiS?P@coW]8I>;c:ED3M`dh>K=InG
8kLQ_Jn0g^Ho0`:kE<_j@07@^;4j4oHMAgmqfVdOm:XnN?84C8MQOg@23OFdg`:W
5iA=cg1fo[=jAjO13REGVW@9S6b1c9=T38gCflJ5B92P2BCWcDPnnPX_MJcM`K@6
:k\TIgJbm=mK]gD?8UF2L\ER9AHRIjlX58LGf`C5_9WA2B^7cDPnc@PL]9q^RD`d
BkDYc04X1f[g`6HNSDk^XC:K5QdUCW_E6W\Z?_Mf]4Ob_J51cTMZRQnNFW\^bC14
UYCgdG]^^LXIgNEo4M0j8AR0\c:7C\0RLBaX9HMc7gTfBRW[ZNRYcS6JFHC^2TiD
U=@gdUY^^LXCG2UlVp@oLk9kI93S74UTJGcGO0IJZIc>9MbM4>ge5d6QhS=hfd@R
X@_]A9Wh^7lX5fBXJS@]4;VHK^@G<Z=bkSja@Cof7lU2]BSEVNke?hmnIXDcHV\L
o5G:cT23X;Km4jlXU;@;OX`H6C@G_Z=bkS;2A_SPpjBVZa^bNmJo7o=MkfHK^RjR
^W9[8_nS6=0j9mbTYT9WPXokAJfF>BLQ66e0hQoIQjNf7I9S]53^l1M?GB=g8GXe
46=>jb0Ic40J6S\=JFmVaN[S9DhJVMTn>nma9?o82j=a?n9:H53kA1M?G]SI?iYp
lmXf?BYanae?UD<5\5lnWNCi2elP[?OPhdDhM2hi]mO]d_@O3`G`UMn7`6JDED\9
l\3Fc><FTGoOPeA2BCS2Y7C;8hFJOJLCfd\nmJ<D?:3nLQdQ^5MFK`M>m6Be3D9f
lRKfO>;[TG0XPeA2<nbGX7pe3B;e]86\9^`HF0BkR;eU^31\TOl;V1S\>3]=I80A
9ZqGc\DA``YIO4J[IaWd6oi[Z`?ELlOmFPlbHi;m2cUA3X5<aI?c:5]7MP5BIH2W
TUGGegi1SZ^PD0hc_cgdeFSj`EX14f6dDS14H;5@=<1CFDfZ6nF:a@W7X@QNY[Zg
T`KG[YMFS`ePDH?c_cgAn@2Hhp<Pdj1DP?L8L=8ia=IVj_\^<]RdQAMmWkTZ=PC:
@PO6OWMHll<V9P_:hM^Xa56[4m<JS@XW][obd`@7l_1m`Hn\qLG9?IhqjcZ>^60q
<g44XVV]0R:oAMfGgeU8<KSaWc_UmK@SJYRGD1?TaJZfSKYlaO]j`c2ck0^Q]]ja
]J$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI222S(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;

//Function Block
`protected
J^]i]SQH5DT^<E[:jh666_OQdB79TD01jOH05jZ@T3K><FQ\Qmd>HZnoRbMB7WED
pQW0SCCllACBdQDfn7H<eTG;@KH0VT^8PpaRRDa99aSChEbFaT=d=VGeNNTW`DM1
g_0:>1K`R?LcS3P9<SR3`J1Gl^U7oapkG\NaDqB3mUVMH?MBnBN?KSe4<L:i8mb<
9`YC\9E?pMaDD64ZcCV5:KMUX9EjdJkWAo_nW]XimeWqS\Tj^WaOVB:Le_J:TYO;
QjGV7j_SPnkRSoqTkQdmYiGf=Xbl@HBSHhbn^JCD>PaXTB7:AcRp2fJQR?K?9QfY
cPXhidJ2RS<XOb<QMJ`ToN:VYR0q025=>;Xp[fiYZ6qH@kGnh2><EfnKPCiX;eXC
md1HaVZOmLQ7H___G5qmbPR@jK7WoN2b\Ta<XEQBe9K4Z0fX^0AD>2PH4J75l6E5
40lRWVMW]L5dSK5K0]8m@Q<WNJ:aoejmDcVNPbDGeU9fKCS7TiKk>Flag5iFa81I
T]9dI9oV?I?ccFNj0^8mcW\0N0Ja=eGmDcVZFV]aBpO[bVCQCcIDaPG\9fcYb9j]
mO69\agngD:a;=S`Xn?9@L_aP0R^h6G3I[SMial0I]OaPNVN9oLhoL:U5>I3^2A`
H3FhXKAX=C>aj\BS8@l76_lE=<1eC`0NdI@EgUQ029OfKEZN:TL`PQ:U5>bb85T[
p6U>[dc`4m?XbaBOQ9UYL?n0KRjMc>8BR]h\FdYSAa]];[DkKD^E42;VGba\\UYm
?6Ynnba0IO?9Kj?Pfj[<SA[Y>Mmgjc73Y>hD71=A3?FXNS0?QGA7UH6N\M@BKAYZ
o6_De6a38OQA5j?PfVPUk?YpdoTVjj]_bJ:KM3XU_;^KE0PM2:]M;P8_CiQ>]5lb
]06SnHPa9lbbcKCmRKld`EA2d>iKJQQKiJF`TZXHB53mR_2R?:n134lgQi40]>SN
kT0?dokiLKGlgg>PBYXZQE:KddfRjQ0di5cJTZXHo0MBP4plod3TQCcVi3O<lA`4
4daE<kOf7k=[[[]Y1>c85L4NH;NO4A^cUW_CaIjF4_E?G>1ll3@65nCnHjG@647l
ik\4eek5k5VJMRaN1>3B43\_F=WnVIOaG^=Hl4j=_Gc]G6>lV:Zf5oNnXdL@647S
68B[WqE8QOf]IU<j9Xb>2XZRPS2M`A9:f4TUAfBaPq0O\kh[?K?fQVLL8Zc0VT34
j0V<4^0NX?I:>MLJYdmlFfRN_lSS?4^^DQS=mGVbj`0F2FKjddBfLRd<LLEjlZOP
B>G<SaLU`ni:m70F>d<oblB^]EPD7_i@Po]hgc`bJV0@_K@jY]BG;id<LLC>[0`E
pYWLG7Ubgk1L^J[QTEdZQQ60H9LCGDke=g1d?6_C4a1K:kQlE:`6YSG2jEi1ZmTJ
nYAIXUnlW\1b3<PZZniWi@E8@8bA]@jcbg1nEVbb>im;Af0S6DmjmfHlQCaoG\TP
nY5P?mnZA\Mbe<PZZ:T`9RJq3Yakj]F7k:EXD=9GGa_BhDa3WeY;2L6@BlhACXXj
P00niZaFl7W^3;NK8jdjEMWJ30E^NC`OgdGD;5NDf45`_CH@o=]GK>LQ7ljULbQT
7=>b2d9RjI<`c60`TGEaWMnU3mN?]Ce=gTm?;5NDXB2OJlp[12M\k5Wf4h[[d85Z
3aG9CYMCkI;J5_IZQ06<I2SDR;A]EJ9o]KZGED^5a^^@ajF[6]QgXBZH4Tk\QT_\
5kmO?WZM1:jc4eQBQcnIjSNAaNc<6_nR?jV?5kMJ3aOja^\[Y?]PXdFHNb\\QT_T
V\P]GqonT;=SL_VL53F1\cGVJH8on=1?oBAA\A]5Z_TZ\;a0a00fUdL[IbHg]Da=
<>5l`7ojWY>VASoL\KobN_]1ck_hqFe0]E9QPZgj23PUAA]iaWBa4PakoOoWY72m
kB46iR]Zf\VoI>fnIYK>G85DE^h1oFYbQ0CRQ[SUCM]1fU:?G;_DV\NNSE;e8B2m
eMWX67HETQ:KcW?BBTY]l9E?T_h5PFYn1_CoD[SOaM]1f_jL6k>q@3C^:dafm9NX
2;HEVZYZ;30g2L_d\n@`FPKkP5=\mkkC;KbmVNT1\WeB@0lN6_MF@Ql`oXAQDL96
BV?2NijOR?ncmOWB;JA=NPDil9I=Fi;G`AoH\kLYSaDF6GDSc_eZ@\M:SXVJDLnQ
BV?2;ST_Onp:UVWH35_9TkE0Rd1=TNKe_[CnFZmEE:@Si>40BeoWXkJc7cUmC0N?
M`ckbYhfo;k:n0YnlF>o:[=>`6gB?SL\gk]W@LT4c[MHi4nO33>YYTjd2Xk?DGi9
b2079jjHobb:=YF[l:Io:M[>`6gbE8oLBp3:7GPB63bC1O@D<3EPBERSN>i5WlaD
`4cBPJ=EF?e>DEaN5<nA`XEimjc1V1O1Y\3H2UO9Y<2Sm\RDLCh8EfJNmL3N@JRE
VlAB>Pl;_:goMFB2]eYQaQ;RBgEB19M1;>3Vn=>95V2SakRDLCOY5J>9pPh2Pid8
nROMiLYffKWH_@mFhQ@2S<LAQ48Fb1V@kXiakTiIHKUqDj12iG9G>QXWm\P\jinC
5]L4=dlaJ3ZP@hGeE;[g4b;kO:c\K022=ERcgN=_0?\JDYJW?S]9TS9jTa>0UHY4
2XUg0f55iQO0;hE\@L30:fJInViQgeJ;5Oj`MN=U>?ihDlF_YS9:TSkjTa>09R?K
b^q]5\I>LcSFJL]oEIPdhJL`DG6\YYN;fo4=KR]bf]L>:YQSTSJJ=FZel5OY2hGY
:G=]UMf4\MV^^NcIWcQWdMMkCP>^?`AAWYnGKiOFXC\KKH_C5jZ]lXY89AR?]=P5
:_O]dYFC\4=^^:OIWcQCZi8]cpNjooc_300`;1olAVKKWhP=NWHeLCj<O6dban?:
0M;=U`helK3CkDnTX5G3;j9@70NfVo91fFcaaXMCZP=8]D1l2g4Go6]o3=dbZ\X<
4Gd;?COUBKUZj363BK3X[6I@e@NNDE;1C\cagbMCZPP>lL0KpgGND>M:T[`4kfW]
Lf5B8S=<YL2i_Po>KE>T49R<oQSY`HATd6CeiJj:`ZZ3R@JE8gjUH`8D;OYBg9`J
MR1Sk[eh6m24VE<76R>Fh_[jXEd]:nSobGj2an:iEXfJPiJcJgdUnc8>GOY`g9`J
MK0\3H6qJaa=LjF9_TjjR57IQji?HBOS00M@cT_FdfSJ52Yo92o3G^9;lG^QiK>m
Wg]Q>`T@Jl>f]<S<AECWnmCO6Cj\5^WY[QZM`MG:\fJYIJ[?3G1:UDYL=C;2M0RH
?Dd>c`2VJK;i3<o8AE5WnmCO\9[Bc7qK@0Gf]?EhZbBiWX=knH4@kNX>6EX6^AI7
cG0I0X6Eol\ioKXPP=719<oef<Bcd@dK_\d;dl52>SVPF=g]i9UfIqkhBWE=T1l2
C4n73kX@YV;GWAXnFM^;icGh;fKB^K4i]\abB9RNLSc^dni;h1?`hUk;e0WMkZLb
f>eRTnVC:Q8QRN@mBJ_<UInhkCK\m`Q:eDUA<=eM?c4=:gmG;f7`\ok]jC^MD6LR
6GeRTn_Fo[?1q42UffBTbNU<el??]2PUD?7EgXj3WSHb\J`CW:5Cj=5cB1=m5HZ:
aCBdmH`1l054B4e>fo;=>6Ke7ePLi?[NPhHLJXC]jS[nHF`I_feYOmoO^cF3Me:g
EIh9MDRg=k59T437mm;DF6ebEePLidC8MM6pRRKW1\GQmgW<PBAfRY01Z0@O[foF
4@BQ75\SGlK::]E^@:O5AbWDJ]d45l8q`=]2;m`hdXD:7ll=mn03UGa057TDIi][
SB7Hjmf1hG0Z\<SI8U0`=EEm<o2B21`l`ma[DoQbDbMfPkO8haL^g]Fk6bV;4nmC
XB1AZO<RTOLK=>kDSd>Rf<V7^h[:912Y`VnVJo=CD@8fPkO8Dl3\L`q6?>c5o4K^
`35lE;FdKh<oY3@C5`hB6G8eL@M]5<kE_51X?Rmfn:`=1Yh^fPf_3C86^6C]kVcZ
hld2FTZOe<4fmE?XahQ\=em6L@InB\>2@Y7TM]9eE\M;I6EZZ=6M34H6dS=3kbgZ
<d02FTZB<cJ84pge[lO88I_L<mkKoQTc]d?@H1[?o=GZoif0;93kSD7RE[TM8@dV
KZYAkHe:_fB;m2gC@VDm`F@b^0e5CbJU:c>\PlE?1WiP5Kk027V\Jg[hkDA;8U97
P273kAmC5=[;:Ug1;RVmFk@_Hke5Cbn@=L2eq4N7OAbOFhKeKEhGj`kkjW<4gj8D
MRR1AkbYhY3Z:g@@RSo25FhGNXgjEFQi]JhiT4Lhl36SNPnClJECMOd_\JBl@b2h
U[H2P1bY9bPa9O;NR1S9m[BnOk9bm^>fVHh2H4Fa@n6PZPX0mJECMG6c_ZRqd]EH
j\fEkkWfbmef2:lG0Gkgjh:l0C`Xe5Ti`U]@klcYITXc5e2C9Gk8[U;@V=9^d:4i
GH;]7]VfJ;X<5SmWG6U?Jk5G1I8U15XHG6?aS8gTR>lkFIVQON3f1Od;l=ZVd<nD
8Hc\7>COJ;X<<3<`Y^q9a[ODbod`KGhbO>N[je^c?YD:Lmk;QhCjJ\`Hg;AX7_X^
lH<Ae?6KXYIDS[EU`1^9bnWHhZC7[\V70E^f8RBQ\?Z0LE8<5=UPJfEabZjCClkm
GoePNBAh;k@MUj=e`2g9>MG7hYf762I70E^G_BWNkqS0S;\HG4E^]HC8mLDgN?c=
BDgjY;^Gd`CZ]NaZfajI@]\PT:a<GdcS6>IKMA;bW0SoQ=oQBghQh7TIaHPW<[9:
h[G2V]\g=HnZ2U?LO3`H10=97JkU6KG0N<m;5<Db3`Sd:M[QnUhLX2TIaH@FKaSn
q5AC3bS[0fdb:mHT8\MbMlgW8NGF^=hd[heaO0d6moMji?3Z;c3OgaK^dof7RLn=
L5@\:m]DFAPVjcGo2@II`\gqS=R`U13]XBIjM6ejnVS2nWl<3RR<aZTH_XA\Qj0U
7SH9ghh3oCO?k>kYp3a8dCRIEPGF@g9W;14\bgUJ_3WNMXcUW`;YX_9m:5kfGdEY
gCbIZG[K8LCkU8@9V3AVh>_mb0OXgP`<dGlMo6\A7DOfEa`d21;[0?he:0\MAg22
5a\i@ionGKF9B_@QN37EOV_cU0OZ=P`<dJUN2?Tq91MK3c[]248<h@X:8IX=cG^I
c:gnG;LMnE6CBNJ7RIRP56ag\`<KjNfBFW_i\4V59_i<n`dSKmOa9ZEOA:?_]jTZ
e:fG@I6GZE^3mCn7Fk;Zh0h0cVa_hCX]Wah4J4?d9Vh9R`2QKmkF9ZEOU48Mg=p6
Fnm_g]I2X0J>F3^3KU_F@]88Q^GOdd2>RbY7<He5eJ0_\g@ggh_6Qc6^XV1h6;d6
@>8ULgUbFHU9bO57iZlX`0QGQ8k1l6;BRf5MKi`cea=TWnYJ\\f;E9C3joAH6gW6
`=DeL@RbF3c9bO58O]:ZapV@ecJ<IKM2\ln;bF^LC1g8`5V_E264KKQjVFlB@3k_
@9=hOGZTJWZ:D2ToS][MJ]VPA;NnPOmGKPCN1a4PbJOo66>hfc4SXIij^9cHh6@n
BOKaISl<ID4hk0P`<UNMN?VeTV\nJgmG^2CN1aSPnN?<qDh2e2bNnFU6a?0TJi>D
QCDeENVPN7\Pa>bMj^ZkodiM`J:WHl=@;_J0JWkC5bM[HD4TWCd;DbZoNc`3Nc0^
Om0j?d2FZIkBG\bX0=A2jGIG1R2jA:8`;fV64VfjQZMI=D>ZVDdAdbZ;Mc`3N9bM
hJQqcfPV1b8EXQiIhAD0K6bGRLm\[]NXmQ<66m@WGKV@im3bVVCFfFkDa9d`bbCK
>[Ync[jDmKRLGBc\P72`?S@0oOgJK^\0ONSnlmeS>LAYDj=Aio:fb2QD2DNQF<7H
I[d^cPn]0KN2GBc8P72`6f:4f8qPEZR]c;WZc06nMNSQkfgCQ\RhW]nkMJTLRg8e
SXnYKKQh5kKk]9RMgRc1elInLl:PUPgn6mkj_E5M=R11BabW@eP_Wf]?L6^0R1]J
DHPjZ[l`:>:\PbFHI==?8]WgLM6P?JW36Gkj_RIM=R1DOD3CCp4A3MbIo=LI1`a@
ilOHB1oX2nJ=dLP2AA8m4df^fVG72Nka?QK5PHkNh[HM]lKm784j:1c7?jAf>_QZ
6:0f76[8[FMc?m]]OM7mce;3I0mC]2:2:[jhd0OM`1>7l@\mRZ4kP:07NAAf:_QZ
6:hlE`3=qi_RF7>LMR]n:TUjlIc`g:QN8nY61^oc=:IQ4WkN9>R\fjnF8GMLdjVF
F4m;7adR27FbAq`B_Z2b5cb=98?;3[KOkMUhUo>Rd^;D[n:eTJe6H8PKIk\^SM<C
>AJ[>^GP<ER`L?`9UOfkgdUjOm^Vm4XXd]CO5fD_Vabjm1@ed[HCFPIQU:bL37Ol
7[ShlT2?55C`SU`J6[@kSmUjDV^Vm4:I4?EQp_nfSBdlVI<@FfQIV\MdQURcFF^o
RGM3S0o?2:33lA1D?DE]CFb?T5SLWEbEa:fNY_NoP\0]X3bRGh1?i?Q<VPQpS;e>
9[_BB=RRaYMnX2@]HoDEmimF_\oZb5e?JT5mHnEO8j]6<G]IIWD5UnQg;<iZRjah
3n;2]?`KS;lAHdS5b4JE>ki[9IeFVL2V9c5<4B;5OJVaKd:R]jFI;ij3?jHXCj[K
3lPLI?jRSAd1HdS5eBITMGq??B21<YAUBN<_LmI3[<[gCQ82KdBL4DGng=ib8IJN
@PPSGXfgiNLeaJ3:\J:_O;4`SAiMhPGh?[mdF<FCGElg=hO=BU]0`:UI=lAkFIVQ
82RAIW@iWAc2dB`UC[FV:La4S7]MWXAN?^kdOB[CGElm3a8QWq>UPLFnhdLi>QW0
N4J3m?aRgVY808_Cqk:Tnm7ig?K78>A[fRn`5^ak;BlNQi>4hJC^AYcPH^E]oG0O
GVcR2ZbG1<;mmhQSok=o];;ga6S]NcJ`>dYB75Yh6>B]OS^1WbC\OT4Rk9UU=:19
R[eaLgZeJ6DR3>Qa8khF;S;@a6P08cJ`>Lc34bmp322Jf0j`E:@n3:_4<fA_Y><[
E?EWlhD1O?d3m2h:i_8?J]GMWfIc<Ra0h7<m6SZ9fBK>HoS8O[09L^WTV`WOP\0^
W441VaYXU9LdJHheLZX`a;@`b<>bX1UG7e1]^FaAdBW1H7o_k[9nL>K9V`WO:1<F
]RqR1iULnMY0e=j2Y\n2YBUU@[NdN1U7L0mSYC3=QgT3ZRO_<16e4jVJF]OIQW5f
RmlIXC7W_Yo4mI_OF98jeS;DXb8iLgDejQJJG=]h^Q[]G0HR`bjV9WT6H=TU]U:X
mGePXc6W3KODmVdO5C`jeS;9fL3`ZqfcA[U[cI6QX8Y2hj6`Q<=9FmLDVg?hn5im
6UANAhMRNQZLo=da;V@[FinGl@^4RWIQ2J6E=W=N?^Xo?95?1aXdMaK7bf0o>Ho4
7@dj@3GmB5LdMG\ZHEeXnJdBVAlPYK\Q4Z6I4LgNROXjAc5?1ai@iZGhq0J5FaDm
bHojUh1bDfe>fDh05mOW5>13hMNd8BH_hL:l@dZ5f[SBdZiSG?W1EkC?BCGVU17Z
GHVZk8?<\B\^@]5d_OhHAhJ[<7OI][omc3=YKGO_BKiVH:7^D6PH:\Ui\OGHD1Xn
ORVVH8;=dB\^@El?NBCpe9acO4V>cbfJg4Z=j;c<Y31B<a>KGlCKhYNVZHE`8RnZ
IiD89d5Cmg0eieq>o?KdbniEO6ThFjKI;VdOe:QhNdek=:_6fVU\Xo0LjA19f^7F
WJI9H6YjinHg<>ZQQkZ39Zm@\;5I\[l`d\a=IGF0H?h;;e11D<CXloD[dB65fDTJ
>4Pd`QJlmdIJOoXMQ7h3?H]D\m\I1J<`d\aXjoQQ>qRKgKmc6AaMXkgf;gLEDWF:
_6NjFJTQob3jg8OnbH0QD8lTmW]BZR\F<I@:aYYOQ0C7T:3LjRO1NGc]H0VK:1Ii
iOLAdED\D<SiGQW;PIJ^;HfgH[F5k<H1]g>V@E?Fc]]7CM3R^1K1^;cmW?VK:1?O
S4R4pi9VQmm@[NhgYan8F=A^jNAEFT@>@`N7B3PB`a@c=Olb_cMCmR2AYLemGdM[
_nFPX\U<kh2U>60jTXN;[UCG<24E[9?p[I1h7>D;C^B8Uajm7C:K95BNNCnQ;IFk
DDImj4iFjhVF94:ec2LLE_aCEA48[Bd[meG5E0RPRl]KUeZZE5\e?ikP;>;hW`cD
fc9RQG9Z;ZU@;QEJ^@dkZ2E@UJ7mJ]nXTe<6EK=:>lPKUe^ZE5\eRF>YJKq]?;?_
jL:leI]Z9\c8<d\Go7m4SEdQ5CmUVW1<0Sd7]]=[nTl3>K:ZKfj42GgNS4>DJCdg
XKAM7?F77FE^2?S:fH222S14P`F9lCD8\Z3[BBmf;`O]C5H;RjFKB>bVVK_cJZYg
?8kO7E;77:^^2?SS\kZV\qJ2bB0Z=5eDJ?5JSBQLI_fgE1i7oVVce5]_C33PWZb=
>LZiNAKYdBTi:^^Z`7iSe78YK]2=T05ZTkob]79SU^falcD^@kWRZlGedH:MQ7A;
PXhL=S@[j?4cPFF?>8BD6j5YL12Sh5FZ`;obAC9SU^\^c1fnq46]0MeAlKTlRgOS
LoDH;U^I_>C=gQ0N4a4HQ]HC;NDBm0KJnSDQZk9C>GlWd2SQfA\[6>cO[E3h0j:Y
BRRgLI<fSOEZRERSHJ3<EN>ClHHaOYbN=Kd?@lmM[d4iQe[6lg\hI>KBnW3X\j:b
ARRgL4Zd_blq1o`BlNL?GSX59PPg8=U9AU`VUhNddC2HmXiLGeR0kFhdK9ck99MO
BY1^I?PR24`M?Hj<g@Nd_0_9h_0W[Ca0KDjlGahQ71gf;9@cn3RZ]];\P]9538MP
33@=_=[80<:chHY1gK[oU0LOh_i5[Ca0NN@?AGp?aGPnmmRNn2c8\eJeh>3:@oL^
m?4Yci@`H<jV=F>1c[1fn[`M>6lj<lSfJ7Y\;>mj\PI3iSjFA0HBmKG@CU@:gmDb
cfhglD^nNR:d?=0m;^a3LWY06N8ZiBQi?J^i6nhP\Df3KnRmA7EBm9h@CU@gR8eL
9pHT0260BYYP\YTi68>k^Z?cLC;d]SoJJZi]Y^f724m1Q[Q>qDE\JCGk?]1Vc`KB
fO_WGeBl6;nh9Tj]PF81SW;WcXoJdm62nLe2a^<D=XKc5VffPm6WU=_VG3KOBAbl
R\GmTlibRO0RR9mCZYCUM9EPjgQPRfDee__3:jN?m3Z;R3b^KA6SU=X6G>K[\AbK
R\GmTLF?T_5p[YIcD53QbRAZmYP0b[48Si^OP2fBcCJkkikS^i_mcNm1^WRiaDgA
f2oFWUigN4T]8=5V5PAbfmGAOg_:<\b]Oo?CJZ\a`E<FCd_NIF_ggfIFnM8mQA`B
MFQe9g]6<j:Md=7i5^VNGma]Og\5<\b]7LM4?Bqh\3SZ4A`@:k8JXH8^^:N98<oD
4YZaEO2QJSB<LJb4bL@UM>YMGQbUFnb?khA8hBieRR3Qckj@F:=Bcbea31IAWhKQ
e\nnHL[9\PVF[J=d^46a8UO6S_QI_4FO:9;@e[XdR7?QZbn^FlDBc:4a31IcYZ@0
7q`SP_1LK>bJF76h=`JLhWMOJ9QGW3OT5JdEC>cF0_=D53E@;=9d_?4:>QAcg1?6
d\QYX6aGafHNBSSN5An_JZ9dMjh`p5i1jB9p0WCQKIC$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI22H(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
Cdc7cSQd5DT^<>\h5bMK;8^Y\eSk?J?O:2?_kIf^1o4d211:mc92`e7AafH4PhYn
j2iMneFSB;\khfWpN8c39_RhS;3K:UG1\5c4E\5V:oW10RC;Gcc?BDkI^3_AdS70
\5J5L3Bgq@LYL?ChX8NIDl3C6O>fWhnL[W2VQUiMImFXW;KT]MU\P7L]>ma9nSf;
`WdebU<W:QQB`Imp`AL6c1p948J1ZTVfm2Ie6kUE6Qh:CnL7ZLG`@n[K6p4@XdN3
>[`Di08j@J:j9=1e0MWCg4K9Lfi6qXM8G>CeBl\eN1V_1f0aKj5c;C=>]7Ea`pm;
XLdi3qOTQ9SnpW<A=W_aHCKUTnH0jQaL\kb`\M@NHN9nXWhFcjlnd2K1XTOV_[if
VNG2RELGhaP\NW[nk4Fg9XJJXk5Bo;T5eC1Y7RB3ocfD4jhPHf=UFXSIRnCXXRGn
W47qg>R9bMMD]@KXQZ;9IOKGalg]03Sn6adkk^=BOIkN<lT_jOHJKN4]3MkaA>VY
m^k1gBKehPS0L@P`oIk]RWmLfgT\`7hgeD8la^jX5N4Ldj?6NVOmDBMA_]pC@fVE
<G6De=linfhgf;a[>of4UiS>1^7lP^]MHX71de<7DQ\0Ok31Q^21==Y]kGdCWnK9
C40RJD86Oo9Dj;2N9oingPjOM=hfPXR2:aWlZ4h6=S2Vd:NQSqenk\36_ech<OPD
EfO1pm5Vl=o8m4U3[alT;N`H0b:P?dQ?Rn9g9fNIK52d=]ge^[W?MZ\S1]NFYUF2
D8VYgmNk<TjlWZ^7hYJC97A\bHYqU556RbO9n]]n5gF`W?Z2jdlL=?AVhgOU5gBF
00cJ7\aP>kfHdkjP1jnHOcL;[fU@U6^W62H[V2hKZoc9Q_MTiW=RY[61KiFh?gcR
BBA5L3Y7oJigF7kP<7piG_XDeJKbIGi?^?bgX_2ECS4MSHk?[2Vk<\>53IKYFS=`
iPMa>3KWFiV]>F?@CdmiQmacd7YMIV2jcUmO;_]=AcHhIC?6BSPo<E@D_1WkgcDM
^A9Q5Q58`pB37i@BP\PWj[ON=DndSG2^FN0_`?fTMZX``\LOT8KTPo6Pc<oMY3jj
OcGdl3_eDSBM20;3<0Je9V>MgRb:GlEHQlDGQkg3?62`GW@Ci]lbAc<]]U1jc`lh
qYm@TM5R?GY5SAiL;G8QVC>R`mKIoeT1SYZa\KNB2TSQZVJh8Pc`HS7AlhLC=8Ne
5Y?2<iQL3:X<:Cf48XoN?Mcq0aGV36eUEVWfK0LDD`7FYe`TUd?IeoL5H4;SoY\>
G=P[Sm[]Y=GYWe?OZ04ZUP_U0d3=UJ73`V:]Y]3Z\@h3LDoW7`@S@97@o4F]6fKi
iB]I?1JP\e;4jEpI^bbcM:^FEoUNG5GV=0CRb3BSC7h4@5h@9XY]OGdhRb?^0a8M
`ZYF9WB[>3JP<S9I`2@_ZSnUEQSddPX>h`W=k`nUKGGQQ\619_Oo^CU7KLoRiGW>
P2;7bpYUWm0?kefJ>K;FeLOdk]=eRZP>Xc:INbogW>TP@;1belDNFQKd<NA:m]XJ
JnTfS?pCk0nfhN5=WcSGC[h`BHc0SY_GZfeh4ke<gnVb4YBUflO3ILDAe^K5aRR4
Ug53^^2CMWWY>giKY7OWTT49WY?0V1Ug7gM_[;JOgnV6DGA<mhkObIHHJMZUgp>_
;=TNdQ5i0V_lMi@P0oBl=_Qh6PM\S3I0eMaa]>3^9@D^[Q5XYfXlbT`:Y;OD0;>H
<G2ELioXMne0J0_=BHl8q[nd`ZLJ[NGhg5Oc>?0So4b9eJnG7Rn3RODe[ZMZHR^0
IXb?YX0\D<0lMRP@\f\hQ[cadA;\B9?dDHlUi3?olH;WRg6flDm1P@D1Nk4OiYkT
gfC4PX9b?Ehq81Mj=5[f[IaA6NeB``?<\^lA<QFXLDA^nMXl3kc9d=mKR?5dhf4Y
]7A5NY5Imkni8ZTWoni39\K=jI9A16Lf4@j94[Y[dAZgHM?DEUaVhSE\87FD6[LO
B^pFMf]A>4dG[7IgQRAjHNfYfg3TF6FE^7YgIGhXISVi8nL=VS2Zg>^A85EocnSO
kn`Fh2X>ddb?^^l:4D7IDF@SgTj@GX?_3g3EImC6268TG@RdV_HklR\B9p_6KoAG
bcV8bG7U>\lZgP1=99^S6c5_MUF3:gPJSLG=]jPa<>:_cc]NjVK4ZMZd:A_EPRbO
]BMeJLi\TL^E?nMbp_BHO?Rp622NWDV$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI22HP(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
eQdKHSQH5DT^<jfY4oAVThMb>UlQRCS9qndiBi?I2UQlAn:4T0Xl4fdhS<<QE:;c
BL:ZCPIq[H9lfIm@<2dfOlB=mId6C_\fiN?XjWEa]OK^j]NnR<Qm`k[BChjWiJ1A
=Gfp9IFfLmqOB5<=>PT^8n5@cfB:nY\oI;:62G34mC_1@q72Sd5IZCA[A[ZVjG7W
FW]YOJceh49F48EdqhdJbaERigWL2eJSL7ob`F<ffG;N\XAlZpV8=j5cAqb^bYOd
g\KW\2EJdeGTl;fWIiP1m8XK>DVh:HIg5GbdWcd@CJhbKpWXFCD1p5i5U:Bg8fLD
9hJ3d`0]GZVjBHl^SR7cGi3S@_c6N]H6idg\lK1\k26:8^=P@__Cg5:=;3D0jl`g
D>GKM9TfkiSKO=CBQ1kJ;53SRg3n4RQ:1f[HN@`]^?CqBU@nB\dZT1QX\3V>Og:G
R2]h6SF0YEc=PL=Zm[6FIDK=fe4`C38RI5>5=<BR=QSNB]Q5Ueh611CCP9MQE442
6k=99XQU=LG^DLT?[ZVC[?iUdfc`c[CDE6qUkA0oRV0_mSlemm^SB>oYXon`kX@K
l3B:]fED85J[UQn02mLjDZaNlH?0W_W_0QlUZa1Tmlfbf]PnQK@X0>IH;i4Z]U72
\ka`]]TR]^P@CKTEQ8b<0\SOIpoFohc13Y1SUEGUmmKD`hbZX_OR5N0KHVc=ZNbf
i4j12G7<]hJcMkKFHI=X`M7S1`o@lD]=MJcR:NVD\fIL>^2oqVj_Pc5\eO9PCb2:
LbDKD8=CjjhC=h\J:FX3eEf0;I<:C^S8a7ik?V=>CIVTldSH\VbU`kU=Ld^U__HH
]<3ZJShc:VDD;f6mThXBR0U1ETTCWZbO]JW\EJTpQfTPM89c3=>jDCMOnTB:<Z:H
A]7fcQ01<X9C;E3Y9<:DIflN1a[84>R<b4TA69[[Q>REFFb6;=ZKlGj4SEBMLJjE
aPQM<\P>FX7f;B7co5g;YJcb46LaK5qbRVMbfZZa67hZ@iS8B:53J<l\5102`WUo
=:C2C7V<3Sj\P7]dSgQfDPJ^@FGnD2bbP:QC^0EG6kOKNhW9g0@0ZS;`O7m14N?h
=;J\\>UPK:P;YhC7]MR?4p0nIPVOVQ?IQSo>n]Q`akoEb7;I`85?e`AUK4N3jGoo
cSa\>23g7A>VhkDP^4He:U01@0mmQinIL@f4Xk]OJeLhqYINlO<Jg:06IN5]YYRS
@S>ViAa5J9I]ZOW29pPA0AfUN`7K7lYcg>[^GO<gEbiYOBYLh]d8k^iT>K43Odh`
iZJ0@6Eg=XWF?L9O;FPffjmOKofK8?2`GEg?U0R529LoPMn`<BO8IeToejOaN[[e
`7]6GWcAp>7SIH;7MMlg:o;\5gX9?O12072Lo``]W@^NbTQ2^nbPo<Zb;BkX\>AE
WZn90WfZ:>Z=MH;]9Dl]`7JKKIBJ60RoSl28D2F7[0^=C5YKX6N`_5kBo;EYmN>q
U:DIV5RU=GWlcA8ZloXLlBmS=\cS]]f;8P?6X2L9fbOh;OKRJ_NJ<RUfO[4QAJ3j
U?jff^V;?]QhUVTaJ6?9QjlIl\62aRaY:P_I11Y76;;IB@nfD[egQBq7ZgNlmNdl
4L7j97?X_XWBJce1U=RBF3;g?PG`Jn7nQd8[T5hlIL>aek=KLmD8eiM7WBR5eEH?
6eFM5IDDDfb=hqGOl3OT7YA`@lIB@i9P66__]Ih2MEklgbA9\UbZ7fAbUgU\dnEU
QeNe2aOJNqE4oN1leW@D08XPegocKbeKc;Z<EHi54_TJb8WfWAYL3dYo@OO?Ad?J
]VD;?ShToLEhUi^n^RGBnPi7?UD`Ll3>Wgi9^lXN[SEJR78WRa1K\leG\:oCGmo<
q?KGMY]<Ken1Z:3^:\abPOmnM8`K9GE9Og[;T<3@n5O:j1K`4g1L0]imXIdUfID_
o?O2e@M@`VE?jIEV6L?^R<?W9l`UNF2QQb[FT?mX8gkAOf@l6\OjI56qI=1@jh8I
V;I7hA]CSEYaANNBaA9:B9meJjgINJ0BkK^P3H3nj`S^TIf@RL\=2YUmI47<Kl\G
O;IBPLSE\<Y=G39>KiGJ=FNZAjZlLVci\5_^Y5?V]0TQinpL[f?TcQW?5ETiC`LH
bmoON?1ADcGgOI=\?ef9Y`oC9jUd>?@:Y]X6NPH5SEi@7QFLPj[M:;Xn5MMH4N[?
Tj5Saq_O]WjRqhT`jDoK$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI22HT(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
64L^QSQV5DT^<LaaiPCD6L2o=NiRIGAFH_BKEC\^TS>lJIqobJjTWQ]Q7i\S>SNj
VBk\ZCG<OkQ@WDDNN^KpkNWAA?4G7fmnO3OdPd^J_ndl6i9=\FNLdb>?lTXg0R<j
80j:iJDehMC7]FNXBjhJ^dI3ebP;p`OdSnDqMO5V4i>[D`S0JHGeiX8W[^geIYXT
eXFPX0p>6M3W:3@W:`hUQ0=EdIWm:O\HDSc[F>RWBpb0OLILLgk=O<JYAk>Ceff`
G]Y4_6kP_KqLoP4VBm1QG[Ne:@@cmpAb=e]gMqLob`g<p\[Ba43adUWbgnX1bSN?
<I99fCSGD`Z0@lPAajVd]Zn9:QW2BTSZjo[PbAW4cjJ86\O6J1Kg7@m]g^_j_5O[
mF:6Q3WC\EEm\SP3QZJ]B7aeQ42Kc^Jo`>_pXY2eUfNEbO42VQ8NW<D^eWeGb?WY
`=DF1YJ_MnP@HJeR4YRc=eHR6<R;CY;n]?ZKXLFVCOXP9O^RXHRREK`T3BoSa4`o
c;:AcYJVmNLTC1SVb1l@860\l5pP<dWTT29LGCFH@TSf8M94o28l@Nnd=1d`I94R
]>;FP`OHUOc;Z96`8lh_BA[Hhc9S9pGBhR_=b=[J0VCOXIj6@4FUa5?lj@20?We4
o^g=25:0_7iO0TDPS\7RmW^ILiA]?HG?^O@LZN>oU9WDFOd2@D=iooZb<SbmF>h4
`mKhC\kjn]GT^E5bRnV5q[6;F;6CmM8FQJ7CO=[njdMOFE\3jVl8l55i=Q;3H5WH
T<h24:5Q>o@3SFKBfMDgL[\\lbc_kbO9L7eRMGPKAS0pXgG<Ze^kjQo?DU51[kQQ
mdiCa]EECoOK5OiL0KDg>12A1ek7j_d?O`Zj=BVWFYmYX<T;84;:obV50:R>3KLG
RX4MBDSYlfc9IOKdcPEo4dNB5fTPk\cbJmp\HKH@@^Mn5`^>GlJJl??_dU=KLY9T
I[:lUi53bMMJeU4:`4j\APqF[<Y<gijbFR_NBH`Z[Mf:`46j?U`KOE@h[WPB;fH8
Cd:Lb\1mP2@gg\Q9^YHPOBQF1QCOGP30FZCL0Ha6^MhbhGMIT=`XKofi[Ybk@O?E
X`D]f_jRK[@QmqeM;AHhTCSZc8ZLSQYfI>X1lAa2IWHV0DPh>BAO<HkREh9`nb]5
1[8UUbYDM:3:h1eRf<8gPNVZF8\Q[ZZ7XR2D4Z\`J=DTI==h>9h7ReDYAK1CJ32=
2U_Cq4e`kE_fkgb[58;]KX6H3\JSS@X6U?aeNQPJd\m<nfUPL5Ql`kVR1k8B`fGo
0Ok5l4ACDmRY[EbkEEU^;lAJkd[pMIZ[EAcZP`PU58QCFgEkV8>KSRMMikS>NMN[
JC1oS:M3ol7akW11@IWF@YY43:bPMN^B6i0iO`0nVdOEPbnU<G1`EcCTo><MLM<=
TmSMK<jOE5[?Z7::QmpCP`\c??`jfYLleSHBHfQjQY]mMe\\VH=0ODXJURmiZFmo
Wl_@jAA9KNe8W5Bja9LC1]ZbJY@UfFaf3LN?k\J\I=`NMh2<j[IlO0^kRKV:ZVJa
=bbH:>1FApQbT=KLfHC\j]9oUKBG:afPgGL`6h6Ae;Q]8CkCkfFNaR2aART_I9aQ
CYDWn2c0NmQ4];E7:bec862en4CH`j?>cmo`EgmU1J3]LLhdXN3c3EX`\5o`1IbM
pRScM`B7<D6T6Bkc?2DnRNOcaDDGff3n\5aY6IIF=O:7=iF4M3al>m6VP5ilmhA[
nRc^MXW1cRXDi1PBM`^HS8:pF:JfWYDVhgjViMX>0e:GTEWRQ0GV5XWHmc`[JjhV
TZ;Oa`@D3lTjR=iJ91STFbI^F3iHll2kS[1a\gEV8CUF;BeAPW<4Ac>^0c3;14Zn
fiL\`S6FDnQfbLp@IIb?D6JCL7N9l=Z;BUldj?ocWdT4]4_n=gf5H6G[B[S`aUpD
<YnQgl_In[I7BdCF3lNW6VQRY5:d`94;TH<Fl3KTmWOjV2Zk>KXX7B53YAB5dKSD
9o;bV<L16R@olGchfb]<4_SeY4aIoaUBTeR0ZB8lng_a;WoHdiCP2qjLkChP4B6W
2G4EVg?j;TRDkMc4i?<n6?SYAK0Fo_cJAXCV[Ad[IZ[QVfTa\m1W2@jn^TTal24W
PD=B7Va@;\<FRQ^Z]7JDSQZY551>HgTo@ddJC856PM9ip4IDXdF?YGWcnkH]Hm06
bX`eVogFdK7e@SR3lRXifb[P^GPcm2>\R88NG44eRRWac4SFIj;[iFW`YAIj4k96
V;XqScW^kCqfN]`ON165\XZNnP6SWd:l1cYE9mfen_a\SWc:fCKF4OaOH3k@WT9K
Ck9mo;if>\;`H@qQ1bB2o1$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OAI22S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protected
M3IVVSQH5DT^<AIK0RKKn3XLIBnU[EAJVb;RM7jleX==I2Yneof5CZJ9=_9p37[B
R[JHHn>GQ<f_QWk\S9YcF`O_gDD5[FDQZFXT:1:9g7AVK1@IB8OjJ5:OFPhR3iJp
Ra4S_R7eN8cD^PY_^bi_co=iZ_]cPG_Y<PU7n`RoaGZGUX5@8QBOBmIB1gMao:h\
I4pgT>Ha1pN2See[ImGR<E8g95>9U@dP78Y91[N`i:Z3pX>T0OTCDNMT\jOnUM;`
480a1F@nNGn;laOp=7`02@;o2??MYO@6l`1V]eill_8FVBWAp]hfb`7YqFJ<HD1p
;C9^:o[i[B\X8e?@U0SgG12dRPSVf[a?8Nf8c2XUooKJaOHZ^PJJ0nL^]`^eDj05
;2iLGd1j>B=C22]ER\KlCmogJhDU5\D\6NVeE_?[@CH_KRJQT8j:NCq4G?^d^`3]
l2lA^5K[OLkmo?1_TPD@6Y6:_3PdGKA3RJ5jW[bFl@k4@n4K8DA;KTJ4;1<;bi`Z
l9Ih:D9Y>X[FB>Eo`b4;I5eW_nCiK`^4]ZX=7kTk`PEB1pJ@jhd1MWF7U\`_`nE4
[HKD2be=_]PBQYHaK7m3aYSMA@V1NiYkO=6Y1<cBe\<\T;J5AHkLLUY:dhT^FS?;
[JoC:W4>h3ZHAF1aFg7;l8A7YPYe]Z=HXcflpT=]YI4J7RHEQELP8PfB;Kn6CdPV
`B<4^<RUpI^bicYa6b\od@J?SYdAoi>^m`d1^9kj2>Q4G=\^?bYc<Fmi;RBcL32:
i5PIS5h9@I1GUYPnh0S?;HH1=?ZX\VNq_D]<:WhEQYjgFD`LnK4:;6`^72F4g==`
mISTFUY8;bXm[dL@V8GH^XP1LM0PHf6<_>kQh0F_57K5Rf@gDV_k9Th5R6^H4a\?
gIY5N5S3CnD9m]1MD`<8^VqQM2E9_YoO\``Rb=g8aC7`Z@F_WBKj3Z81mSKD^RHV
R=Z2KCF:<3]hAe^YdSf;o_]Q[j^=0h^^2Qol?^_<V6QZ5oaQmQDYlHX<m`Ebe8lZ
mJFRl\fmP4aB`qRo18eP8S:l>bV_Y6gMnLW3d[kOaSl1k=_j0P<]dfAhcNd1kl3L
QmJPc2e4@NVnCXRdRmQn02`;AZR8WG?RTk:MFEhFfaB7ND1j:;`>8SN=[AV_GfaF
I4=`p\f1ca><amYi[_fB[]>4HG7dHA^5M[Pn;jb@bGINV>O8m>j[oaEnI_`3aPXZ
nbXk]\H=C:WB04UJ572IF@m:X19p5D=;:DXbABSl1dgon:hFI716@Ue9IIcK3NIU
^X6FdKUUGccY46<2ThLannocOe\BVd;q5:ZNWCl8glJXb@8h6]oO]>?gLF5D]2gM
QCRO>389=b0foXZeUZFBaAN:kfX<mP>S5l813;UD0O6JOeC]a0X^RaTCK[?mo6mD
EC2J3;Ve06CV[;VkTkR?MKq>]5m5=[iWb^UKQaOT;13XN6Sahg2JhONR7@i?1_Mf
k8GR\Y?YRB2mk;n3OZb8njE>Q:bG2n:gbZW\5camhJ_mYI8nGVfA1Rk\7=ma9`nA
fdcK@`E\9Qoeep6OBC0h;2V<_e?]L<lb8a71[@2DPo]C<O`h`=XG3>M600I4KY7E
Vo?eOhcmUBf]L^61RHKF2AOdREj?OmZBS6V\@m<oH4PdVAeh0101Q:gCLY^Q<hHO
SWV0pSchULa0o>UUOk3m8LYi7dLVhmDTV82[0Z>MHIo5l:i<U@B1ef`S@ViPmWXb
4VoC[Sa`@0^>K0c0S`lDRiZ^KU?pE0bmIFM\MD;SCHOJBiX2<Nh62UKVCQEoONV2
Q97;I2YG7AZ3?1Z>pa9\O;ZD`W`]DL\ad32VaZS9OAd77`bR0kj:lShB`@HW8c\D
\3JBM3VJl3?V:\3MOa^^MP6ZU`7VVOHgQDc1P69^d1d?l4Ok8=jM`9g3RjHC>Hom
hTbCAl9q29=@Z]g:IEcCjc0W\^S4J?`fWFQYCk]dGWfEb=VcQbX5I4LOjnDY9_\P
XfhhJ]S82?>8Nm91jn0\n5iKJ]H2>2][fkGgSnPogWAd8<_MTeib;335HH]S96pA
\k^?2Tah`6Wg]k?Nj=j7[1BHa60iFdij`Xde@7792mnXBMIK8cZ8oXWgi^XKXQgA
RjFWAb33J5AL_W`eO]KoS`C^A5e[N:9m`e^jHNSR<XPa_]i<=U9kWqMiL5PHC8Hh
\7de?NDQ<_OkX56^E:0=WN_VW3_IbVk^VX746c?ZJjj8Q__28cI^lIMPKWUVl1:Z
Z_1OiTiS2n\Qp]RlhEophPKM2OKW4i5lgYghCnmVm<]h4mC:n<LIadkSG;5hOeIb
qAgR0\<O$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR2(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
2O`K0SQH5DT^<Vd1]YefXRJ`:UWR;CAaX@Lc[M3oPLNgEf0]jClk]dDmFIC5JMDn
`JhaJe2fWgpC^7@`dUe0LMddZb_Em[>Zd;3T6=lFeSpNNK3FMH7[Z1;4_=fOWP05
:TEjmCg?Ul1q4gciX=p:95L\[l4k6FD55D6j3U9j5>1jn[TeIjZqb]l9`fjp@HFT
9mpLA;\U1XoMjD3JVom7d^1J[gITfi2Q2_Z7JfjXcJ50QnielokVm^DRgY=p?GE0
L1lL[E9KCQ6=>dgS4mV@eNPWYdS=bb@1GFDYk1IfW4fmQW8<RSn58naS\O<<?T_V
X^B\?GT8REkIYL<p4@oiPSBkVKno1eW]>d8EHl2iJOMW6W\06BRQomN^I\4[=blH
^7kHPMa2KAZ_>?R24[eBhfCY<`JiHCm^61Xp\Lfn2Zl$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR2B1(O, I1, B1);
   output O;
   input I1, B1;

//Function Block
`protected
ZY<RdSQV5DT^<Ka:Va3HglT:Y9apCYU<O5[TZ=9Ra`lMD`:BNT8eYQ\[AX]oP_lH
bB\p\9aj3>MeiO^G6hM_BZ;>9Uc>L[<k67`qUQ6n60qf`=_:D3j\INOI0aTQCh2U
@BGDo;8DjNQpBfgIgB@1Z2Pd:O5U`jo6RCd09d8pi>oPPj<qM[<Tj`p>flGn2[L[
j4<bEmjC^LCE?@<n`f1L8V]hWTZn<qoCSnGQPZZ`IkO4U8nifjH4B;1dIYZJF>UB
[12h5BmSSOUOd<n45ZQ]4\J:SkAJ=GodJNlBJdNYddU[=CidgqDNCR@R;lmRA9<`
DU`RTJgHaDc4LKHca9H2oQnkGkPl=8L<VWT_C55i?Nbjb;=>j^0d8[7G^]WV8EGl
H^ZV0E9k:q^1c_PHS$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR2B1P(O, I1, B1);
   output O;
   input I1, B1;

//Function Block
`protected
ng=ZRSQ:5DT^<kPHkdZS8HkPf9GlVS@UmOHnf`5Op>IH;6`RCF6?@\7c9\P:DPN]
VpIEa[gEce8RV>L[?R;i5ULmBc_[_g<Z`9ZCMo7YUpjWi:D2q]PdPf:YRZI4\D==
3fF^9AAA3eG5>6<b8qSXQQihOZM]h2>k99T@[T:aZ?MCfpAfZS?VYnlA7Bc=]L_8
m9F7J]m?WFQbBG[^X\V:NF`W6aWej5^hHGp4JTYbS;p:D5AZ^p20HfU`J1TUV^:[
lMjcM5m^3P656CIH]jU\UBWTCdRgmIfUVg9MSEM9k2m^f5lA?R27m0k?1N`^NDYM
F6Sk7qUeU\X90d?M7^WIPIPHHgHgA;bW]`[CS8Z`S1oTIRT97^S7af?IP9_:he[H
jR01ieeGO3eS_H_l3fC@KF7Q>5oGIp=HZoJD3$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR2B1S(O, I1, B1);
   output O;
   input I1, B1;

//Function Block
`protected
EV1E2SQ:5DT^<KLKNKD?<IP[eoXcRU?_\anLlM6\aFd4\K8bo;6B76pG:LOY[RT0
Ml^1fZoI=MDXD27DA11l2QjYZO\:4]UL@iL2>\HW0Bd1X=EYBkSpY[iU<`Qcb3lG
6Y1k56jY1JE=WjCoEGLMTH5Yd_ZinmD?2ZX`dgdHII;Oq2cb]::p;\=fHYfI42ff
5G?nD?od1Ee\\bN;lm33p5d?dI;6]=R`j\I=B?_N=`J0>259qAPK4o=3pld?e=@p
SiD;<:H?ohICU=Vj\43`02l9T47OOioX1?YiTASdAb?IS>7[^k3AABK:lj\8D0ao
S;o9U]>nYL[JK9Agi[DpETQ_U=L:DPRPGZAUPdk[=7XO=23EGDdcJ7CJZ>DV>MLH
XTj=d<h;5eANkc5LZ0<kE4H8admjmMHlj?MRfRTpTbfbhZl$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR2B1T(O, I1, B1);
   output O;
   input I1, B1;

//Function Block
`protected
\`LefSQ:5DT^<Y^Y3f]`\Wa8JgB7>TmVA5m56l`5DD8T:DOMUfZeTkPKHaO<JKWG
aGAp_^R4QFiD[A6mA8j?QhlM2<GJ2f>W@PC0][f]lYp@IN3lgN5gcDQJC:;5G8U6
LqGb<KQOpS1O`>m]GYYIP9nYU7Q@S[_JiCPlgJMfWp>8KC2PMom9iRJiRAc:gI3V
HeAhVp7B;EKDYphfe1mGq_>S?YIRRFoWF;TkO25?4TX5WS;fGX:6kjFSkH6`Af1B
YUghFoE@3WIRnZjGN=e>T_PXc@_LL1L9Cm1]^9XRpc=2WRk5ac?R>3Kokn@fGaR?
GKK\ic1QDlP0U:l\28aDXGA1ZQQR0C^h@j_P89LSJ4@KLQ<JfeY@eJPb[@;1^\fC
qfTo@K^7$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR2P(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
=>`n>SQ:5DT^<h=`7m:6inq0CO^=dl@oL?O>JgNgRkC_OY:CiKZRXd09@W^08R0R
f]<dkDfHX8_Voh^`0ZEgkck]1;hC2p18S\C[ZjaPb_aGiZb1i=UZhZV@@@BA08YV
_fh0PLih3Oo`TFj@iP3SJ1:7ZAg]ELqDY`0X=q5_F4DZAJO26ZLZ8PAPIb@D:ZYi
9MO80NqA>D4>`5p`Wih@>pUTI8[G_969nXIn^PJL?b6@eiO_2ehGL7=XJeAG3KMO
l\4X>HkLLXWHa>hZXaRD84UlKD]KZXhn:>EUd>kZipN9J0AIB_;n]TY1^ZFDnDm6
N]pm4W0ENZlg?UCk?F2E[T>?@H22BdX3Y98OE?GV55_PBXH=_mJohc@m73=9:o75
EG0mdoXkj47^T9Y:758G;=qEWPFg`S$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR2S(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
[93GRSQd5DT^<Z`:[j`2KB45m[gCAh0^h7hp\lY=oo4I;;?k:TUOMPeOB\_HL<0c
XTMfCfEd<8DYEm;XDl=7q=T^=27De=TLS?j<G@g[;i@0>9;VX874`E0hO7nN138_
lilFeV5QP1kc2X5`428k^pcAMK9Lp6nUhc0`>mH1__`]ji`SkG[\n\\\WnggDpd6
7[c:9qO[Qc^HqdfJhVcM04bH95:?o2nJB7an7I=LPgK9=fShEh0];]Ad[J7i_9hB
dBSFDaUlb^N2VdR2m0XL6P8j]@h4Rj0gp62nfaHATY8WRgZLMk07c64LX7gI4dQZ
lYj8b6SK^mCcAi32;LRS0Y;7m]R9;AWF46V<Y652]@Oc>UXS2hiCq_FkMIbg$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR2T(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
dFBZ>SQH5DT^<gWlg>cSGY;GRKh]IQiahPaY1[<PX\i??LR6pACFkWMnF5[?4JB4
`B5KLjQpcMA@\Z;hU8eAjcJbg@E\BEK1[SYD_Ag6CYB]\R0nYPPi_T\17_FmRUI[
e8H64QU@Z6JM8YTop3Xd\S4p0Y73[9?KnImY1mLK<o>;F8VY^Lfcd:HCpH;Y`1h=
pamW^FLqEZS]?XA^Pei@bQ4n[cgJ^2:dk`ncXDi8\XOY<2iAME5L]6_D1[[8DDV8
p<fR239A@dK>]<7iGW`9=5n^9MC3nX5Ob^H7AHWW?PMAIaGgbHHE;ik^8VgS7LE=
0<B87a=hf?3<o[IeH5lfpJIIiKgl8I5\nW8oWiYXWfMWUNgdZ\037BbC:2S2l4o1
@AL7DJIN=92GQP^8WTTYnJFbThL6M<BXL\f\OaR:qZ@NFOOT$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
kOI<>SQH5DT^<^T:A;aeA`I0M`bFcbboZa<2=Q@CDec4M<g8bo@KZjo4GBab9oq:
0KVJAD5kFe`=Y=>k^IQkoB<d1DbPn^1[OJ98Y6qX79_c;AYOo>fGYK`N:^IkBHiM
mGQRXjLO5`ef1qUaE@h`q6lMiWnNYQLcXeH[K1liR\@gZ5Kohm]cj5Bh]i7Mq1gB
PmU9q2c\XU7p:^Zo9D6ihjkVFYm2j=SHRiDcBj<URh\F20l6lXiYh>>@:Pe^Qhh5
Q;j_X_jYUnk>\SEDJYgfY3P\X;@6^U@a8_opUT?F=GcQFI3D]Y@]L^S]5O;[[n=I
RTCF4cT8nADJ6EOkdanUmKRUI5K]aJ^T1>4FU^=a5O2=V3`@e38Y7h=qCUEjLKYK
DVe]1TDPW<5^O]ko]hfc2iMUO083gZAV^lM[iS7gj6NKVO0R>jN_cYoBCACg?RjF
@089CglP`44q\;dBb3E$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3B1(O, I1, I2, B1);
   output O;
   input I1, I2, B1;

//Function Block
`protected
Ic1SdSQH5DT^<b[Ra]gbTRPIBF36EXTSKL_43n3`:J:gIaZIURRb90QIl2DWP2H1
49hjiD0E_;7lpVaCcSeeEUoUgf44GQXkmROKhiiCNf]WU5XCgBPK]AZ6o<3`Q97\
iJn>5Q=E;F[1Idd>A=B[fq6C<L5F3N8aBZiGeYElpZG0P9mp;U<8>80b3N<M\W0o
_fD]Jf9nnR;H_]IX4lLX6CYqRWRDREEAJR0nS@mlUgo<L2XSci\pkME0E^7pm=\V
Ikkk9\99RPQ_L?Up0Pk26^pNh4MQRYK16D;jOGVBiRGN;K]16[A?6[Oho<_g5NTn
Eb5dMDZ0\>[ehTQWcg0<RJe@0fC?LVBZ4N=1m<:F@Mb1PUqNUa[?g5_;Q4_AfEgd
2BS7KCDG<KU6TfVX6@VH;d_l^QXPh>B4Sn;jb\MecR1Q?F?NoQZ9J`^XT0\2T9iX
?0pQPn]7A\NUGJlFg>`C3gOT\b7Z;HlkcSMoJjH8mDTnHb?AofGSIZLagEcUg3:X
d1A`7N9PG<<<M1gW8HY32WfHd?pL41@RKl$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3B1P(O, I1, I2, B1);
   output O;
   input I1, I2, B1;

//Function Block
`protected
=[SJ]SQ:5DT^<9ga;:Gb17dIB5D2[=pa1KKMS0_C8S:TW2CD^Q5aD[TWlo6J4NBh
k<>PiiA4cJ_9LHLE4HPbNUp21lDW@_oILRI4?WKOO6^^3qSK9ZAPqcJ5kn99\J>a
ljkTjE\<MD_I=?8Qd1T?oJS@]d8@q=@:5^E4kUMllnQcUW^lXWhcJi03p=e^i:KT
5NCRn7W88oe2mSn_Y4Io\`e3PelAcmlHkXIjAZZ4LC38>VRL5PfMeq=L5@CAgpg9
dDkSp=KW;^;[C3hOBlRCJ5D3I79?oR@ZIKOfT1=WfFHe3iZKGAYWKGE_D^9=DcJn
PcX5[fK^WimJfN6X[3m0h:OVE?Y1q^F8O\X5VIZmHCIeYInC60N>DEV8fO4871V]
6oK8_\MjXdP?987RFl8N_<YfYX2X_ehmkoX[e5Y[HA04PT^NH?nSq;;R>Ck4XG_l
S2WXSOiFhZFaV=4d156`<Z\J;FX3e3fGKL=oi5l6^8AmL2[He[;:@T_<EXl]ooo1
AA=ORSROSe>VY8N>qGJUaMKS$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3B1S(O, I1, I2, B1);
   output O;
   input I1, I2, B1;

//Function Block
`protected
_8E]WSQH5DT^<SMH[gfjdb<[0[E>3E>HNQJDIdP50N^p>_G9]HkdkTEQe\lZ]VPb
pYJ\Pn`PZ>7f9Y@cEA2l=4:QBQMaCZYWm=7YId3QaW[gRWNNCV5[LEf:]RTKi8C@
d04pUE6k?6qmeE@`a8ZCfZ03>P@21HMKMG^^MeMb?Sb2<0a6AmpIbX:>WeVOABDZ
AQERTEJ;_mJB]7p0JU?lFb:_55:Wj`2f1jK;ciTDK4T7hbF[XabY=LbLUWT8LA6_
o>qDlFf\]<q86DVLWpOQe5YoU34\;A5b^eYN]L0VCo1j_VTN9_8DMkHRmbC^15mF
2<e<l1]_ibF;1HkYZ7TXf`3^=[4TN<Y<:P]6Te9?PpAL]DK>29_o^P9b8?T`K?G:
SApZMD@Ue_hf^WSAJb]\eo_<T]QfE7aH^]_UfI6M778@Fh1M2LT>6D`^l;[3h1G9
CFRZ9D=DDSf60@i[XZ0dNZq[47:Me>M1RBOCgbam><C9GY`hf646Z3>2oLkPje;V
4IhYjJ;Mf1gf_CQL6FFj\;S[?eUNOO6FKX8TigZgY0p^onLKbD$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3B1T(O, I1, I2, B1);
   output O;
   input I1, I2, B1;

//Function Block
`protected
gE`C=SQH5DT^<TFHX`C<23^m;7ii<2GL]caOOmGM786VcQXGWe<f46VIpE_o[XG9
l^Aef>iQUR9`mZ0I0e<J6TkK?ZDDQW;En=oTD\1dMa=;\qaBB_]DnbU^KC_F:@Jf
GK[`T<V`l<cTj>9`__>=Al<W6>11qO;6HO6qK_hAI18P3IcZlKQS98P=aU3a^GH2
DS0G<lDPUSHq[1E;[_c9_N?8J1\iQ2^8ef=LnSjpPLV^`n8qS?JEL^q\Tbhc=i`c
PI6ckaH;JM7JndeOm6XNHkAK9:0Y@>82OiG>H^2aPjRT]B8Rb6@d[7eXHRVl4adR
OC2=mKBJ4O>Z4kq`nF\mE]@^U\]9BkLEb>8\0=\0EOnYILL\@:cJ>WgAY@\\lVV4
ocfFCMOnF]f<PZl0=>5_G3o_TPPS]ZlQbKgYB_q;PU_e:h_Z4ZSWB4^2A=h7Y\nq
XPRXIB]TBIh7HSZoaJ]Z<B<:>F2MFUa`<cnoJMN7oON^^gV83gFJUFE1j=M[?h0]
noG__W>VidDg@Qj98eN]YXh1_89q:g<j_EP$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3B2(O, I1, B1, B2);
   output O;
   input I1, B1, B2;

//Function Block
`protected
E;l4gSQH5DT^<JaH9mbR]Yd98A:J2=lHgIbUThkS68PP8:S_46AkEVCHQ<;Wdf63
WfNE;Z8qj?aXhgn\Fhle_<Vce2q[EjJb^j@<7YgTjT24Ia60G;Y5\@d?7DHloR<q
faB6QOpD:ocEM2Zabj>\clGU][k`=mXP<YTVQ6JIh7lc:CqPSn^W^\YHc??KhIIL
KbfO_\]UoOp3J3G5[eLV;^2K\gd;g1D>QN\qM>O^2Y1paLkUY?pJA_]6GIYVYJiJ
bfbhlJfWAf[@?4@R3En;imCJ8L?JS>YLe]RX<^U6Y`YfRDI^el<JC0;[hBmBhHfY
_[YFk9qk@Y5GNI_iQ0<C4kc5kq_[\bkl<:cAde0QiM`GB`Y<<`2V=HcVBoCa^`Y^
:E]PH2@<BM7jTEMl?iXlBIbd?P_fSii^UNC4fh57AhZ?Hq>gR8Kifc\MHB1CVB]:
l9Z;8bH:c]J]m5NfncDbU><e7kleSMNTeUKO\?1Z^jc:6P>cd8bHh\AM::WcSkWT
KqCAUYT>b$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3B2P(O, I1, B1, B2);
   output O;
   input I1, B1, B2;

//Function Block
`protected
52QNQSQV5DT^<`mHL^OdY`SDp\O?fn`fbTX[^Gl<[G@h<Z4<5O\lc<51Y3=Da`=e
nC6L8hmES]3b^`9VXd8_<Sng4iAqLI4<=WEJoZQ?aZb^DLSXVGmGn\ObgAFCnOYP
DFnA=_Rc\4HLYNBJBdXH:CR5l0PmiZq>bnb::pnoCD=KTB;Pmbkc;fhfWSB@P3:m
i88QGJU\J9SUKqLe^eSXA=HYfcR;71Y1_>L3lG@kWpOf[F_N0oJZ7UgaI8hWZ33T
RTq^iHdi\IpWEa3XlpQ2S=K_NJJ?RI;@j^5meA9G6Y?>Gd]LNYbeCQ2C7]e<SkDF
Q\dLmSnk<HLgnhGi6=:Zj4[^=MNgF_7X4hX\]FNUapATej3?h6P3=:?\\anQb?0j
I=?a:]LmIIf3SNn:C`8JX^aW5UM_:][jFC@\?K8eQ=AVom^D7ZG408on;n>Q41KF
`_AoaqNWXZ?:oKckcSBcKTeLJI9^8=S[VKOCICoGaejcNHMC_FnY<H]NkL>c<jEk
aX`^^`U`TWRPINgdPdV5QHcL8_fbdX2kcq=^?1[ee]32ifFiV94hFij2\hOon3S2
:aOaQ2n52WL_:OLUY:Z4LGWoeAEeQCiYE?qJE0`W2?$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3B2S(O, I1, B1, B2);
   output O;
   input I1, B1, B2;

//Function Block
`protected
3IhHYSQ:5DT^<`2aahYZ>ia=[ok[8VjL3F;1GPqBXLQo=m;MZ2jNap[f:lBQTY7?
:3EW2N2MVX9H6Db?`ckR:Fn?Pi>oZ=fiTfF]8e;k_ToEWN]31QR78h9PQYBCMq^<
L4B1qhSkA37GB^4ijTGaA;U:Pa]J5F0EZj6gXYFbBeWgpJTA2Fla438im7kEcD5@
CnB\SVeGp>NOm0QPXmD^2AaDDADKl7m8Ypg:e^8kap`Sbb;lRKAElTRh1kgB6Eb6
6GhIOHjc:8mX8HhHf]q^;ogGCqLh6R31M_mCF60407BmY61A^03_gQ<3a>Z[K_NN
;L<HC4BKGZn=hWY]<hYl5elRc:LOf@40;RG\k=VaR>4A[qno]a7>U5B1jO<TddB\
<i]ed:^_eJ0QZfa7NoC65C\k9V;7<;Q[\4234Y\eS1jNFNn[UE?]WQSfF:mfOXg4
Hp?2=icHhhM^CNC6a:JDV39Tk\GUg]mC92emXlNgRmUheL0N:f^XHbG[AA>^ph>I
<FLiidcn1hknRZ4PH?[\;FOW8X@mmTBb62j8dSGB?PJOc_bWABH@Fb5=D2`81hQL
mWI5>0nTNG63dYN_p=2Q^eYB$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3B2T(O, I1, B1, B2);
   output O;
   input I1, B1, B2;

//Function Block
`protected
?DiXJSQ:5DT^<k3`OXMC_41gSIbYoe<eK08ZL<IaemBo>YV;i46q7Hl<a562mg@W
gUKO2B[oia=Ll<NfZo;JViK9TAWV>jV^XgUa0Q?BkApCZa:PQkkfNKXB2HTmW^aX
9eTL2cMGi;jL4LhjDjYC:F@h1G3ZeCEq:`EUB`pO5Q<h^hP`QX[3jnV8OadVWX3g
8:GeQd?90e5]I4qiIBn=:nR\gHf<fC`kiUm7im6cHLp1aRQ\7cQl>7]E:Jo0]A5g
oH]pl9S]ciSq9?:045D2h@d9WM=SA?QT?;]aVL8Bo<dk6Oe64FE`B1XkUmh`4g1q
d2IZ4?qMf\=iM\DAPDBS3=7Z7YEm?l8d6JnC5hWOWbV_dg[FEI>MMQiDiXBUOg=n
kj9\49:>hLlS[B7dM_=`gCW74>O52>qa;T7:M54TSbEXdGVlXj]<CR5QPjEgRT9j
XnNAI6Ah_hoH@@gS<\EP\ih;P=ao\WkD7cMZUeU1X>1;\n24Xc1M09?H[4q]FiR]
6JXW2R_Bg56BZjE;JR5aYBV62d>Vj>W^286[AC_^jfCNHK`WFmA`?:h_el^>BniW
iD3?Ph<CjZ43ZYW]91maR<qB;o`I?c$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3P(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
M>EL]SQH5DT^<4MHEV\iF`RoKa>Q5Dd8f9;7@ioKT^j>O>C3_aYFIfn9RbMB7h:G
pMLPG>hKHBeIcS\SAYRKFgHF>FQpaok<f`_KGJ^I@U6PcIqYX:E`?q6eV2`oIZAT
A1^CfK:LGXM^9eUU:^hS8?gkBF]5ipo<n9A2SpPH1O?>p`];ik<YRK2ifZciiI@J
a8oMiXB>^DlKMZV7b;7eZfOiK;X2cCG95lX^jKYkCa6nC>omQla8aN`M[jPZTNg`
IMNlqAK`1U=J80C6AUX\8]E@4V9gScAbl>oOiRRkdj>AeHP:`j=KjMSEd;YI4@Fn
0<<1<Z4T_JoFn>>\2358eVSgjOG0qMS>=_;f7\C]mO?<REIFhII3DICV9O6F:cC^
B6nQ1C`g90;@Da9LFIH8iUQlAgHI09=ShG=_MO:P\LJC`I5gf]VApYLb5UDX$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3S(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
MU[b?SQV5DT^<QRX0MS[\jGme?SPSSHmg9I?1TBn90[4G9hRTc^6iW7]X0f=H7YU
9o4m]MFAB;\kGZXq1AGFbPUGI>Mo2<j8SlCai324Q:1?983Zi6K`cn[Anh;;AU0]
3gR[^Gi99:TafIdqX?=BJ6Km@dK;OjP79bel>`mW]54gQUMe@64=oB;g[8MnFS\?
9a8h0_?Ak1Tgk@3qW;UYIOpZb_Q3R[n7C74\TF>GM[GZi9J>GZ2F9`Z9\LY68XpF
b=N1g?pY^44A<qb40dX8?JK]9@;ZpQBIGnomlU1?P0P4FHj?eoH:dH2ICJ6?ciD2
FBjn>FR;h[77Uc<0D=H>j?:l>@iB>Q2ohQ86]LGS\JS6maY=p1C>chi]9>kYU0Tn
7Nf\l7noeP75YCI8lKbS>H<K?1bRRFGT>jlo;O0DIifQ?binT1EEcmDRm3FRm552
VC9HpZ0mFEoPBc59X\8h\i[_SA=;Xi7M0eHD2?iO`=06Mc3fiBY`8`75Pc2SlC`H
bhe0=Zg5KRY[Q`6@>j^e]0a9p6eYAa7Z$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module OR3T(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
e\ZEfSQV5DT^<hgY4]N0U5Ch>UlQR5=9pcHOKF7LHD<OUa`o:qn60k`m<0nWnfEL
=9QN_LERFLh=YDHbog5^D^:EF9`dUJ=cG<qgGa2eDqNV7LlC5Y;:8D1FAajjZi_S
b;KN7o;^]>O2Wj4o\p?jPD2O?qQPnL?6pDmO?UiN2<0JOO120XJLfP27RH^\<TQ2
^Ed4Ec5ga?DJ1[P2K5g5bUdbnc>kAT;\n6h><`>OeS^??Xi=R^oeK\EgqGA?>aiO
6fa7ooVk62?^\0VkY<Roj1Jc7Hf=1F7ToeCAIHDY^WkiG@IS05`oUdlC6>=5m1a`
lSX0en3PcD9g1KmZp`Pf8QoTZIJeag7k98LaNAV\W2C3Fbc:8X78;XIh;L2BVfEj
?A8inhUgA>d[ioOSc?8P>md[Lk4ToT9\USCH4@OVpS4GASN:$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module PDI(O, EB);
   input EB;
   output O;
   supply0 vss;

//Function Block
`protected
KdioFSQd5DT^<[@i;=>LS7bHiLhVoGVTQ6;3@C\^TS[jLIpXG0ZDJX?DmkV]maNI
XkCZb4VqcBWMoYHQe4fYi[jP8W`K3Hl9e\KdJn]RGVnAhO5:9kof@HMWnC]g:koE
`4MkhMfDD4qk^XXD=qLeUn>CY2?W1WXabo;ASY8a5j4b<_l[h?GBq@VJT3?6pn55
;::pJ[kIL5iIYN4;bT_U_]QWIfC\>K5]4E10L5RRln<XkR5qejEY>PZI_T]6d>eJ
LJV;To:OH\WTSCY24L5VTofT5V3lBSH[<4]e_?JbR]TAo8[JUCmZeZR25kcM>3Gc
`<deQ`\Zm6dD2Y0CLmdl7O^?0fDfdXmTUgKKY8De<3eh`XcQTMLA8G\j=>iii3EB
SODCJB:f5UWT5C;bDM5D1UKd8?T9BMX\m_UD:CWZJV>EP<;YY<R1EdWEpm0KLO]b
$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.3 --//
`resetall
`timescale 10ps/1ps
`celldefine
module PDIX(O, EB);
   input EB;
   output O;
   supply0 vss;

//Function Block
`protected
Z[]dYSQ:5DT^<OW:i>9Y1iZ3LfkFhiYhg?^>7`Li9l=mRBL7;BfeCZJ9N^=p5]fN
H_;88ZCKAI:mOEf:FTncF6nIT95<a8GPf4_E_Z?E];bGQ0A5eTg9_cK_<3mV]ZD9
OdqmhoJM4FBohgWgLDXeJfS`LTGe:Gg8e80qFP_>[Gpf7ka4;m5cXiPdg5U`B@Gb
]`Eah>9_LSLnA4?]O4hFGbq2T;7X?<q2m3NH4p?VO@_nZfP^Q>\mfIfR2JBBk7gT
VKLHUJR^0a01d`<YPGF2KagGRkN1;0ibSghfEK?kol6fc@=:mB`OfB6E8Td:cEE9
b0W=g^X><C7LS1XiFf?4jflQ4_AfggB2f2R593;710f8H@[:mB`F@B6EOTLodek]
Q2JkGBWL>lA5>X<9g4?4F@;G4EAf1lB2S[7b9AkKO;hHf6ml2I_[WPWQW4qNPL]h
O1$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module PUI(O, E);
   input E;
   output O;
   supply1 vcc;

//Function Block
`protected
0;3QlSQV5DT^<=ohS:^?6n8IWoTDnQGJN@i3jaGA@mJBAEW8TOa6MaAghiFGD[==
bJhaJe`PogqMSfjG<Q?;0FXQMNaD__AQhHPf9n\_XOm^1F:Y27@ia`0W]0ng<hZp
F26k9b9SBZ=e2Vl8=T@QqoiC;FLpI13TZ3EZ23O8NgKoFTdkdPPI\9M@RO3^q>12
aX[jp?Z\EGXpkW:?]f=U\07BQ[EKQKXT>YAjI[cVf6NnDL543=]i\]7e3e?HjXY4
C5KcI;5]ABOOfNY\AVS_PMc5^GgiRJW_^4lnW8?XN>K<A9>BEI;:e?GfULE\8jG>
3oVUNn`UlI8RIZdmXfoRn\_G`[EhFej\QYAPQ^cbS6]iCGURF;ea@EK32h`_:1Fd
:bj<8F:eimH\2=PjaM_qQli32K7aeJdY_Blk:DpUooQ_:o$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDBHN(Q, D, CKB);
   reg flag; // Notifier flag
   output Q;
   input D, CKB;
   supply1 vcc;

   wire d_CKB, d_D;

//Function Block
`protected
6F<ObSQ:5DT^<5T:=W3bglT:V4<pcmW:M\]T0FNZh;f8nM^igI3SnN?B5oO\QI5g
Un^`KoD2aa?PkRZi5W1@bi`KDf\;VAphJ\fg2;lDY>`29glM_2m@m__N`X`K25mc
Yp;F;;Enp`bI]]Z>\1RNPm_cj6\TbaLO5]mq9NOJhP@0iiL1ATP4WD5;C6elAXP7
3h_VSi<<d?UUCEG08nO=R5RnnGT59dnU3dSPe1qLh_\>@m6j^M[N8kQ0R0QUdTSL
e<NUQU^qPL3cCZ6qim[a>i3fG;koohNI\56bS2oPXnb4pRm7aAop0UgEGCWI:fKh
<NO8aRh3ZJUDBlODiU^LXm=KQ:TF@=15SUU?2fLL9ohH=:BFfKk>X1Yo7BX>LShT
7bhVe2U_58J:CG<l67mOA?8HdE>j1^7d69p>;Q[c:5BC49i5lF@73SCgD@=MChhA
lh22Zm1JPkS7]KkRaP:PJdIgZ=K3Wg4CM?8>g=>T\[LX?N8QWOhRKpcW3[6hp]Pf
Pb1W=9R_o39XbZVf^BLjH=<MU?CR@MX:@]=0pbZL8PY2HFRgb=`Z9K06G];_WD;;
2AJP[_\UEN=`9VU=g5JUJ74I7k@nNn7aF]ZJ]MSp[:1Hae7HJO1;@2HdJ1Yl=lM8
5e434\7VH6CKQjq>K[V_MmHL=T]7c^8?_Nl`@Ml09PHmJgQFEjETTKOHF3<a;FBb
?J=UJ8dJ]E1d9oR>m;k\X0FB4eXMoZ0<TE?WHkl_1QWII:4EjW7^7Wo^\7LQ07AX
7:;CBdl=]d=dWFchG5qVnkBX`;PaU3a1C5adm0H8JkObYihji[V9eaD_IQb1cMaI
kEXXj^J8;@;eMmPVKCEVbH==XX>2OmZJTkM98ESZ[E_Cm\>Z<ja[?<KZ<Wh5=h1o
?PHjEM@N7K206id`aJKZenqZkjOD2qC<S;Z:^jSS5E\:LQ]]Z=>XEDXC`bYlFDB]
Q5eV@q394Z@<==VDO5m[;GU`k<P:Y5NYfBd1R[YR_>VFU3Jb^fY_Y1I343D2nWa`
ba1fj`mmd8WP3ik;6q1=8RYH\$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDBHS(Q, D, CKB);
   reg flag; // Notifier flag
   output Q;
   input D, CKB;
   supply1 vcc;

   wire d_CKB, d_D;

//Function Block
`protected
J8ATmSQH5DT^<R3bD?=i>R]=fK\Z3fb8mOHnf65OpA:@cN]fCffM9mC0`B15WbM5
J2UafeP8:h;F[UibdKBODRYq1@C5;oWhPj]Ik<\9MRYHZg819P[8HFY?5amX`7ap
84QhO6qn9O8^7lOlG@:0lDbo3mQ96;447qCe5d4a:09=D\cS;aELQSFNnCK=>bWJ
4e81<XSO9Tb2EbBSTl5oU83MfSNE40C=[9Rbqc<:X9=RdCXS:<Aii^IK<Q0;^9MO
AO<J@q5OC1D[fpWk0SY=pDNRh<Hk`nE\_2eD]82^;RG[AEnccc`BScGbGfn=D7g6
V0ROUFMGlK7UiIOijPQha3G\mLQ9PkYk=P=2Fngae75BSMN9e_a32>UBB?CROmXW
g5JqO8^NcjMVXm6HC@b5V=QEkm4bdF3^@[1kW4IX`hZ^UkX8W<4gP2DmkR9lL]OY
3n[gWjMLJlLEFSUiB_S;CZP3IWpM`KCiIO4[lPcHN?GT;e:W[^Aifh^N?m\HYU<q
S8^5ohqNSXjd`f>7Z=@=[>?OIMdS8TP\jQ?lR9_Uml780iqVIC?G_4@EWWTk[KEa
Q4P0UXTQG4gk8U`9m`\q2iP\[J>NBU0<`HWo3><22=C8`l9VWmckm[_6AJAgZ4`Q
XPPDR@7]Qj<o0<LF??kB2I?nZe<k^DLd=:o[h8I>LB45kDIY@44f=3SnD4O`_^2^
FGUbgSMn[TQZhWDOkKiLnPhpOR5JOK0fQo>jh3jOHP8JZ\^26PRF1mFV=YLo@3Da
TaohNUUe9ajnaegLGf2F:K`:OUgfJSUYkZ?AWIhWjM4XTLnb=cnV10J;92_jd0V9
Y[N:E_OoH=^5R^>YQF?ePIJZ2UOqcU[1hMqTR`?NJ5HEI1J6;6b27RYW8=P@6pdb
gg1H0ITL9:W^\:fL0NT;IKW^l9<_Wm2iC>YPNp2jRhC2gDD6AKY`e]XadKK6RaQH
gDUoCFa:ALOK1[kQJYP]^5V\cjIX8:kWO<gAhfNDl9;DAmjMSqAC6U[A3$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFFN(Q, D, CK);
   reg flag; // Notifier flag
   output Q;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
jeSUhSQH5DT^<?2iR[8]Jo?`a[O0>cWbo=JlEMUOHa`XJK8bo;oBe6pZmT]hB;>i
Y<D;h8A[K]PE8=^T3;D_[6`lM[LY=jIpJ\?S^S1k;_:N<NbP0\4T7ZiBeB4?FgJ3
4@I3;3:a\K;CC[ElXEKHmEm9mb`AgITML<8KfZiCpd\@:J:qC:O<k=XD[NU]afR7
YQ00[6CbX0pdBh[i>M[MJ1>ZPdOmQ^@1JE\mjX[S:T3oCiK[Rm>d[RoB_b;k1SK6
OM@]Y<0[72?]O6\Ojn11eM:flpQ>PR9iGpi^L^eBpFPo0YV;_lGhY21h`dRe9eSk
:P?`76XFJSP2b>;j^;SFIA8P6hQq?Q71`=K5kL?i;8Q4XZoV1=mlX`QcX3W7X=Ad
djfKMe?C0BkO1>QK;fLl<9WM_k>3o7US6>S?WfKLii>Holm6P9XK=ZOTcm9jY5H7
=PkAT7n8pgA^6^Ip==^04fGQXJh5XGnZPHGENSWLSf7_ORIc6n<bY9p4M?G>]>S1
jN0lS3jgfl?0V3Q;=XmGX4;`=GqHo01Q0O<M_SESF_eP7bi]EA>J5QA`G5]Q7Kb=
_Qn[[Ma1KZB;ihJUI5SeOYE:H\Je8LcV@dcjAIZ5dAcjUa:3fAbO@<j;>mXbUFNJ
?l8\30AFm\_DV0SR<glfH;N0o6dqAQCMk3HoCn]mRmHR@:Bb]]@aTRnJFT7@`EI`
HhJH7IdZB<QDnB<j?=e[dl9KMi]BUT;:eAj]S77P5@87VUSYBW3DA>nXm`b36BaA
6CGRN^d5LX4Cdin5Dk<meL>a=HDAqI:SKSQhTlQ6eU8`B99dg=UQfngmi>R632DH
DY>[kcFDocgTZ=[SkSi4[qb11EYnq6G[@\T^hbfWjD=51KJWgaaK7\ooc6PL9^o<
QIKqk[1l@cJEjNmIW`bboD[DoE>UIRA>9=9Wfg1D>^p?=GQeN?Gno@iEGeaj9Y^[
ifPZLjGJeUOJkOhkgEZBeI[2eQKGngD16=QdOFdEKH[EDBj`=H5CLpDgd5c2UTW@
\Coc\W0DlAmdfc:4]`45`>I1mQ[fDc;AehO?Nh87AZ4Ji9MflQk?[nAiHmIbd<OB
pnQ7S3\5$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFFP(Q, D, CK);
   reg flag; // Notifier flag
   output Q;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
2A3D[SQH5DT^<HOXjWIJ?[<cl6;m6O8oIog4U]C?9aDG?n:UBVZ[23=2DmO`JKWG
kPGpYc1CJ;\5fP@a3ecb3jCn;cNMa\ml85qfXB`ci_o89dNU_WM5Y469`9co>XPM
ETVfl93?43062QeJV1h1GbICMo[pdhbZbDpEF5W_NO>e_a^EUYZ?Wd81U1S91qL3
_=\Z<LL@>LWEUYfi;lf5QS_k[1ZASONa?bVmci87O<?DNnS?0U[lVjdLF^]kHIM\
L9^SNBTDQHM^qlYKQ^_;pMM<]OdpoKE487n[G1;<ThQWM5o\gJXn^KnCRae:88o7
>k<8jK2@0ZcPNI]IY8oYEXBoBRlN5ZVSkbm;;50<:kiO=N1KUCfo`28PBoNjW:Z`
K[Zm>3KZqDB396kqXT[V=Y?3K?bR;Ra\1e@n8OW7@V4Ob4:KRKYG8?qf2<>?[ZnG
XiPJ245=KVFkl<O8cG>O0R]>lL8mN_JP[N\PD7Z5V^j]a^?qd:ck;WPCkobDNQ65
Lkl<2EC7=HgG2KilYE=pIo2S]OI9GFOKLI:T@oJBI`N?iUXNZH1iMe;I:Y1;MVX]
0X6XfSFga8ZV0`Md?Olj\c\nB:YcBd?PPfM6So5lo8D:m01H@\J6a8iTGhBCMnNg
8E^25YMf@k:0L9F1n@KmplZQ7ikY<8heb3H<\W<cl`=J?k5af2FTBmlWoI>=0m[o
J;eUm^LiV7k]R7gK<I>Y7g^0h^HcHQGA<<@N^;Ia<2]MhiNT02F1XhG2odL>T9JT
kZd?`Ln7eGb]7]C9QpOFmB6iRKL<nZBZj[cMB?_e7^<f8o?]oZJJjWFN:8e9X[^n
cC_imLZbqjZEneDq129b15>=Kl8lmU1A_>NCRFIQ3lK0GYm;VN\D0opIKCYBfPB;
70[:UY6;J<^Rk0EWD2OO21RfnL20^p3Q\`H[i6@Im3NY_D1BddUB^L1ZT\kPVMEQ
fPSUeaX`W[43L]9lBd^MDfec?\ZBD0Ig:K]Tq]<_81Zi64l@]`l>1=JfXlY;m[5C
1>fSd1o^dcC5@Lc\lT[gjH3DYf?hZSoK[Q:Tb[m[dmM;@^SpHG5iTi[$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFFRBN(Q, D, CK, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, RB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
?VbSLSQd5DT^<h=`7m`\inq_R^]iJ<k0_=3?UTTFM[Q<G79CCFjG0FnB@RY;_Ff`
6]Ii]ibmZO`Yj8e1E`V=?@fiA\mD2p5FYX:_M6S0:jm5SAK2nLjKf1>g7^d4k1o_
oLhYCcK5H7eUeGBJSbNk?>;8pP<PPb?pJelk5c]lD^MdCA=070UlAfbQW?qE^dWk
QWc]Q<fD[D6V]An_2?_Al0QR\D7J4=NmaAmbRJoUXWFYAIT^<E<n^^>oDmh0ZDSE
RKEoocT`KbpL_;j\\Iq3NF8XlpHP^:EQZcl]YNNoR31S_l89]9j[6H?`72Z5j@VU
oWTPeVkXJVmU]3SaiBDD<;_m@YZ2RQ[SbC4S??LDh]8^ck49l4:[i4>LTSLIXaGi
PV[[]apZm9l1dZFN3:S8;GmTnb5kPV\W6WQ5?:AH02F637jKmbFO[6YVA9_EPLK1
[8_Qa2DZ]9@1T3??@aV6hR@B\M8T1@f5UZ`a5V<U93Kp8GO;mlpanF?;=DdncU=6
I?:^?7ATm;QV4CGGY1;a4Meq6`mObCmI??Wf0B4Q;l]]\N974d_eMAhaXgn8^h;c
ES1e_:bmQiD=L@d0EENTpX3IYSUT9nCmZ[hCBkSGehLYk4g=AC`keUEVqMBN7kOf
6GAZh1LGjj59DH>S>X6G_H?YUEGAeK3emRa12gB?0k1ODL8Zj[I^1mCDmH^A0W?7
BYmJ::dkkMXaFTEn1D^<CZlJRR<826iXH>8M\94mi[biUdmYF=@[kGDmn6mPD92a
0qX2IGejGoT7gi<9g]Oh@:3ILBC7LY:\M\goD`T2L5@:e5VQHa@T10EPIm17GJ?0
V]jN8=lU1538DQEHM35[MeM1SXI7Q462?T1_@Imo^m:k]l]QFdBUJ<mO`5h3H5K_
TYGcNiM9eLqPd\BS4q5f>R[WkgBAG@nPmD4`9<5N2@0R7`Z4m06?]R6QgU2Sq\jJ
6D<WNYDXNFSmc1ZV@ghEA]2HYcNZ:?5LcIZhiOlqD_IThNC]^bPm[oUZc6X;dQ?8
QX9VLREo`@PflI`R;hh3b7oV<Kdg7]ZP@[CW;cIWL5CH03HSGD:1hhnf5WnX;>BV
3ZD^T4jZSNH^8eLWfmNi_Y0h42c:0dRYUKf;e4HbP\Hq^ZXVH`q`olFIkZNdBUSD
J:LE;?b858?>;44FH9_bnJT9QaI4@4q@MJLZ:kNImA\hAAg;f:\EC@e1S`kbV<=9
cKDq<U0UDelV`VoDaWhE0lZ2_5IZ??:8_>5VTI>UJPpm4RXFNe`cI5IfohhL:;@F
W`8WDS7I`la?H3Gpc30o0Z[mjb@U>n=GkUM9>SL?1OiJ>IFiIH3?ZUaelW:?hTko
njYOM=S?oje?CRbaNK=Ii7[@Thq9NhgNG5C^j3ibkB7<ie0mMHMaU4od;=ol4f;U
=AZ9@mpJDAWWcmFi4^CiXFHPL<eb1^ZVWcGL;F@lYJDo=9[mSHMOT4YbI>M2_h2\
Qa08W?UImW1m14EhDp:f@dEIJ;iHACF3oTOS4H1OOBlC=_X8i4@1AbUaSK4LiZlB
@:RQi0B80mgC:4NVR0\`KZRVqnBoG32c$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFFRBP(Q, D, CK, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, RB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
o^3STSQ:5DT^<nA`M>`DB9D^b?gHAh0^M74qGXWJGT10LG7Y>nqC1hJb@9fj4b7m
RTVl:TLRSWHN?P44`jf44C@kDTomVp\4cleMqO^L0V0g8Yc66@ifBdMb^g<DjJ3p
S_iRI]`<dlQ1A>WlEn3LZ?93gJ>66YU4<fb6R@kLeohZC1U]ofn:gn_G<ARF\OKU
D@hie]@G3>Ga:f9q3mVZ]^cq71;8CHq5oBfCcdL0Jn@hhKV6mIdSj4XmbCOY3c`G
Y;[nBGb^;6hFfhX5nKhGgmQaTq4QV;beBjYlB:;X2ccX9D>AAag7JlCQ<>^\okR5
Yn6?AGR0;g?@8U]QNAO29LDIP4efH:g^R6A0\3fDXFBP2?fdIZkk3MDdL@EcVOlC
F^bgaUpDeeabL`hWm;]]ii^Q220lW99D@naNo@ahPf@RCU;FNFkV1G@Y3>ZG47A<
Dl:O`>;Dkeab13ZS08hlDXjI7if<\I8Ok>0;T4oN^W:p7NDSl5pEJVlFN8HA?^Nb
JI<W7DH^C<BU\;_MCkmZHHc>U6IClee<VFH2EdV2af=R_Alp>An6][jK39E4><67
455idQHK5b<TGBW_1fW0pEbg6[e`K=3\PUkn8V8TIR64?>QV_`@keBZoq>2KA4gi
8OP>o<lJ[3E]1kcm6dH?GLhjj_cYU^Ram6FnIQ`@[OmKZKAAf[m4\lSF_nAk^b7h
o58V8DRa2G5<>JVN`DTn[^6ZhdlXnP1HW<B5Fg_QHc[P1Z:TlO_hRUKnd3g`A49e
Rq_aC6dnT7NSGjkClRj2;UlLD8=9`o`XlBdSV9U4Y=h;:d[`R3L9D4RGX_N4X:bP
13KD@XO2OU8Oi>XcR^Q4NB=B`EXFbYW`:^0jH<[eJfZ>Bm92hSUTMc\SDV6iI1UQ
6M@FnamEgWqUOY?Z^pDeOahA?TAP9^eea6RNeV[0HiV_G[LiY`:5Z\TYbRFjp4PB
mJ`WD6KP\ggMmH0EGc4I[1<6mij9dF^@aCM3VIGqTXddF1Ak8Ne8QiKl=\hL@b[f
]8;UQmOp5M0WD<el@0OlCgC_=6Cc\Y]ka;?k?ejdQdK6NlmSK\iV0XgCfXZl;AoE
:F<@2KVQj2l4oa8Vo6Nd9LaG7:><_Ld[:;[J[WIfPQ1^kL6LaHbjjZcK^?E7?DV:
[m[[7O12XVVpm8OoBSqA7`2Bf`:VI^L<E>9]f43NLHWWVjV1S`H9o:Bq2XiXU8`m
l]b1^kBha;IT^>HD=]U@8foC@2]kQ^p[ZhidOQOIN2cdNjc[?KG?mpU>CX^=XKAF
S@lVoFX1I[@VV_3T6_fLK2UmbjqS@1h4Rki_cL6mD1ZL[M5SPWa<BI0E<\6oQ32:
Sn7gWaWkmNV9aXO`^O3?A?ekBTThGgf4i8=0MqGkXCYNTa6@_G51^:ehX2M^5CjY
]N^0T1Y2BEYdE1;o<8`Xg;=@]2QkaQnIIFQfO[igXff_TmYoq65T[:7\@bV843cI
YVL`AaGTFnYkn\APDcZN7?SLP3J3gpW;IaVX[GcXEedRGSGhXAYK]Y[`@PBFddGS
@JBblBBn?6=Od]Jmbg]57TM=d`kLZR;jH[@lX8X6qC7@k^F_$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFFRBS(Q, D, CK, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, RB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
FmEWLSQH5DT^<6FaObia@0B0RkbeUQa5hZ3Q`h@WX\i??h46qgM9TCLR564k\?g<
oE[N^mMM33O^36o;5NcCK8JTlZ7BjAg:j8f227WpRm6>F<?QcYNVbg?n7^Pf^?ad
^?\09[UPA8\>e?Zi[RiK_a1epDhO]d6p5F\BUVgNFJ8kjkBV5LjmIF0ec^qVQaT:
VW8P[NkPX[=Gm;4bJHndKjC4hjn6\7S5kd>>Cj;iZC]g3OXjcP@dQ9g\cEh7>2Qe
l[j<AT@@EgqA;]IVcApkEcfBXqCoIFkMg]3Y3Z096==6D^2o`6Lode]_\Qa9OVOR
632@24l6Ph1V<h^fB@U4hmdONEWEJWAOLb:k9G`\Xhm5VbLL6aHjfLjIL^LRc5aN
U@IP3@qod@lcef<_l:hN;765PmeH:T>n<P6_;LVjefnZ<7N_2P75Ol:?LjAdHlbi
IE[IFQ8o2@nc`InIGGTnMYVW0g7NRdJ9MI8@G`P2@BoqhFBMjlik?Z\GQ_NL1MbD
U@i[JB7PiU7RI=_pg8m\;dpM?<k]lVlb7l6V^IbXH:BnTEbH1`HAaP4l06_q=9fE
VC^gF:khlKHDkAeU>]MlZJ2li>`6C:^pE4_F^ag=7RDRA:]0o44B[Omf?_7@<dOk
H`4:CdUb7QC@i5JcllGKAAb8S9e6;PNiA56oKo\ZCaT5fRQIW63\Fm2L@MdTd;NN
POWOFG`@Y^K<m^_joB=TUF06@=;_J=5mAo\hf=U2qB_XG?dSlY1KFQZfL2PNkF<h
HRUc<9R9oI?ml:c;?32`T0`Ai_fT9C13SFgW2RL_=V4kPFDb>R9G>62?L9[121?5
3g__cS9]4FPVfZ?nnCLHC<@>9ejMnCdA5P:>F6@>NQYii0F]oqhbQojDp?nTT^FI
S;l:l]@Wa8W?d`3;G?Tc25dfWma4i;JLZiWqAPO0f;]BDK6648\KAb`RqoeNdG0G
k<3HgW0`oK3ik00E3EY5Io7XGUHI1;N3JM4qI?B?Ibd\_;2X2l13hBgioOS:m]OS
58RG9a]a1lSOEUD6l\<lDWDB[kE0J?4cj?j3gh\1jg]Fmdj<C7[D1F6O`SF6Ij0e
SZLof[ah^45i2o=8MEljU@:Tn06>F^4fT\A7mUKqfcFCD1pW?hALgc0Bb1i9=U^d
gWG_IXEX_];kBf`B@YbqLY<Xd4X^ebEKJ\9IJHcjS7h0ne\1jPnTghePWTq:fYNk
Nl69F:STIR9?Gk2lQceQB[G;ocVlEE2qdQ<mjeIEaTRNF\oo]j[MV]4nSiF1;iZ^
hj6d>ZV73>jSG5;jdmAKO`[UAR1n>j?n0aNo\Odn\;qOo\`2B2jTl7X=02?<FTDP
`YYO[2H9ElA_P1\MR[8gPhE>h1Gl;LmjLKHSJQBV;H_BWB\S1Oe7np>W<1PWf80d
Hhg35@0ZP_YU?1PA>9P4Fb]HV;Qg>_dbkAf5;<[kVd^4L`HHNZYe0ILHDjE:pdj5
ch9X4h_`T@Q2M>n@B?J`b?l_=WfFk1jZ@\IThaXDqE37QP;=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFFRBT(Q, D, CK, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, RB;
   supply1 vcc;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
LO:P9SQ:5DT^<mN1PclEU7Od0Z26hJ:fO<9Y4Q_GbYEIa<UkKiXKfjoQGBZFKop6
Y_Mld^K^UJ]\dTH19N@oh?JHlFednW[^k;;8KcfUj07FgkcbW8Mq3MKiR5^AoA1J
^6S4Xh21hfjlO7Ma;djMpdJg;8Lq@dX76F:SB<]P>CoKh]9K;[nKnQqamF?KMXC\
0RYg`^Jj\BIUl@44PiJa_iJkCg>`Q@\;`0O3jHPfXD5m4HA5ol2j2b8Ml[6Mm5>?
F8a]JHpoIC[``GqiEAN`WqGO7b2508b<d\<U<<dKROW_Y[n\V1QG2a]5LOJ_:gcE
`RK8;AL8U_5CV@a]];nakXF2JW_6g:MZIoR9jRW_DF67JBdl?HVYPO5gOAL1MaMX
B5pTUI8dld1:oGZJ]JEo:MJUP=BZ;RkEKH6@^;Pe3hPU8Ik[F=lh=MG^jFlIJ4eW
DagT<IVdNM?N[l@MWiSI^IEkDnAY_=Ocb9^5NojqJ?`8nlph[;igTQUS>`FH=WX]
Nf[ANai_:C@3]]XGB=PqCV`E1>jX`787D77GciT;:@\Q>Zo]>ljjVJIFd__b;f4A
h_lfak1\3IMU<f2<1HXI6AlZq2>>HI72DGL_^k_XnHBOCHJk7P4XHPO3On5BqJi7
HTeBeg=B2F08KAiXRFJ03Q01D<gYVYTXR4VZRI5UDLW2CXhQBV]KklXPF1Y_P]?^
=KUX3ob8ab_<VVoXKobce;JTE2n>18Jm`@FEWkiS<aHnn;<fHP0YSoCNRKSVEP2D
:jDMVpH15_S2bl6A^a`==213?G@>XGb@XeWP>>`N<CHTO=OT`fVX25Pmd?^0n`ec
@HG<KCFL_9[OQHY`7SMMPQc8mkOb:8`G?l2ck;On59]P1HYPOT_O]YB8;Xo3Jc?`
@B5M9e=9dkfI6IqUDLEn4qiU[nA^hg7CW^?EQUE4^_WZb_70YaEZ=E@Q0CR63;B0
q_J`4_S8eo<U\o;1IBX`OQW0=m]<BVoO5l1I:@7Gj4do@<9OH4nBi;<e^PoWOT;7
?pE7c\15i7TW`Q>dffNg=2U2ifo?FVMCCJUi@klj^ilTqVd9N[FjAORFYg1nNK3]
5i]i1RjS1Ba^2AhPcS;]KFgb4Ql2?P4Q[U2^Wc_JJ>^n^aMOL6B`NAh`;=\JD<0Z
BYH7CR9Q05Aa5jJObKM0D3KnD;9MQ^@8dPBelH^NLaQUfYo<p0fKV;^p81?n7C]d
WjNIn?QDVd==<UcP18:[@oMQ5H^mq=>OVWMdSL=ORJ58@R5XHgn[U1@0Z`OSfH>g
@Nkq?8WF0OAW2QKjZgM_jJAQ0mh;Jcl9gJOjRS>>p]R4TNaCb1BnO4BL\7lm^PM`
ic9INFJUV8JWgU9ohe_cP4i\FkEXNlllMRQSfgEP[CB48\GT0daqdi0@4b@Y7<D9
\G\DJTgS:Y]XqhLffoWnf7abPgJdQ`RB41\e4PEHcKBk086DF@eMj[@1MdD5XiEc
2@F7^`2i]b:aHkcP1I\o7SMpF52g<^ab<=9Tnd:WCmGcNA45MF\OoS2TT;ZaY4O:
BbV=oBcD5@YoV5`=aVkK]JklUJGSFMQSdbpH`[1H=8$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFFRSBN(Q, D, CK, RB, SB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, RB, SB;

   wire d_CK, d_D;
   wire d_RB, d_SB;

//Function Block
`protected
NdfGSSQV5DT^<J<aZCLMdMkIB1IFSKo`X0@\?j;8NIFUe0V^DL9U9a0?@1^jP_5F
cAUEiD0E_49LpYmJ@fG>7f2l_??pmYig==4cI9^=CL1mDnbEfG^[RAdZAT9KKN\B
JN]^4naaASB1^9YUQAa4:hfqZf7Lh`qBVhjgSAdi^XmcKN4^J2;=[kKa^p]MfR:U
PLdJ5DOZ3YG=HPD]6RoRJTm;K82H6gZla2jXQmIo:P<S]HnA2fB<hbP5S6_H<kR7
`gQ:5OOObBpXZ=UeIG2j55DH>HcPZO\Zl2\b8P85j_;a1OLQ?Y7la6^]7qEKbj6X
9GOYkIZoP7g>4<1Z3SQZMFahoIh2dnk=F3mZ7dpFBWm^:XBDIe8G1Z;;Gne6hi@T
d0X8oV>e\<0^ZdBPK]BJX6a3EhW4CTcqj1=5_IN40lH^YK88?63i0O0QJ]mQjcTN
m][9^c8a2Z@qE?^AU@<8=10<B8<38kMOFS=HKEhL436FcXfdQXZ4DI[2Vf;8HWO;
8M;EfeUN=;^`_Al=VT<N0mK=ehjB\3_dNa?RNcQ^==Nj0I@TLGZI5W`q=eEhSUEp
C>EiU`pMl7RY_N7K6D01\[gX4:Z@fjJ\[1a03UK`BPWJVfjR>JaeKEdhh6>_cY8C
8a;ZY_k\T4FD7<iB]DlmP@cMYQEoYJOn<7mS1Nal4eIbY]09fo7pjIRKe@LgiWP=
l[j6f73V8ANgiVaE^hiP?K@hDMV[OldEdaXfbHRKg_=95QQ2\g:Qm@UYqGLJINRS
En41obmRfX4W\5MWK]`Lo:U>Zd=h0B5C3YM6I72<WnCQn7H6d\GSS[P^kGgJINgN
9QMm;GNH>kKdYbOGWFWjQ`SJmh2Zjq0YaI`BaJ`??`INho7AIcL[E6mn@ELM71\O
=`DiBaEWc`g<kb2F0dl1V6S0EhgO[=9mmaH<EYbgC<^NX0>6U^l^d5SUF4OeoFZ7
;Mh\5kpcV:f64q`f4bini;CX8<2NM=dc>JYdcHa8c?BQa\MaGcpR1mP;EMIK8_0X
PmD65:_0K=b2]bXk<bbLU2qnITOc>OZ`19]oAl;a@UmE=4\g?\9YJ:kl3\853mM[
@49m8@8UJp;HF5VSKQSJ=K[Y\HjII_TTbaj?fZS^Pi[JKCe;]dhY[\E9bGm5hYXD
8K<<>6gci8abQACnEc0<FFcVm`P2<B19@GjHUN]I@hDR[NQDNRhVdXbPa\b]gaWc
NmcfMIYJiL6W3]Ae75;i=HZN4Ncg2[p\LQbMOB;^@NF[f^5KN3]2b>GWle3_C43U
W6OEbckm:ke>>7<J8ZG6^gOa<c@3ada=SW8FGTn:dV[0cTRm?obZ][R\BonEAW<R
la8UC8L=<J5R^m@Ab9E1fF3lcfTH6d4aFV@n:PkL`JQ2Om^PlW_q0VgOIhqGhUk4
ld@;ZWa;D[0J[DUTZHFGnWNb>8V]XGUM?MHP@qW_@\_idKL?NC6W6b1;;eGiiMED
5W^@6n;EY=mlbJODp<nCk0:TGKMk8U5m96>7`UW@Y>=H;g;;@\^5Q1?D8VJqbc<C
FgeVG`Yn_gCD1c`4<>HB=Ib?1O`iZPqR>o1:;`A^I=13^=aR3=]DW^JUNK_@hVdD
n@`54:l>bpn[HOjSV=V]JY?BLc2a1gA:A1QXQS0Hh6?=1oTBf:4]J_@J9^_8Uadl
0AhmNB:FnAEDYZc?[K1IMYMNYmKVkj2ljCY=Pc\<]?MbfBG>=J;oT<;ZR?mCeCI>
U\de0l\0>56MhqSW4_7ZfhgdmDa[ZeRQbM_F;bg^P_]Y1\4Z^m3F6e5^O\?m^BF2
P`i56JZ<7=WGM=mQIM=63jNSAaim@L3[2KgAiDmULM;PFbR_=XdORdjkVb;nUQ>n
eOFJDG:NE;J6N3SGR3pJK@gC;q]\a6I6eTE0cUnD3SBH>Zg>JTi8hVM13UVc:\qJ
SFkL<Rfk4HQK2p2dfI^IQ<_o_Q0OI>k^?DSmGabP\VcVX]a7UXOgqGK]A:6CJ9bN
^KN^ifF:QHGT?bdZg0GNT=^A9`aqcVnO=[CgHOT`YaC?4o5E<=eg8DEf6c_Q:D2D
\mpi^PKW_BEF;=iY8=39_lFa6@B?>INhPeSO2\kL]R7]SCQhHYREdA=MXlh3GdPB
RXT=c1<G2R:7XqYUhfn4n8E;hFF0>D:<H3L<TCchm7j`6U<HhM<=kX\\QmSbgMjI
G8Dg9UBn8S0>Zlc5h5UX`fLPq<Sagh^6Dm@;;K4n?lRo9HRLTNcjLh6?iSj]Z\c0
0Y1_`P_^f[k::YUO\eUR?97V4T1`PdBmZCBp37>g]<gRPiH]1QL<Ei8_MGkaYnbG
`^k[BM^X4k@b?GIBhnA]UfQT9C[j3<`djWDKb<afRdqAB^TcLA$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFFS(Q, D, CK);
   reg flag; // Notifier flag
   output Q;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
W0eUMSQV5DT^<9kY610eh7daB5@2[=q[JcZnOZk>9dS\A\iEbbW`f_`X?>RXCl9W
GoX:KW2had7;f=14icDbE?lpgF11OKQC[IZ0M<4Gk\=2h0GLk;B9T`p:=dO?6pDM
mi?9<;@K5dl5EUOcfCoFcB4Hp=Bm14ja@<=>0n2k8inaca[Hck6e5eCn2mVXQBFP
YJgNQnH<5<2D[GDi4VkIXBF8bcNgIlmol2FJb?Gq9\N1o>fpPbh3A<pD:cda]MUk
28f0US_BD]5=i=Q]S_?DFQi6G72?:VVLmO`l2<4Tf9Y_B1Z=b0f:lZk7<K7OilhR
c4]b5W\4DHOjT4kb9=Me<C\8H6ea=ZGK=GUq7i3`M12MC<U?\GkOBAA1FTFHHEHi
IF8eobcV9a7O7Ee:^U54e=X9DDWBqPE9B]Cp\SfUVQa=?6m3Ek5m2nA@<fBal5Io
ThF]?d6QlCq0CU55HA34MkMH\dP>BDW^V`;B5_k[ahD21ep]n2b5UWAQc0TgSCbH
j8Y20m03R<033l240VFi\N[oQ@KTP<MhW>F[aDbmW:[LB3<G08mAfVPc[:l:ZoXD
@o1ch3^cnSfKH\d1=PbWVRm\Qbm30QI7?Rc3eY33DlIFVQhpNM4YDeLGmUA[]QbU
=:XX@DeM[SCCJ`i2aHGAD5nf6VHb3Y700_ld64`oUiU:X6KO43]QSTi;4ZhUY1Bh
;5E4YkDjd[SNUl;L>;Ln[c2I6?iTRd9m9PfI:VNg4Y^Dl?k_pZcXBFYpM>[JW<Zo
0VJDahYaV`P^gK<n6@0\VcMbY7Y0BRqVkZKlVjl?HMPJJCMFWFiZDe1R?Sm\\ICa
1ZXB6q[;a@YS`WLE:d[:MTQn`5i3qTbVLJ0i:Y4neng3U?hFCd7Bmb6bbebW2MI2
R^lj1^HUcb\DOnV2VaN`^h[f4Qe4IS@cW16qhAPOod95H0_Z@mmLTAZ6M\K1k18E
>^7KZfLnSY5fTBY<F4m9_HGQ\Q\1kkjgb`ZiD8mJA]?5?MpPI9efAg$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFZN(Q, D, TD, CK, SEL);
   reg flag; // Notifier flag
   output Q;
   input D, CK, TD, SEL;
   supply1 vcc;

   wire d_CK, d_D, d_TD, d_SEL;

//Function Block
`protected
?[Un4SQ:5DT^<of:Sjf@6\K_f40D4dQ\_AJNIdP5\Nop@nca<hX3>1m5;FmZKJe1
?m2H[919UOTjh1HH2>>:BPH7io__a`=iqN^V@8flIblVY0Ro0^]XT9][<J32m7VV
T[m\@oUA7beZ;CRGXdKW4:Spa3o>Ejp:DmR\nXnC5:=Y\N[T\f]\ddD>OqEKQKfn
NIOm0PSbbH9NejkXRC:HSE6clL:]FAo^Y@?S<B9AA<LGT<g:ZeDioe^MW?Z3@3^<
lM37cnq`X9U9PT5k<Y[U?42h>^jXLgbZB:\=F[OJJCOLb[@=\hII8H4;K^_SdjWi
>;eq>cioHAUp`fgG`7ql>2PS`f;]KLnl859j=81?=2InBLDe>55BNVObnlKJfbK9
nbE8MZ2n\;=c?Kh4n@9hZi:ac`PkAYV1^hKaEMf\mNN1HFg9G;if`W@TYA57Ng9p
0ikZScqS8Tg=d?FeMBcb9OFdL1FX_[fkkaf<eD@eBQgZ8q\8FOBnmJoF<mcIMjch
q@^l3]3n?=eVb8f6=F8RY9<^QX;:iiQM09AEp3QDj]DUZk2?Rk>ITcLUVQQ`]_JQ
G\4>PEH[F?;<qk:knkAk5Yf^IJSL>?^AXBkdOYHnFm5mbE]XGp^7dSYW:_RVF6IT
IQ5?G^C7La6gBB99SX]lFlJ>\jq^A7C8@Lf80n>X6dkYn?01F8g@=UYZT016dO1?
6p4>Y]m]Q02AE<YX@:5]]n]JC9[_6]=m3P\P5YV`=gaFDP[gD7eKH]WebIdk@d5i
SRjLUHnDolb\U[MfF66XobQc\RnTflLYYXG6i5kTBFTOMS<Dkgok9E4Di`1AXKP6
Nj?I>A1jNYm:DqaHK^e5;mbg4S`fn5c2A8EXf6H7>ZmB0[E;3]5K6nk4UnkL2oEb
HUE6@ANle901WSE8OSpc]bW4C7;mT@<1a>J53IB?`MnFef=C`Q;hfZf]LgCK2o8l
kKMD_ni[\Y9oDbLhBiO>VJ:ajHN>o5iSCgTAieXQW=m3ZX88OeILfaPFnI7hT3mi
>]n3RM3dWdA6`ZP`dJHF5DUa`:Dnfnp^AaD16X:CnF961O]H<Z4RGWR_ngTWL=Sj
:B0Z`eWdkoiWH99B==DUIo^1Ok>oiBK^WZ>ciT[GQY2FnREIh;?hBDVj93[dbd[n
3oY@o^_l17_YD7BhB_XZP5P9klekNj6igJ@@_XSH>5GeV5BqF@Jl:NL08eRBb7XV
eI<:ddRd^0ZjSb6\A^CXFOBM6n?OGF2i?WLgVZ`VY]def\6[FZ]C`VE3HVfIShAP
][ac^RF7Kokmb1DKoTXjA=bleTcFm0T1kEaAk7V`A=m\3oj<6P2]lA8271^\H=ma
pRjPYGBP]RlMbeDAGk\j>hL>cV5Fa6KoHb5UAb2ID4eCRnCIQEfX_kU@AaZ6TTHU
Lm\lG>a_1m?1CZ:1l32N:;GhNPE1=Re3@Xcg3jJ2[[fTdaF0L0;dN@fl5hZX19mY
e=1AdY7PK9<qaII_Kdo[5kDe>]DYVZ?7gWZmEMCJj@FXZS@[hghcVlAGNZXf5P:5
7Rhih>2:Do<d_k@cLc`UhaLaXm^]@YmPYL9h5lF@33\;mkdgN]bTDgh7M6ENj5C>
EhD6PdC<oG?1mdB>aV8WiBpKYKKD2pPkYhc7YBN9Q06FBJn1d?g\lE\m2;e@]`m6
o^_aA;g<U73l;SqeTn0j\8_cIkbe]da^Q7D;SbFKbbFCW4`hN:BB`qNS]4QGP:YW
OS[3GJ]=HlKRPTCQnkEdDIR[O?G7qkUJFG_N]ATX?WmRRVWGLJ]53YA8faX`=kjO
Q?YKS^>;PO]a36YF\ISUGd1_Y2OKB5CRlHb<l6CpSP_4E4i1Zb=c8M8;T_n^:Q];
<bSXP=YMpCOF54WQm9LYd>:N7RLX^V:g5V2aPb8V5k\j[P\oeBJBf<j]dJjlViIW
_6ZY2Wlh5c:JLM0d9jkqH4DQSZ1$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFZP(Q, D, TD, CK, SEL);
   reg flag; // Notifier flag
   output Q;
   input D, CK, TD, SEL;
   supply1 vcc;

   wire d_CK, d_D, d_TD, d_SEL;

//Function Block
`protected
DXacFSQH5DT^<NUb<LMQ>i]VCoYn:B=n]f\h:c2J7;SAVlmhWe<f4PiIp@MN_fZi
a4Xhd4ZWfS]Q\i<LDALaVjT@L2C[WTI6plH[JG^:G?b@KPXJTA2nA8S_gREJE@?U
i]TT5U3ZVK7M<pU5jNHmqIJ?dbNBk]2GMPY0HY=ahNO]g>1pNNHfo6^NF7M_`=l_
PMY7a3_MeJkhPdliOQC8[7MVANo<?lF>Edgl;]j^fg8m`bI_gOMkbI21bS\6qBXL
IgMImfmb4D;:C1[O:<B<FAc<VQ2PD;;J;XaM\[?InnO`>`mU=WkBXCG7jp@CUkIL
[qTA>LA`pcg^g?bKLckF?kVUPDkKBAZ4Xjclc8Q`V36?7m44XfXF;WmAd9R\dV3o
=SlE<0jcSP8mdL<JeXi8JJl@hnP:CfIFU6e787oEJVaPf28XP:jihqN?c?hA7^RI
_Xk9J9P0=>8NlO5i;6;KVEU3@_;PRTSd1;4MBTjD@hUcanQ64IqR0\Y@cq_hi2M6
5fKcMb98oPKSiWI0?XMINnZQEXWde[emqGU^2?Le^jAP:_nZUmd801GnSJTGjd::
^J0CqMB1OOT@A3:l;e6CFeV\m[2kMn\OeUcm]34EYSg`qGSmW7k5]D\GHhenW<I[
mk:ifO<OMnPg4[;U9p1hNVT9d5`c3j:n0;Y>SNbR3A2mn<d7DVP[0W22Uap8@HZk
kPl7?mf7_8eS01RfonH6`8ke_jXNm>6:>qS1W[XlN`5cS6K<oN`9HF?b2gVfSdiT
jkcWla?k0W:Vo:TUFVjX:H`=?WiR]g6KIUX9c6E7QCd=\UO8EHSmYan4^8<nJ84_
A<;Z1dl?Z`Ple3mLdARg^nJ^fV^Kg`a86j<fj>lg;Ef4jp2EhFD<XgeCAf48dSkZ
C4?be]f\D6Hl@Q:Mb;EBAm]5072LF8o<^8:E2BnAa;l6F?M1p:f4NL[=_9dXocQm
Dc3o9AmOB]V@PHXNRf`JVGj[=Uk`6P?`923HM[=KigUo\U4SgTXg>;F8hD[kHH05
ilQn@dW?XmXl:H9_3SCFOjbAZLVYRd>1?6eB[1OAHTT_KBB\m]f5_OnZ;lEIpBm5
SC_`edX]20nIXaLR1Al^QeK_hG^jLi]NYdY]_OZ3bTEQacHXnEo\LL6j^g<cLB`e
[5L1nDUQbbTlT@I2idTJhJZXfI9[Pl<fUHS_8\>VG^V@f3on1?BjKF=Td=]6RE>]
a6[c9g3@^XCb\p0M;ja\FGhiRa@T@2]RMPT91e;\WkFaPe8GhN>]JK1>>c3S:Bd7
agcLeL:Zl^:HL_jnW>dTAF_^PLBWP@H646in=>O>\H2f[B9NAD]:X8>mGcO\c8j<
Lkh74RcWEgjm29NK:?Xb`=JZL8[QXWJ565pZ6Pglo>cH7[=4O<a6=R2d8_k?GgdW
E]YUk4N;W3CmK17NGLl2D2UnG1iZf[En9Q?YZ1iZ_?>7Y_:2fMD8jhSoPmbYJ:mA
2_Z<d2TioA>B;i;h[57Wfc8G`AJ><l;64Ck:J_DRcA8SJpnIQPFH=J^[OQ6W]lkT
VS[VH:PnE]4ki7i=[Ci6GkC?mOP36Ge_D=EoG1d6H9I_:B12hkmLm\`^A@AFPFn^
25IT30PMhB]A\i@Zj1C\J6A3[AHhh<5dF3KRG=<P8_:Q<]TB;PiafIE0pYV9B9mp
^AAHZN@m6jP8[41BmS:Fkf5em3dkiJV5?^74aZq7E2?<Uh>aW=HX4UUW[f]IS=ao
XX`>m?j5`556OpfL8M:DCT>EF^8mSbZ?agTeHa?M6EG_Sf4i9hX?p>@d=7MFjN3:
oSi44O3KjOG1:M7G15Db`?0EhK1;]QX:[LITJjU21KNAB3enPg8kZ[gmT[Pq3Q\`
H[i6@Im3NY_D1BddUBl91Z`l7?cKXL>Em3]@L\kPZ2F]c_QS1K^V4OI1K25H7UGn
4XLWDlp85[<RY2$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFZRBN(Q, D, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, TD, RB, SEL;
   supply1 vcc;
   reg D_flag;
   wire D_flag1;
   wire d_CK, d_D, d_SEL, d_TD;
   wire d_RB;

//Function Block
`protected
mm8G]SQ:5DT^<GmMJE5aGbN:PI66f=<ilPE0A9lIhob2X\HY7EU]24CH:I2Kd464
WfNEQm<q7L1KQE3<S5>FD>lUcP8ZXb<iL>B@2@^FZ7N0jV;OD70hbAYBgU]^ND\;
eTCqX63mbBW8G47T724Y]S@7FAi=OU:Kc_PIin@J94pM4W]mGq5jH@=oe3E\hjeD
HbRK47_PHT>OCI_?1544I>pVoHGM>Pl^iC^83`[0ZJ4_U3;OBqAm_9OABWi2;PaD
e17H:;MLLh1PocXjBoUdb`6j7Ha\Nj]`H:d5F0Wi9=d:fe:ZR762ZKjWRY6QMBfd
p76^5Tm`8Kmo[CDKYG2<U?YcnDKm94LX6>9N_XWDLXfhOW`l9fjYl8IE?ec:q?F[
6hKi<mm6Bj<cE]V;;RJ^c_b=h328>4[q\5j\`RlmUeOV1N\dThM1]`e=hCF4UIi@
6XcjE<?pY9Y?m3I[3GHD2ghLD?=;=_gGF8b81Y4f0bV4fLEe]3XqR[GBJP=p2RZG
aaJ9GOQ\Y`cb\019Gn8K>_egNiHp\KLNW8;H0ZD`[?f:ncYWWXoM3=pNTPOa^Wp6
5WTRfSCJ9N5\=HX6:]0=2KQCD>q[mJkboal1LT>Q`;1Rhl\j<bf3[5>n7KmoO4hc
eYQYA:RqHNUA\jmqmD3YiZBq8m]4`[pNe@>D;@AmRWLK@cE19P7S5HD;:EQiEYll
U?oeo4D;DEE`NVJ>]C>C]D[YDB::9XE<L_a=VdU>?G3>T\d4S_<8=bON47kbUj>;
:neeS\U2g9RpiLI\5ZND:fCgoNAh4bg=J^B9B0`d6fgS_A7F[ed96SYjk7;UgA`V
D=\I;2[O9NS@ihI05<Te>a2=nH0a7Zc0W:6F6`bQ5Ck;:E5Wp<JLKKQpeCfm1J<:
_gL>oTV`?AZcMbTJGGeA2ZDkjdF604da<P7h[iAP3;^2VYd^lVbO6dpkAe0b^UIa
GGZAVRX14PP9Oced[M:85^\UJ3Wp]L4\UgRj:F;3T6lOf?gMo?MQ3m_=XGT@@\Yp
D[_dVKXNT^4>C\Og22a0NZgP7aGACB<I<RhI]f<pW^aQdn8J_E^EZ56Ym1pQLc]W
2AW2PgbGOC5c6Vf74EY\P^lJ42keonbf=qYHOD809F71\Y<KYaW=mgZ^eZSC:7g4
Bk;LOnnJpB]]aRT6NV?P>=A413kn?`aSlXDCi`J5_SZG]q28hG4<:d5nD^[Y\mE>
i6`IL31O7:oR^oAWd@;[X[8mRR9>IMHB8i5K2HAQ68XSC=IF2>@O1OhkQK29]8cO
0=L279?4K4m`[WAmBhbcLUb_6<Oh35fcIVH<3g1Ti>Y@@lPYgj1Po?6gc3XB@VKO
mqDd==CTSNKPgCF<EAYG;h16E>?^DX`PXbRj[4ZD@Jn2ZaIihR;A0he[W?3U71`@
n^E4OY>1H;VCQX43jh79V3Ho8?^];eVKLkUh2UDYF9AeISeQ>LF[hIFZ[]`oVJfj
]>G@7l5]\Q_D?kYXQ4Bb9qT6DTFU09R`\FAXVkMKmY:CPJc=V;li`HDL`Y98RmKg
EHff2KeGGUX56aG:7L^ElBPkeghR_L66K:Pk2<d=dmO<Wf<@R]^mQS4;RDBkU^]W
ecRI4=dm239dlYVTWDejIm8AdYA?SeXPT_:g[lP=qmTk8Ro^[^gYMD:jgNEkQ8;_
R<PN2Xflg8Q5IA@BAEOl7aUN2_NaG@Fd80B4lQ4FQQT^aEUn3idajJDTgDFO5bKJ
\eiDo4_<R0RVi6LPj>1g3QGLDUIOce@?^dRXD\Xd;MOEf77QSI7<?NnQ7g;qJ^oH
e3AYV@_`3b3XB70p5W850m2IVJdofAlME71PbPcGN:^Qn^7iWGN`:Q:f=l234cmE
^biY]]?ILGAfnAlJ5=TU[@Amj86`5^e\PmY5=?;ge1`iO3LoQ_Reg^?dACa=VY=k
QLd6l1\W60?O@=Em:9ndIg\@c^JO@B3d>oK6ZX^Qpi<77Z20j^`V5eP`4[<e2QM1
kPbK0mWI89>k:KSVJJWb[hDPI:K0o_TON@d4c7Lm<WEKbLHkLT?kb2cCVb>j0M8c
dS_e0aE:6Z^=NkacAgLCn_CmH`@dBfi;m6h@Ad=LnRTBk`[WBUENX^dN_lgRZKPi
fRfX6pWRfOmIqn\E45OSSQC>7`^ID7OVSLb]5IG_9O_HL?lW`nW;WMgpfiD?1[[Y
]PoBID5]IgQ1Y\lki7k8XoLXcPn5gh;Dl>p@l?DOmHEI?;RhQd\Lh70>3<nFoM<_
aPARUjAC6EY@a@MV\_?8gknR5\jIhbjfhHQM<2fZilGL]Yi>KPU[oDGSDK_QVN_5
Sl804TMk5;W6m=O^<]JATDLACfFjAGQ>?X]9J[BC8Mhpo??a;la39[?A_1ajcP^A
HNP`Dn[49oL=e7Y5FoWBT6pmb6F:?p`?n5N^E[ScblhU>C2bZQ_af0=a^GdISY_K
>HqO^:N3?fRD6oc544TRe0bJL4Rjk]fnGZ_MaM6U:pAZjEWoGYd@`ko5B0^Bcn\[
Ie2Ka\dM7]N7_<Tcp2BfSj<L8\dLkCFKDDKN^hA]735HTSf2di[cOH2\H<@lUX18
>jia_d]CM_Ob7<BBLQ\A^iH6D4lqD`kaaRi1h[^`XoGB\I6S66E=2ceUTdj:MTdG
gnn2jWl4a0Z==9Y<E0mJ6nB\bejoBN8AlIe`hCpROK`7_7n2QdARF5Ph^OANNeYb
dbMj9QaO78Td=\U2KEZFm\K??4B>lLTZo[`64bnm?`Ehjq[U>IG:IK79g1I^A`OI
?`aW;iKG^<EljofgGhZnHdd10_8`0RI54E8KddDeJeK@TgXM2@EepT>XW7V`$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFZRBP(Q, D, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, TD, RB, SEL;
   supply1 vcc;
   reg D_flag;
   wire D_flag1;
   wire d_CK, d_D, d_SEL, d_TD;
   wire d_RB;

//Function Block
`protected
5dCMfSQH5DT^<E7bL^OdYUe9p0MBggo2jN\?T^h]I:Be:o9dN?SSIM3Qml\=OOO]
ZaHPBZ`]n_QoWdj2Vp;ASK_9>K\RC46lHqnMfZ`Mp6Y5mW]CL0MJjeV5P_K_LNbR
9SHP<a]=^ah13qFaVcLoMF?=gm4<FY_o@`\9iZeGph@40Bm7AR6@7=?obRcoOo7c
QkWVJ;je6WO]k;9O@2nFC>_R0V4Ac9<N2k2i8TiNVMMHcl:XT_NF5R:pHeW=IZ9N
PFIEC7=AJhD7>^\YPS4T@^RJchdY5J[0<jOIdm^UR0LmcXcZnW5qc6b;XK4R8ZXl
o2d`@c_FoY>6R4eKg88n7>qX_hYIM2nhY:EmV?4MfHliMnNEK>FNR@oTcTiIEApD
>QD12Qq=Delo@Ci_CE<cl^iRl[J<USkPJe;GSj:^Q_:fk4L@?G?8V>3WO?Y`>545
oG?PSR>qe:m:ZOMRB9oX4h6??ZJ<gOHfN2bBDUbqV2UCclb_4?<GkS^F9=F=OenK
PdpXf^DQZmqHi`AJmbDUMKaPM^YO3AlY:6KWY9p54?diDCqNTm1BN;qLM1OEhpY4
FlkX^Gbda;Ph3i5b>I>6TSCE15WKdc5P0Z]k?\]X6fjl9L0LSF_;2jH[4TC?P449
9YcbO^026;o0\M:`T]je\hbB_LnlkGA0]A9D3e?2HSqnWTA_jJV@j`Z0X>T:g?nn
4JOIIfK]b7@obPN>DbdKJ]UB@PW8<Tc<^p>?5]c6DlkS[@QM_LKKh?@gOilTDgnU
Z[eYU8jPUVUP4iTEH\KQgjgd>72L5e=lRN>l5]cHX?P2`3TBHQZEgfoodP7IMbPg
58>aRMpnd4eH]qI]8cRj<c0o]TiZb:];3G<9\l::VoZ>DO:<CXpmj00]QSPWhd`6
1c`f9Y1I[nAiU:8nhKloJUq>k8R[9de_i\Jea604ARJd]T:HYXP9;[WC\eZ6I>qQ
akSBgJTMIdS5\3jV<EZc@\nP>H9oVCQ>BiOg4p[F<F=N6j=_8JFo=I\WJE^TQkZU
R79JX5mHNDl1O5o3q3;9B`7B?d`KTZ=ABJ7VS3=T>KRHK6SB:N8?J\nqEYfjZVZj
UAcck8fKIAHV;4TJGTDcQ[DJXPgIp2`O=Qh4R7YGdc_F7X^Q5R4VT;HCA^5LJNmV
_?nTWO_Z3OLN3lT>7SRJQZc`gTCTZcf9_WT?L2o?Zcn9F6WZo1Z20JmB_1X70BV1
67M:QHJ_^N;JYhlT\^JVR=O@XL^PJ1?R>_>D@hG4?<QQ3GQ@p54mmQ<Sl19:[oh8
0W8WijoH:B27op1KB0T@Nf5nb`D35F7R0dKAE^BX2WNP=dJB@WF`X04KnRPYNd;>
PB2aC734koIEWUSgbKM5GDbke>8>g^kfR;>KmZWKBXKMCk?Q]oEZfKF94\@<H?`[
2Pf2AHkM5gj`hcA<^QX;UEJRWSfGJFMIeq5g=4iIEOld`7`56<TjQ\]T`Sa0S6db
Y]0?=g73LhJ01e9I\gc_b9I4GKRLCHaaWYcRd2D3]7mePF8G@OOKXkk98`Vnk;Po
E_F`6mcVDDJ9Rj^U@i[2d`JOaCHZPeUCh\ko@PL13UQU3\M5DLe6p2@a<QIm2LaE
<YNQ;I?iMgQ0WODI`gVZMdJ4l9=ol@SEQa`<QD9;?fe]d?]WiOA:BRAHR8?7E`8_
JS`XU6XV\UB1ASTVAYb[:79k2XFkX61Z<\=\Hg>YD8Q2MXOd^BhdcX3;N8JJ3JG>
@T^]D4lqd]bdh556k0dO:K\^ScMM_BGB2Ybe6nB?Acm2Q<>>hQ=jaWPl3^0P1QAL
DJR3ioY:dO>lZJaRh<O891LDhajC1Jlb\F;M\hDPhMNfE_WAd3gG?f>HHM:;>SQ8
?idMPRDS447Xa7Wd<PnOKgkCB5n\`NH<q\53@03;A==T@\CW3];H4Q6b;m>\J]17
3C8?1:_BDQC_KAg@a=0AoT`d6D8HfaCVnbD?cD]7T8m5LA7e>6cjZ_j>Xn=9gG2<
7JaoL1loUWCc6ESXB3XR:bTVFL2B0:IB1klU\5\Ql<7bSTkBfjJ7OoaF:A0jepa=
nMZ]p>0S1N3nMC_gk08>0dQ70R@97Om<p\O:0<=QAd\:>FiL6IaPbPFHPSgEFa[1
5L_MlXYhGDhq5_<5]5gHD_N9XTdEOS]fl<A3eC\B7m7PSR7Kn\fZ>6pGIlM<:JgS
A;I0BL>Fg^^D=>C5j[fYia<JQG\R>E7GGUE4Y?lgNaE=WenE0cUockSlV2KB`65R
5G9KIRd96aHClaJBYmM3G6`Ij[27M5?PH8;m8F?]6D8>T<`om0?N`B[KDi<4>:gq
E>K_UT?[0eg;[a2Y0_1KAa4GAaLE:GU`6BG5Q6B76EQ[8<Z021>hH0P_bMohp1]6
C3?q8<fa7A01DUGbnHMVLd1L_U5i?LCGn\1b\3H^pDH[Mh<=@cc1g5\Wg^Cj1TWi
To0>N@gCU@9?Am=pREc9kJ\5lELDP<e<g;A;[_V:6kI?=9nRAK:dV_DVd2WL9S0A
C\XMd@I2L`EIQb6IkHqEmBOFLm@3AZUSO1Ql;i\20NAET\LOnCFWWFS[MpD8f>cI
g3[J3lkOGUT08a6JSU5gdeSZ_6R`GV;iIeGHb\]9X:gONVljM6R>6L_fgOT^@W3H
VRg?peA390\TWFR7k>?XiOWX?YL4NE8d\U_^[0Z>3@UAYBMD9c:[KF8HmhMALR>?
<7RCbcY=SnZ[<?hpBYlDWBT;8nHAZnn=LCO9i:V]:DYlNdmOZRGa5:05KEK>PUGJ
VO?ScLaV8T@0LQ<Ccdb5PB7jKmq1Um=]O9$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFZRBS(Q, D, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, TD, RB, SEL;
   supply1 vcc;
   reg D_flag;
   wire D_flag1;
   wire d_CK, d_D, d_SEL, d_TD;
   wire d_RB;

//Function Block
`protected
FS;Q9SQ:5DT^<?YM]1f51iFW\QJg<Vj[3F;1GPqXPe80LeXXPgbHFPa`<Ofe_]_b
BnNX>V^H6[OK`Rd08g=3E26WjE`OAAGn=?;V0oFp^oQa`Q`?>g7k:PD>^]nn5P<`
oL0dYcoc:BX=?gcT2=Dn?AZ8>4QF\11R3LPpShTWEHq?YPMkOBmU\=5Zn3<FF;EP
onLE8eRjgdk[f]6plT_hcfRgQLA30SE;E;m8;n8Lglp@D9nARbLSgbP6NoZV=mUj
><5:ejYeQ]co<9MDSdknSbQfkL^<Gi@bm6dc;^U;kd6F_N^m]]OX6?S5Iq:eneiN
CUHmnS]1Mb@H;K^b4PphQHnJ?5oRnEc]bP5D\1^;9m<X28HG]E8a0[o41E@ac]Xj
3JGP?jd[CB2YfUqLC:8O?488kJF]BQn7e4bJ[?8>609PX<AUmpDTS@n1<hbOVHW`
@]H`nSP5i23gP8\EfbaTYmjRop>^HGBOAqIMF?iE@16TXOlHL:\mYKJGXPbdBJCH
lp7^2NN:61KYULcKng<oZb43f:ZH>K;5CBPFE7lIPJh6O`@94n:b;e\G:8amGoIT
7IW`DHCMXp]d444HHf6\<o>eFK11Z6bO5l_1pCK`M]LKp?k[c^4_c]RG<DC:iWge
P><cUm^cp;eoZX`XqQ]MfOD2p??f3Pnq0gb5MUQ]EA1;W;e][TFE5f<?8N?`UHk9
:PKF[IoK6a=7:]2:m81YpEKbEA8?c1C^UAnJNWEEQSiH7N?WjDAYnn91iSl5HXnE
6De0W_ZaoRZEF6g0QThP2XD?>[:ZV7];2H8;BQcmP:FBXUja6l\XIhWmT?c5NG6l
8q5?S2?k\jPO<:1?jOgh00jg]F^djVJ7S?9\6=OWA0@e`L_1@^R92`m;EhNK8:;;
XW5AS2?GlZcmgZIdAkPZV:7Y33TenYf1<aLiL=p80;eU@p2HPKHaWRlV@AknMh9b
6Pb:Nb]Ld@;n>>g6_@pB2Ef:C2WG\92QFUmTbD:][V=1;OFfA135fDq>EB:YG6\=
V0GJGGb5_Rb[Xc5Qn@INRSnhdNo41Cp9FMl4H2TaQ@\OIB8^`JZHGO_;RQ1K5SCh
[3oR;pkc^PkI6=7FoZRBPOK<CJfAg<_K70l\HL=5mH7kpTj?^`L7Cfbk7R1=T^Xl
`llbi1H]qfFkeKfo1`K?RoU`03X`P?NQaIZ1P3SSeDI:Qp7XbeHMkY0Z@B9U]HiH
ec1;9[FOHQ0\DT_7[KBGS<cBdPPn<Mle8b:NJiEoJRDB;4bml1nS8UFUjX]3c59g
en]MZe4iT>@3[\N_fEQm]kEE6_3jY??Kd@34KM5O1QO`hR]kd\PUXFYGUP`On\]B
gq3n7``dKQ?2`5J5C33Ukf<l:1A5jAb?VD9=XOY1V9kB]3^KR]d5JJ=j5XcDFcm3
ocA3d:eYXM9nRa<9<?\5k3e<^<\^4RiF;T96I_?hh=B1@\FfIMK`OZJ`LBIXB>VM
F<XmPNVB?@N>iU8fRVkADp4WZfoJTZPiN2kmi6g;XGMlalH0DhMI:JZgjY8I[bZf
VX5bTielT0mEpH^e5=?c=4BbF=4AVBRAI`VXA0>ZK`@F_IOmQ5aK6>;faT`U`@49
VHA_hFFG=Mil0aolj`Em6i1\PaL;BJ5FJ4J6N>Xe7N6FgC=\\?\?B8[89XFC^mcK
Um4dBF[lm^K^Amf:d_JdBPaJMHdLS4`qHGIX0W_E1C`ejIWJ0CGW:hLX10eYVCK9
O?Ydme93DX8bf_bd<08h7[G6[K3Z>d;mYSeI3QJVNG__Y9Hh:kXl<OIPR7hM]UmS
f\MH<Jol;f@_n0?jSZmXgI]jf]ZN^UlMLFhOZ4UkBlc8mn^iHdp5a;>Ek[Mi2T:Z
TAm@j7oGEJJ>8PEhFmZ:]3JjQcGnD^QYifJRcNWV?@6LGaNa?7]5=W62^1A<`akQ
1Yk5d841B<RBe@jkl9aIZGMJPjGNUkY2<I@?WnI[VLJO=fH4gX2<7]ihQF0F126i
BLPl\b05TF4q>S7H7XBB]ikGZW]@a[3KoB?X4T09gR=fDoARRH`7cI5;CIPGLGHc
@KQG?Ugo6UY9>cL5bm0IC3[RebkFWHlK:Yo@eNYmBF7gPM=F:cJQ@\n:^<]QDCla
JP3l7Z6?Ee4_4gM1fDPjTFbWMI@^6beoPj_DQomipk<fZ>EqSXLaV__f1nU<bWcH
jEfUM9>;W7o^UY@UAGT0`kRP02pd`H__ZgaSG6VJScY:U^NdH=J9l`@C`5RQjTJj
g_G4`S@R_KBQ?Eb:5qbcEZA5QeRaPGo]BcSoFMQKB^736F=F0eMS@^Ld6b=1qaS1
Bo\N?82>LLHjPm_<mWCL8M@jFWXbHcJlJSlg2;?6i3k>MF1^U99dbEgK\0VY\AEi
fGmRA5RZW579RZcRGaTVRlDAZhnJiN2BiIdo[kAl4<jCLZ6<OeP@8Q@T5R95Z4PB
BFO;MpolUNKCqfQ41I7cVO2P]22`FXVL<?m^fL55=RW1:I\O7qJCKFiX<Z]CUCVJ
6M`h;OP\kEJQfC`3Tc@G@X6Bq;A2gMYciaUh@m[oTfNk:khhe5>KTe9d7e=ZTHCq
K^SY1_WN2Zo9gljEiQL<iIO6jdn29H;179JheY`\P`L5TJg4bNQ@AUjCVIZ]cRnV
Z;4oFdIK__qh?:jBgLnIJQn\T\DnE94XI@4e70KEAjHdJF]AcCcH9Hj^UAeG5c1I
FnG>g9<9i\W6ZcKaeS;a^q?e3i\Q14Df]lc[_9[m>=m_eA6QHQh5LcnhPjk3ep]P
m[a]i?8Qn3cKl83FB;2cQP2F\S90Yb]`LRI[0@IFI8?8_G2WTO;AHdhXJ15K?S4e
UA96pSZ3nf4k$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFZRBT(Q, D, TD, CK, SEL, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, TD, RB, SEL;
   supply1 vcc;
   reg D_flag;
   wire D_flag1;
   wire d_CK, d_D, d_SEL, d_TD;
   wire d_RB;

//Function Block
`protected
TOL4TSQH5DT^<P8aB10SZMl^QHkX2<BM=bI=3k^Pc]B7>YV;gh4q>Q1i1K]N;;dC
P8ZJ_`\m3kD8G>`TpL_oC05hB^0m310NS6WZ:2LL4@07iM`?9;>mpSM^akRpAO^^
YUmWl1^_hEh5?JI@`5V1_mFPh7hIF]>fqW`K:VKK0:9e0n8FHZZ8L@T8kWlq@5;3
`B>9Z:N?Pcin38a88UHDmXDb5e]3_Y:3d@IY1San@5MWaPHYcSjWnDlRZMa4=iET
dfn1c5`Ph^plL3MTU5D?7MIo3Q[:DhbeTTH48D6fjaT[ojbii6`RNS]o>K;\Mk=Z
eHYRmUqCM_A9m>_J14IJkbhB0[S4?<]TPh5QLUa3_q\3<]Me]>\XkaiLcRQ5ZWDT
6e`0<[?IEHG]@<Jn;pCF<QgB=p]R@M^370X\i;_O2iTMThiY5EM2Y25nmqZj0>bJ
lZJD\E`TL7D\RNfld7O]aeW:jZMi_G?QM3@5FIGL<epG;dfg1U[?j07GX3XK^E8:
0W3`<q8fIeFncqbmB@:=T;\SDal<;fehVaUCbBN`6pN^@XdFlpbXD@]g7S3gWZ6\
jO7M6=o>=Q5bMC4_3=cV1f`X6AW;GdPbUJpJM[d6V[p0j^Y^[pZJmcH8FQa5>Ff;
HPYF>_YdS`J_<T\:0oAldi9RD:DRb3>AZFjI_Sfo@na0a0MGUQgDPohBSn]RGB1\
a0]NVlNdmC>HB<W8N0h>BlQImiYTBgp9>V@ao@G:>W5Q^Q1QaYMK:beJUKMDeHKL
FKQ00>okYI3kF`K?RFOOcWlQ;HV?]]fBLcm0[0pZ5]K^mM\Y:dU0WV7kYQ[M4?Ba
TBlYgAPF@?fiXNB=jYBoefB3ejQdI5Ik6o0Q`NdZ8]_^XL9PYgC[O]N6Bg=A\97R
D^2>e1\M:`8pe?gI``q7\K;OY=R;33>]XNg>5e84gY7CEK@\GI]3b@kpbZ@<mBKM
^TbJ=8P>mTi_`dK3Fb;gMj[]n_YqTW\5E82^8K4g\`eaabHfiO9YZc14@=DhhDO=
@mZq5MeW6^\2DRTJ@ncP4^Q]7U5ah@I]coYS^02cl`qa[F=IJUCD`<>WOVLJRXG\
:PlEPLI?cXh`S0[HhqL^?h9QYI6hBf<PZd`SQcQ8RC9^d\ZE?L_hgEqTm0L[bR:Y
U82?be7V[F8]_]5Vc[V0<[PgD@@4lG64UPPa5pW6k82OOXgLE5kH`0;RMFa<EOLV
Jc4;N8E^HK8]`]12hOZbTHOc[JnR>m85C<EMAAEcR70>8]>MCnMQ:?hfT_16?NDX
S22bnQKS?L1;e?Y2Mdf8@3OXUFUW72m3cDXh8GT@jFWY8F=\N6RRRQNRJq0?;lJ@
e3hB5837h4a8kQGHP<QkK7`[Dln25`Jh0kBCgUSg>cU9mgPV;9=1h]QX[0736_<_
[MEG^F^:FAHa^2@15hOoZdE0?YH?ak\FQme^<570YedgB6TmVa1bl<WC04Hj^4Hi
AQEM;Yef0LWAepX4COY^6FD_l`k6aM:Pk3[bD7QNEWe2DheA1@bejFC=WK>7UK2B
2>XUD_IY;c\\Sm[PleJfJ;eMSU>ne]G>UjMOA:AGFWF_K9JQBa2PXL;K<6o02]66
Hl\G_9=8[0<FD=l\9QkTL0]`^<n:QSlIql5>VnJhfYF>J<j63`IMhGW_317IaYM6
AL2b6SE\>@UFQVE_cZjfImlb]TI?:CP4qaC5E:HMlU4ldRY[0\RefekENUB;Hi?[
a;JYgDcD[Lh0AA^FADN^diZY:U;d;S2]H3Om0NfGFkfnmcbjJS@S1cJY7YlmK_dU
6QadY2Smn4;4nHb_BFQ>QfVMn[^O;2>NS>0M0]noRQA<0YgJ41mphFUXFSCfWcZC
2Vb:E]odX4Pb^HI\UHDjMXCh=[JVobWb2CCF[YVbX9O]e[hXH@EGhElJeG`^\OWM
`K405a2DSBIZCXN]L@=]W<kHFdYVgG2d4^JT]N2X;28hG@Y;;Zni2mHYi4J@8VTM
=Of[<1<4[LXapSgl7RJ]B=JkmS9M@8DkF1a5[Rn96iW;Nca3DOL[RAR`?PSG]k]8
nedND@:N\;c@HdU42OkN25`4OkfHl:=fCV[Kc6PkTIDTmGL7TM4@1<AJheH3@hK7
8hhX]Hk<H=B[Be;;3Ra0iSm\egF6NhTkg^2=]fHSlqTUc@YapQIKPKSUC=DCM1fR
93b9ZZVDBbmE6cB^_;ljFY;V?8<q3;M]:EW:mK:Fl]Zej4jolaGIB1Q5>QXfb=;b
ckj6Wgpe=fI@8l\R8LoY\7a\BlhbDLb_[2QPGTcJ:672G6EkCo<G5C7N:dcW]mi:
[=XA^l7A08]YJAQFhcVL>\aQk\\XFi:nXUk]?GlgYOaI>HDChNe4=KZWo0_MR<G^
B@C]G_<ah@^9E6SqHlD8h1D@@NcQ58K@jXPJFOc9AYJc`KW\AGKLbM1C<^P_Y=3J
3W7S`oYCU\URb?3p7OUR?6qbHA_?jh[aVVSPk;<\LO0NTP3=KK1M79fcHjCp9V\6
Z00IVdkD2K[J]?ZUJb\^:J1n<oM68E@gkdqaE`2kJN`@AW>b9ZQoL3Q>FE\Q9ZK@
j;e6be4T6q8LZjY<5H^@8DNCWDS8\KPTd5ACj1FS[AFP@?jj7U=Z7N]EVj_Fji4L
9O0lbdO[]9J>I?DeWb;SpjZR`gLf6_7\Z3XnACQEi1?PlAITC1[c@W_1i3VcF1TF
iWCEB7T5P2kR_n3J<_bo\8BUZPI:e]Xq3kW9jRUhj1gWHZLZM48iE>G06<I12h5c
>S;3Ien4h6V4W7QRRBm4B<KQKBXJOnjOSCDY;LkGbJpTVLXWA2o>JCh:VHi<[_UB
]Qnfie95CV9S;be2g3jgAO<L^2FEC]fTdmMko<qYgDP\o7$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFZRSBN(Q, D, TD, CK, SEL, RB, SB);
   reg flag; // Notifier flag
   output Q;
   input D, TD, CK, RB, SB, SEL;
   reg D_flag;
   wire d_CK, d_D, d_SEL, d_TD, D_flag1;
   wire d_RB, d_SB;

//Function Block
`protected
lGlM^SQH5DT^<lQDK5kV4lTSX4=?G;37_7=K^g?]A3S5_bSM_NGji[V9RbMB7FFD
q3cC<MnT7lN6X8jB[W:mq\NIX^3Va`C8E1R5gQZ4icck\Kal1M?h]d7_2R\ZV4f;
g6M?XaYSj\oDaaXafIkIIIe?W[dqdKIV8Lp[5`kC@]V`ECacAV:_Ud2YLY4ekiS`
bgloUagp[Sf[kEDQ3e\KBHIeo^hMgI6Ti<p][L9Ofh8Z]R4eYd[TL5Oj?gOMQ92a
EDODa^P>\IT9KndS_QF4SRD<KQm4V8Djn?S@:eTjgkYjf9=lKfqAS>mLWAaIoSPB
5EN>WUkdBTGelh>_fRYVXf@HMWb`C]dMZ7Ubmf]WNXbD@iq7@i^AA`oHO7NmFCo4
[6maXld\aPWob0b6WKZ3chVP=GDE2qcG2oJPlA]GGL3k`8IWG`jE82oB2nf5ekXG
=jH;\gE3U2pce6D:\Ah=n68OOVMAJ;RceNK:@Q98QioqB7O3TE?TO;XWKOSTljJ<
?H@Ll9\`k_fk5^63R??^lf`[?69[PGUq^`032`S6j3;c:fn`<5MlU^l=lJLPDnlj
Pk]3Fmqo2Qb=B1qOSIR][D0KlABW_NlHAZ6gdNN45S?1n>qc>oBPYe=NHhbFddU9
eX8d9h7dIpG>V0jjDqA01f5N01^43cZI4[2]c_;HLi`AOe8h8hBE@;j]IbB9fO0I
TC7aMM]@E1T3?f2Dq5DPF=MS0NkJ^::fLE:nAa5m6d9MqKn5Um_UqfJ`^M34UfOe
XHcP8g`\0Fh=mJ;U6T:WU5UgAE=HR>an:_RNh<Z0f580LpmVi\J=D>il@dIMbGV_
QUS=`IGGD0aTnF[UEIfj_=gX8<U<dIEbpOQLI:F5jGOfO_[IdnEnJLjUAZ=;W?2@
XW9Q\]OnD=aQg7h1]cO?7dRm`lC5W\l@A>M4X@M56UR@L3><=]Am4X[YQ5jVBGk@
6ChQ@15nhRVNpDB2HeaEpCSH3\1pHCg=H9CDSAXWbXI[7^i8Q4XW`0EiC3CAe`Lo
VD\^<0oD\8jAe3UhM5i64^n_\^b^jT``fU38hX?[OeP_;]Q8Z[3:VgonlElWRTQ8
DbB@3=I^pg5]b<V\]A]>0fIo\dGo:]=6gH=@glLO>Z45Un[8DnXNaM@A\W[nRfUC
;kELX0FheSb7Hp1GEF:`ASH\1gU4OV`RaESf?iAC3;H[1d2jC8a5kQ??dRAAKe6i
cKSJo7I0O>;okX>WiNN=L7KYFMj4WR8TLP55Lj<Cnma9W_5Yo67L?BpM0?Yc5A8V
gc^`?6hN;U97GlGA]1<d[gW=2Rf\dll2mk9mOngjcY9aOBNlXnVW9IMM7?GchS]d
Oha]HB8XDiS2][NJ]49l^SJ8[d@qcdb[IhpB8390XfeXCc`3\LRLI7hKIE9MVH0\
5iab_l5pji4Co8M;h\I\I^H[b?:G2<n4PmZ588V67GLpY8ni\QSI1WhYII?fIYec
>jK6oiH8AJ83miOHS8Npf=<Q@KO9@kX1OB36WNhVe]_EOJIUl1^lGK:WH=qMc>7h
V=Oi:@V_meB2EC^i>m`Z=Xq6>KfoTb0Pdd_@oL<mE_90YWm^^4meO<8N@SikYq?3
;JXcoC6ZXJJ7LgfYD05gFEIR8`THAeF94FqSOn4YFI<Y[ieU;AME<cRU;HW??G??
k6;FT2B@06IY4hm@MnP`^<gO:P^Lf7jAS3hdFnFc`S;bOHiMPJ7NaU3EZlEQcEFO
`IOoA:;62:Q>O2<jPbebgoRcCZMJcf:oWA>IT6VFOOTY[FiDYnKM1]Wi1hJAF[II
[:qU]=I@gA0goCJN6\Q2`ZL\Dh<R\YYi:IcU5PF[@_;?:a5=[4K87XVUYV0QRVA_
YCK>bWfOTaKPnU0B015a2<F72=j:5O=:h@b7VdOY7eHe6dFZa9SS?UJ1n29iAA@o
U@E];;ILP5ZSkZD]k^_=>g[O^]7dI3MQ=\UK;JpOh>Lid<]CGo_7AP[ThT1`FcLm
V:5KLG2e7CVdU_SmIB06m^J]2DYP@;XA3^@b4lO^@K`^L80f;cU@P\O2Ik:m98k?
fA28Je3b3HG[hj;PfOa3LXC0^89SJWYaEi=>0CIOiC=NAinh<G0nbX:2o\Em7>?G
m271cq27?2JnJjCD9gPKfd1`Fa<dS]:L=H27Njle7[Ak5UYf=IU0QEoP2?=_I7Sb
GeEi@QMcQ[l]]AZiOfYiiDDHSOU@c;P9lXoI]fVgIT=]ZWX<@\Nge1iU3=;12Dc6
`VFTNZ2JXPS7ZYkJME<O8:6gO`n7Xg_QGD=Cqh[2LHfh3FiG?3DR^hSC40=9mIW^
bT[0^U5@b?DM0`9`OMa1`f0h?0U^c^VJ;mIbIh3<DHD1DZ`[YZ^^L:eJMmNH@G1:
NhRCJ<]Dc>E5>m2?AEaK\aTRo6fHZ2Zghg[]\Idei9Xc;\mXjh5n@LNb3;8gRGbV
DgRUbf<Q4pS^4f52R\ZY379QN7_\BbXHc<b0a_;i2MS=iEM5KT05T=nH@82WhQPI
YC?X2NhUhLjkWGm]OnbVJE:iQ8ajY6YZa_CJ[5RXU;e`>H;da>eCl:CgCUD>n0Ik
NL;bO=Rb4I8aAMMb@5<Y3:<XDJ:^5N5916;d5XFL>A6MSRZW<mpO1^S6ZmA1jN_V
<W9NX1eBcG8qDnCB:aq_aJD=?eI6_PHCdnGGlidRSOme0[Scgi;g=jNjX<S9XpF>
`c?ZQ8;18@gO8GUSjA;G<6Z;KSSBCg`jKgk1^4kW_pYY0[jmIC_2d3Ba>c2M[`nE
5]2AS;[<1<LOQQVOP6^1p8TSjRLcM`\3Hlad=gHdYKImol0]bhM0GAYedRaS>[T1
4K<V0X30[Hf>SKI`7TU>A]>\fDWf`qbU59J[J62@=A`WYFi^a]_;RFhQ@CeQcX^N
l6VFEE:iqaOQk_QEVOaEkGNGNO<Rf_YAT_DcEojQTc8O\k7?kMX]03Fo9\GT=:O8
XX:OQHfLNX]5:MBWN3FgfC087DLH[KVR8O7Okl0N<ASB\3[<Nho[eT^\mB5HReM@
f5;9]BcOoD2@\[i:ap0O?h=]YfIjACbcla<EhJ:d@Zn3cnc9CHMbRUL[`Zl=d9>h
LDDfIC[c[aTkNe;B5kGfgWTUX2]7C?3@?<^P\c7BE>`0_12?5QBDa:;3FHEQN[>O
V6`1ZoNRIQR8Pkc?O?D4=ElfSkOlpI`M9d6pTLc^ahj17i?HNWQZ]eVTCJBM57I<
OTR6j@Gbq6l71Q0kkc8>g?aIRL\W;Z`g`DV_<e?el@c\nOWqOV>dccABlSO1QW5\
fh\Cg75oPd3Zbb1\UIBnE7pX5F4X_4A9;1i0fP]VK3\:dGUYCmaF4Ilp9CCk<G`]
dE<QQ\kYJjk>=nDSY7Sm3eF:34[PoJpfecU>BdnbkhEKe2]jVD?aPDaXJRMNdLn`
1JSnX=0?414\[e]P^;Uh0?^f9]mLVQTCOPZ^OdYJCq02C^k4Gng4;_nmNdVkMSb9
IM\6H\0TA]Gl>kT]kP40NPnoT]\ZYP?mA=Ca0JG8I1jTTeX1UaGNpI_LMn^7A=mJ
@CfLIWiFBbF377DIPBlcSf8gD_PJPb\BIPYCG0k:ZVT_0HPkoWlNg5PLK;jFGAXq
D9nJX\i7X7T>>mSK=`MT>K7l`OSeEbQ@V`6X?e1K_8H_DPPc9B9bb1YK;5O9\V@U
NIDoa=qd3I2A;d$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDFZS(Q, D, TD, CK, SEL);
   reg flag; // Notifier flag
   output Q;
   input D, CK, TD, SEL;
   supply1 vcc;

   wire d_CK, d_D, d_TD, d_SEL;

//Function Block
`protected
MUfcZSQ:5DT^<OCl_1YEK1n9lBSH6\kg>o0UNYLoea7Y:lY9:XLSmO8kacCfgIYU
mol<TjF;B;\kEFXpQ[mIK_OTfRcDB8nT\=fWVdfh;E?VoaLk\]]YSl>G[ljZGVG0
lYH]ColK^EXk[_P733fEp5mG7=]c9UeNN962i<?a?^>TcWSi_i65>ASn=67dPB5?
gIBqB][G]OpgOGV56P=F`9`3f>T6TOUdScV8WpdBUiNQ7YBTRi=ZFDgVOi7_XjUh
1F5GCf?Sb;cD^^Xb:lL[^]]W8M9Q8ZSiC=XXolK6h2[n[_eMK^qd\KPol8[XSLLV
lGEhSklkbL8\b_?7jh>FJS2dRnbaj0mn8G^jS>KQdOl^NW5pH4g5FcLq\S[8I_q7
PTX^`n:RZ4HZ>0PK^8_KNJDlBo673o<>cZI1@UPL:bl8`IXQBJ>P4CVj93MGho1\
_IbMF^_Hj4APPhFYUI<W4;F?US>MfgXIdPhFD@RYkGApdY;LCQFMVadb:H3W@G?S
HC3QJEaRnULqh:;W0dpcHZGC:>]ebgOb3WJ6N:;N4oDDeA`5QGRUb55V=pk:knO9
k6bf^IJSL>?^AX_Eg6hbM^=d@:O9:qGD^C?2@VAOHFT72CGiR[g:Ed_UcabGWZXD
dD_8lpj5HlN:BV9kKdYR\T2V3R`GODQLQ0[Q?K]HJPpGCLY6_KGTWDIb<J^jh2G2
PjWB4\Lij1PQ7SKKVf5qbDn=K]U:gV16kkk97oY^36X`C281Bf1bja]4eBq5PldK
[d`bj8fA;UIA24kXE:oZnJKF8GGmc<hK1<7f>l;kLM0:CW2_3IWGK2nll3IlCGa]
hF`[I_N@P2Qa`>3JUjmHfFHn^AO@41Wj_:]8`K\I@cRV>gH^:Xb`j]o=7=9cbCam
G6e`m`p6W_kg<hLN`E=JAU>mnAbS`d^HV>1G@]iDY9o06@jnKI<K<BZVM8eX7efV
LSF0jL2FO5_gAI`O::Sl@h3RVOjA>==d=R^kSDJ7DS=jA52=5ml6K:^DEAZm_9nO
Y\bESO6eancnTHdN;Lpg27n[ANK1f0ZXG2bI@CFm^gZ>3a2NI_H>\>A?Fo;]AION
^DgPS3pW;IaND12JXEad=iL\lV98?HZ1aVn;>UeFBUATiALY:0LJ\J>eUYQ<>oBK
BHieTWhWI>l]a^`Ma8J5Rk>EoRT7V0=>WFYL:VTUaHKAcToUnWU\i:=XU3n1D8D1
fIeCO`Ikb;M<M@hoGf]VdB_phUjloGl9jZW>g_K_VO68h4VT:8gkEK1>ji@0aF;c
LX5M>h0Vi]NeWg1IJ]9eo\CdhOlZZPA3IRSEHF9MZChGHN<hLFf5_;?LUW3B=DC[
ahkaU\N0BUSLfR]U2@?U;a[UohfP=87@@T;1ISGRpZfe;C=h?g1@Z[D6<mJLfeja
4^iV4GC>ihVZ?9<kbd^QSNKXHI`]L?2iaLN3PI6_^_=6<W=2_ZHnRl>EfLN8Vf>[
BH^i]l?`CPE^T:4;gP]j]1dWK0F1^W_IKOeb@E01oD;ZjGW2>Eoq03K7l9_=\C>P
d=77g?IW6I?kZc7U<dPO]@851HGD05]LY]=>Noa8L0`BI61gLWmX=3XB<5gJ5NBn
Oi_k7Gj>5mmio7FT^k?b>`oh6JYkjSE1F<SohP]^3KC6GFSedTkPdVQ2\Efm^2qi
mhk_WpghK<fjP^8>5CEQ9MVH\HI@fDa^fAZ8i\P@nFpkLdo4CQe<FG3WB06dTVC<
DcCQT7DW]<`3A_\01q>A>HVXODT;n=S4WF>6miVd[dFG@02JVnAXgXI`qIl<MW`5
XnllgP@0Th6\W;J^oC68^gEcdYVP2F5cEa5j8VTZOLOXS@mUNgeCOMDmIY[nJ17q
lgI?:]]@oKKPW^_ETDNClce<<dmX^KlF`ah6C;3Rgk1;c4GJBLoIhkWo:\9>>mRV
@eLeQI^F5Xp0G;C7N=$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDLHN(Q, D, CK);
   reg flag; // Notifier flag
   output Q;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
e[8ioSQV5DT^<\WK41D>=6PY>UlQRca0pCU=fEf4P\3cL7a]kgU0@\67Alcobh`1
\b3;BIPR6L^FAa011VgFX[HSqc_:Q7iU8PGZc=PiM]MnDXYMZTdGDYHgDdfQ9omp
jeRnnOpa2o9^PAcg6VKE;3mRjFK[aAJiHpba>Z=ZdbeRfKK@HB1?G`9<X9T?C0mj
mFWUO8]lNDU;C_7<_G_jGHnL1CD4EO[MFUb?>HpMe@<;=7qdm:SU@qd=We3D88C^
koE?Af0GfoK1THVoRAS2F=gUkcEiCB:fh?1ae0OXO\qDNDISjE\JI?bO]^6R93M\
lh0SW7[WgfT5h6GBYm^An=aKbk3BD3GJXZ9?Wk@jSOhEJ@QhckmK1i<4ZR[gOcn=
Q7DI=m]l:go0?Y<2A<D`64DpWIYAj5^ZOCm_kP[;H5C@T[gj7U`>CFiGD8KWh0PW
X66a?okIHEWRIB;_76CYE8:dWWEQQZO7c\1CEk@K[Kq<niK`Xq<>L9\[]IdF]@O:
6>bUjDMOS^Y9ea?j@>=>94R[qOH3cBWTZDRV5g:`Vij@:SEaLR]7T:@FV1[_pENB
dRQg=W5CBZ8JOP]Lid[8mIN396D`MF`M[k6?D9b==g\05@\U6@`JaY1AQ4ED7co2
<1hbh1cHd=]K]@kI>M3<fl2L`6D7JFn[YKHkPfmW=E=IOO2^NSRO0eDXbq042I_]
HOlKKcn9Q8hZ?c4kLD1=lBn@VQc3>b6AToCkAOB\kCIll0C>L11Z^bACkBlP_d3K
e1hR8@?6I6e\^fZf:C34j:kXbWMK6k4VU:ai4h\gRHIYf?mKXa=fJ[oPQUqj7jId
kqKDf]49:O<UKMF381mMWh7`6ecmjG7Sl@S_QEX7qDEdTbFE]f;``bf\H`Xa;mn>
7:iiY3S;b]7n@TD>W>KNSaAHGWK^<HLPcm>@mqiYTG99ocRR;[R`?X@8I^=41GHa
?PjRGaS[1VnSM3_bTSgXnbT=2n>X?7<joD;6G_2Y]PU^q0RJWBKY$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDLHP(Q, D, CK);
   reg flag; // Notifier flag
   output Q;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
bU^TQSQH5DT^<OOl2<<]D72aFcO0SGlTbIh\?C\^TSIlIIqF`oXk3E0iKfY;f??]
j[A9JH`Dj33j5`AC7M>P;KG1=>IBY_R1h[PhWT;TIHTUXkg0;Ld390cqdAImBD\Z
jL4^PlC[9:41hWO>NVJNE3<2o0i=8^E260RM5Z^gINIP4O6FmPe6gYj4q0I<gIOp
;h2NkP:MbVXm\dOR7Yk1DL>Y0dpbgo\G9NhTg7RXQMPKkJi[S2OSSZlHed_nhLXE
dfC4S[C^L04^:Z6AS7KgV@ncd`ebU\@qgVjh`mjp>O\GGaja8oj6YRe=?9?8F51<
C\WSL1b5`hh5cc3S=8BbV__Y0;Qp\k8GbDq@OOZZLd>G8\VS`T03DeRmd[Ki`87@
iQe5OjkkPRK7hn5cSlB3TM^mWn`j6kMXNckETcJlij@Cekn<_XS`jE^<HV?HE4=m
I[nR9Q<kYJDfD=gpc[`VjoF\lM@NmTk3>VD8F<7CmLYVoHKA^o8Z\9ck6[QQ`=mA
af^g:G7R3Ba<fa5=D@Z@>_1j<@H_`U?FNJnBWoqUm70gSp9N;_QNZ>`QKOIR5kWF
k]=e]YMh\_S8E^AF6ffXpd_=NllO?R<UbVam1gIAU]3IIJ^iV2;1eJEopJdmDC[A
E^A5obb6E>U[I[DQD[H;^S0Z[@Ck7\hZULabm?[gQ@6ESPSQH70g>ik[fEEb?FI:
ep2`Ua0A^aG<T]C]Bbci^Y5<03<4cB]2=^a4UI;bX6ZC]=DGhog1fgn:gI71ZmlW
lBXPMk6c9Ko<L3R\TkY7_]j^PP>Gf5@f3`HkeHlPcRYGY3WIMRClo=e4KRH@S<5>
<LpJWEc`TW13Unnho7d`?o55>@nGo`Bj5TAUYhM2_0T;8LSlf?7ld3oajjD6\BWQ
]b0M:c5>Ync9Q<PYi@LFa5S:RX??7W4\]XPNa9Z6=3_WN>Ll:H>O?`W0@g]:lK9l
6Znq4_7]:DpkD>C?Win3WQ0OVkN@F=n?ejKoH=V3lBI902FaUpoCVdmU>Ig7G4m3
F?\db2AMUFS8>9S77PLj8>B[1B5OMF`]=bY?\G;TMRX0Q^ZoEAcA3;ge;Fd=pJR4
2RXL9BB0?a`c7CXc?ALW1H]V3dLj?4VB5XfRYoPJ=Kb@UCK7J0?6W\WeZFYi<Ihp
XcK9^H`$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDLHRBN(Q, D, CK, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, RB;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
ngFHRSQV5DT^<`?YLDF^P75j1>[M_FT[dS^lMTDaH=^emkKFh1foCZJ9ik\p3BNF
kYU:I0J`Qkpd`o]\20aAC9Ug>=BUk9gAMC9Q0:me4Z:V<9BiB0W=BqEOL_i2qd8:
HLXTgUj4FBJQ>3^@2MMKk0GqkAdT:c4]jEXj]HdX<jZL<UPcJh3]1:HYYHFHCled
3O7H^?WJhEG\Xm5=bg0<oRQ[\mE<gmpiW1Ei3\qnM0h;Q@>_K6KeGP9FF_Zh0ccD
@e107SP<o@0k8<1BH<Q0G<mLV>J6k2>o^TSX73Mo1pf;1VAoqAXjj\7@ELZ[e<EV
=VG?1IVZHJR:gWhhlTm5HFg?Gn?l2KRmf_X7fkSiU5Ne05d3P::JdNJV[m1dZUin
@>Xid`WdIQ;W195E3\>SIVD<B`;a5pEDmE>nV@AjK@:N`@ko9CDPbZaV;ZNQ[Z;d
oL3ZW[`E?HVomWYU4OgS22Bki0gm]LEa`=Y6GnSWacR4mOd;qQ@5BNa\3VWmjeD5
69H?9K=GlW:i<a7`81]XR\_dHAB0SIdS?bTIcC5\:8Te?S9o>YmV_XKO\3Pc\CgW
?m\DgR?1p:Qb6jXq@6IVO5ULUB_eAhO?bk0aKC_>lbUn^Xf6c]Og5SpFN;:QLT6Q
@DCc=^VTaF5]FBVCdYFclX6]5=pgX0\l4cLi=WDLjB^5I=dZ9c6CNYahV3F^AlWj
OMSj9:kELWa84_<fK\8ARk2P1p?C[aKJJG>XbZml^HggNl]d629IUa;MJCTnW4[l
eQKMDZ:7>CEh`@6J5L7SBCcFQIdSY?k3HajOGV>7R6amHUaX[2[6RLSVB1WB<69o
j6RBfPf_5cS\0l]2XLHbD\BK3F6D:oCi9:pO0g9`lhb2=f@fO\b7oL?IPE=S5C^d
kgWK:BR>37bUYV:?[>[gcFnjEd2]V>FSWlYm2Q?0I8LZnPb@GU?;T?oVaRA?m9nj
1In>XLNj49aWidTY4<mfG^E>h:T>`^:7D>Ne?DEC[9VqX??AfGq1cdeBJQ\NRkKj
_GSI@:C;6WU__hfCB\XXW8`6N3<=M0p;DITCWK1`lffU<k43FmK7LC`e>^I5Ym^X
TLRom0l:5fgmTcPLBaK4e_o^<]F[8oap`=Z[T3dDF@DZgVO>NjBfe:]Lf11eknR9
IF8_^VFmkV1pTh<h2HVeS^aId;90T\>C=G]\bUVQ8Z?^Y;JA^_W3dg11X2>ZE:4T
l4eL]H^[gjoO\]kdTBcJ386EVn6icdo5XfWBB2a=7Z]4Eh_3S:TEB9Eo<^QE^<:X
[681N2p]PHSiJq:JcJ@DE0I@Y34A;X@[^ZVSRjHPg1m9;_W<W<3d>PiLGe\STAIZ
Z@M_0YA7bPLMXpbfcEmN?>C9Ufk?Tj8LGQ>CLKXUZ=eg:WE6_a:4qe;fN\EilnIQ
`\b_c[Fe>_0dZ`@oX1O5m]9mI_eqTH[Vc84mon4DX<4_4HSXn0<S1P<8GmQSS0n1
a>M=gM9BIJj51UTK:@_X6?HS6KV`Ze_AMc9>7NpOK:OCZTV]HD6O?;c\SBoJb:NW
BB[Ol;6nHCiNgDR5flW4^RJ_RZai1_FB;iaYN:IVFj4E4GEE2qCm\@4^G$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDLHRBP(Q, D, CK, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, RB;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
HJ>aBSQV5DT^<?E`X>H6KnC1PYFPa\^B4n;hIGSm9CY1HF3YaOln7bad:iccifRU
VJhRJe3fegp\X\CS8V2KXGX[=qKaT<n@WN@g8WD=RKUEeeOCUFab:i3SGkZZ[DQO
R4@=J<5OL2[BlqPB_^Lmq]Y]cGJ840i?5ERJJe9LQWdo?[lpYm4WNK[I>?O5aFGQ
`XM5<eWc]n]:28j5lQbgXM_33V?V0mD>RKfChD@e8`@gZKDZFCMMG>pV^bF:TUa>
HmDSH84Q6k>S]g37oj5URb:SS<?>f0nTJl3UdHnN7G6IIBkS<kqJYDKDQ8p\hQ]Q
?q5o:WZTRTIfS?fPRFS6XjXcbIfjii[Y@GJm5A`[ZdX;RTF]7b`ec6hBQeP``DNP
m02Wlofnno6dg[OP^;29PCTGHdG_>E^\Z3cl0fZG`VF:LEq?ckTl^RDmI<[9n@O?
Ud3^R<8Xn8OCSa]e:WhLC;g2IO8fh[@Xf>hDUEAFG`HBgY3h09`<QadQii45:5Ja
dFn23ln`1q4acYnJViQ88jNN<ThJOJYbTPBRIXcF\5QJU:@I<Z;l\5adG\Ln<XnJ
aT:1;]XK5F\]dDdTV]ZBkidA85[k>V@lEpK:le]>pMmDb]9RYf<@3=8F:Ulmm5C4
`6bnD]fWYngo7_Ap`]Z\GjmIcPl>@FPA;cZ:ReK=n^8;kiSODILqQ<Ui0c@ohUMT
O1R7_`<bZ4BVI[VS9]ej3a\XEcV_^iJg7PU4CSaKILTMCJ?8JHA2qh[daQ6IHo6L
WLbgb4ImckH_WGFW`g]Uc5Wj2FP?PW=7kO29CioYa@UiM5UZ`AVCd1Zilao>?3=n
62F@@OnVd0InLC0:J=9U\AYUao^TheJGL<]KA3E3Z:NGf>6o7co]BT=[2fLafqHk
YoNDK_=1Vf@@=k63^UddVZ1W`caeJcOXIn<=S[EInU4JAHIY_;O@k1n>XLTQQho<
W3Y^ohYl^04_`2N8K_@eklIdP>jlJ[2]3XIK5Hk>J5MUg>;6NccTn;`l=IoDWVFm
fe4[@Oqm5BbXlpd;UNK8J\7\`75WCC61N?2FFdJcJNi<8R]:g:IYf3W>=p42U6nI
9UIEK5KmCR71:cN6\Q4oiNBCT>gdVUW:\IR7WqC]BPGdE6KXOOh=6>6]P7JoVLjI
Ko^Y87R\5Z[UQJXm7=VnR[1CMX>jT3=1gn7PBnYGgKJM[o646VY2Ab^TkeKeB_lN
Jg1m]=AN5G2YfdTS5JVANFRRBCHO?hG9pe91J3=k``J]?`H:D6VKKY7@ij8[Q4:b
H=h_Uk]I5B6nnOl\A<9PCeOg\\9Y:O[RAl1^ZV^pmTF5b<qD<]EB=KlV`[<ndGIR
DN>jW8efYG_oW9L7==2m4qHKPO;6_\9oR>^oI8[m_XdFiNfi3Li65Lh@AE\VqdV^
[VBkF99bU:[NGJJg4cOf5e1F:5fG`Lb:TBc<nBm<<A`^RdSVHZ[2_OX?U9Q5GOCD
?:DBUXCpO[PK30OjlVkilL8@;>`>h:i2Xd1X^kmBC^6fR;gPDJ>gRTZoGH=RTofd
<JMYHkO_=?6kdclm_2p]lammg\CB5NXEWka78WZSj0LOHCLifL4@7m5S>>HW70d0
e41B\0JRD\=@VHZX9QWHYpbS9i[H2$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDLHRBS(Q, D, CK, RB);
   reg flag; // Notifier flag
   output Q;
   input D, CK, RB;

   wire d_CK, d_D;
   wire d_RB;

//Function Block
`protected
W:<P4SQH5DT^<Ze1KV3[glT:i9apY=Kik[9DUZjEe>LjS8o^8lD`d4BRCU4NE?pO
dC4XI?c2P:8a`X_SU5lU?MTU\9W[>]?=<Z?`HTNq]hn;60pIeRB3l0`3;Y[[LAQD
KkSlFbR`?pP;R3nR;TQX@N`j_lYZd`d]OCIIjecG<9Sa5UBV?Sk5@gV579A4?TGF
A;;2ZR@@48MnXQh1q<BnY9F<qAGeY8Gq08D_Bj9=Be=VBVU_h>n4<XNnhmn\l50m
\CZjEL7D`\1RIc4f7EobSM5f;Vn<``1LW54S@YTX6m:5[AflV;:M0P3Y>P0dS3EU
8=C>mbITD29cpL8IPJo^LD^;aj8Pblj3A2>6_N`6a1dH^mRO]\kn8oD2K^[RUeKa
O>_j?EX9UCIX@2H<EcFX11MkBKc3Yf[nA8GRnoPpIg_FK80CcEDfWM:GcL:a?`dR
OQma@DHHWmPd@0nZ4XkS8KCW^R_S\bY^h1AO78XU]aYI7G]WIg\R:Bd22\JDUADq
o[n6F>p;2PUSigTEe8R01jQ6Y0imAmYT_mY^hP687mJ6iTff`^ogha^]i4ZpF[17
llO=8bj]V`MFibXS5kMOJF?[WEJ5JON<WXqRK1DVd53VoeKI5;0f7P27=`2EE_]C
W5a?0op0S?nfnR_cHU=V42U9SVG2O]b`2ZCK:?FhONG1R1BYBf\VhE^28GP67FWN
624Xg;ZCYkCehlmJ:n[X7B<nmXiHhBGFd3USAk2k7Ie_L372gEWnLRWYIP;U=a;c
Ncn^b3XaGlam?L[pOm8iQ6`ZYJm5\]>8CU9KMe7a7W[gF:k@flYM409;;]nWOn;5
84]VmUaJaGZd1]e^A]1oLCIT4Q1JH\?J\FkE9:3G42IX\>kTjk04`:8ckGQJE4UL
a__CZ7KDb7P@;cVdL70U@TcMq7iR0ZBpek`^5gLA5[Un_AcoJA1A[T@]T>7YO4NA
mWFJbnkN4H0qgAe9YQh5b2R[bM>P\YcRn29P>_[a>S6_A5g5=U@:oNIqQRMLM8=M
BR3:Mcj`5W3:2>d1Qa=o_8oP944P]:Xd\H3WHDME]@heOdAInOh455cf=m0ACB;K
^eTI;M8[lR3LAf5c^>]G2<Vm=C1@;1\f6j=VMZVD7CkmUXo^?CpgB0oEhpA<@jk`
P1KKHbC@Ti?kaB5^DoR`Wq0?RD:W7\7<Z[ZSF8Oh2hfJS_9kG6L;h\Sg:ncNqF^l
VRXGN@nC1kUS[Fc6P]H0N70:cX>`fGNX@`hqFNdP[F03P69C;WaoN^@HfFoF]\0Y
d\YVoL`3IWFkFdW21cHcMicM:agcmXHH9>nQ26?fDKhQXCq`o4\M7Ai^eVWYIgk2
4B;kVT4QB2kh\ofBjY?fYkLf6D8FgChY\41@<P]KiiQHF2I^9Ml@k1O92p?]_:EK
g$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDLHS(Q, D, CK);
   reg flag; // Notifier flag
   output Q;
   input D, CK;
   supply1 vcc;

   wire d_CK, d_D;

//Function Block
`protected
Uh79XSQH5DT^<^N:Dd4I]=dPf`g3F@8lmOHnfhQApg<dVeN;36G2I26DC;W9`5h;
mUoTWCWjUM58O3FTj:D8Pd5cSEZG[IbSU@`hWn5O^WQOBpOI;Z^c9@IT66^X95Qi
?3a>:JX3`X_lcTi`XUiIC72?fKRMEk::@kX[M>SefOoFPmj]Ecp1NIc:7qAe2ea1
93Lee``3=J]]7YCKaTDXpeP9O7KMUTS2Cbd67DE;m4SbiJP;KoJMPE4:?X13Va0_
>_a4YO?]PbiZR_@hGbUnGe66BqX3AeakBqQXhYCopL64B@g8?l\jSNSLEnIc\fAj
b>32G?P3^R?n\j?c>CKj<:iRZFiMG8f141n:j3HJMLaWhI?80DPJXZYaT37`]h_k
SG0`fTXWhI4VDG8QRmK4lp;gfZiIkJmi`P;CKEHfj]mbCjM>DHBMEBemM4Ce@ZH>
N<6k1i`aX^?fMkk8?XO5[T=edLZdQEEUNl1@hAL_TDnIpgGAC>k<bm;:gUdbXR>1
XOC;JWTg^_aL_paYEWXlql_e6B4mH:k7oDgU1^1jMACVb3^kln`4CcWMTRCq8a9]
e;=9DGT@M=6=0H[XB_oE7nXR=m=iUgCp][bel7VgT[S74eTVDVE4DA@Cfd640RAf
C:K`C`S;BbSP2MlVZR3TE^^OK9W>?]OnaWejUUCiAdiYnfM1k>nU8\mXkiP?0R7f
Led[RoNV:GReBbnCNb^[S]AW9fFaqkkB<Ub1h;^32Pl60doldaoS70BQ;KdbDecc
=PMj]LP2>8M\PoGP?R<OKX==nC_C[eLI9bLggbWmNl@0BmV=?@4oWjknhH_5g2Ze
k8g_3a`a@R3dX>9c=D;8?ggXg>Aa]q`gVNh4q`bnZKQFRgU7cMkIE^FKcK4A8U?S
lNZDV542`aQq59D5D4;A]KhhUR:gReVHOM:YjOKoU?>BJfnEV1UnhNB8<JPiS4D3
A<\DJQ3p3Y3M;_FQnfmIN3nYW=o3ihlgZKDm7\7J0LT1i0?A<`mm[X<E;ll?`9@j
LAhOC<`M3`8mhBqTG=B5K5$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module QDLHSN(Q, D, CK, S);
   reg flag; // Notifier flag
   input D, CK, S;
   output Q;

   wire d_CK, d_D;
   wire d_S;

//Function Block
`protected
`YEeWSQd5DT^<=HKSAW7;N:`^MB[ic?4ofdK8MSON?F[<K8`o;9[L6qHL9oiOPI`
L`hVW8J?kGi]kqNM?;4>]XNNK>G9h858V4\YKNW\Ib_`6PRDRoXO5g8<6_h4l\oM
06<Q80l=<b50qaJ5KEjp5BP\iNa>g1B3;4lXLOlBXmf3=fP]]ZOFefUYk6[:b1oa
e]Sc@a59l;\MeUPH8GY3j7lpYNNIZc;K`Xd1jX\>LQP<h@oHClqKT\k09O>QcQ]k
jeh80Z@d@[[XN1MqOBe_Xm=qEG`U5935^ngWG3SpT_^U\6pNN7<^mbZ<c9>aDU7^
@<eN>O;k`NGje;eEY0PEo8BC>TjFLCnCQ@W?f]F<=H<BEbSn=H:hGDDoXjncb313
lR\T>XfJPo59TWgh9i>_M@j>iRKqjocB^H84b5F2@TiEL3j@B3i5X\L2gTU\KTb^
KDd=P8ZPH=mjbOk4Ro<l5hjUo0CcdkMNcLEn7j7hnL:In@R`=epVIoD8`3b?]Rml
jb_hQ2`IZ?PgD<keI];d<6M9h9c?2hlZg:74Bg3]`[Y[dObdmiFZ[XoT;d8JU<Wo
_GBNma8Q<q:c<dkCq]`_fnd`[dUf[iQhAZ8Y_9N44PGFVgYbZY]eKBBpZMkn`nj^
f[ePihDLP6ET988=da0e_4^\M=I6mCbWOAVnm3im4>Oo;Lj4`b4\<cK5ANT0FVfq
CK2kaV\aRRb6fb6aAGi093M4S8m`lo\oR@<p?YZLd_8DY:S1L0jjL9VcG_ldK?@8
>lk0jbJd;eY7LeZaO6g5P1W6mS]ng:P<8VI1gD[MOSEZ14gW?G8>i=d=c1\65UW9
>lNPLN?JYF?1VTGCF[1P>GF8b2CfI@ck\W@LCM4bh<:qWFP0n6YO9\QCdgoP7YY>
?FUHjC[iIP_;FV=oSA?Q5S@f=Y_XkGoWIbOi75<HISGfcRe^Ci>n5C8bGfO4>ogC
a`Om2j_>O5PBjjELWR2kJ3Fk6hE2b<j9S8L\\Zf7TNkGCGjcI]_^A:m>ok0qZ\L3
?kql5c=7TkYJ9TSTS;4F@j3<CL=N4\1@CW?]f_E6k2C=lpKDBL<BJ?L<6KSaf8@j
N]<b09MFeg:K_W66PW]<Nlj1pcTXaKcjS]X76VWG?4N2S=bF0ofci;EBJ5SGmN;_
=55GBLITW1Bp@?01JZ6Yh1Qa>ndP6FlOSDW`k=OG5`mWk]1eAj8i0InHl:ARlIHH
N<JPAR2SkPijm8PQBCD_NdTTUUTYMmjamS?f`Z>FR^11T=c?h1k=H:_Zb1e>]]7D
gL70DP^q>SU]>4pT1L[b2Gik3aEMm[2nBBW]gDVn`ICgl:f\kY>dXqAS6\KE=7go
5Ob49lHQ2qVAB>gB1T]oelR0CS9X`DE58eAW:3Ye;OYfV@qLOh;6YZFH[8@MUa`Y
7^T]Ln9JWm8[W3LFTMVGnnKUeGMEWSJ1`];LUK8Dmk<9MLY@26ZPog>^Yp6XE;]0
K4?lI8jUXHWP3VQKQNFn?cmERRJl?QIIM5Wf2@VWPMmj;T=U1HHFh8mdc<0jI_iC
?Vp:TcnBP3$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module RAM2(QB, QBZ, D, W, RD);
   reg flag; // Notifier flag
   output QBZ;
   input D, W, RD;
   output QB;
   supply1 vcc;

   wire d_W, d_D;

//Function Block
`protected
jDmMoSQH5DT^<<PYi]HVRY@DOWTbN:[@e=hUG37^FTQL8<<giDIa0SYmb75YC\AF
Hl^gp;0TdFV8a@RlQZRJ`G?WSJoLX_:LTXTZRZoiK:Y@?TECDi5KVY]d;9Gi4gQ9
OaQ>EA`p1Ig2X`e0Lmn]j?\lmdaa<NmAPC[7D2BY3Y[E9_4RT5>ZMiBG[KPm1WTi
TWUefkbp2[_<:?p[kd7n0HVSPT644_H3EGhRAanbF:m0d7cTREUo]DH1TYaC2o>_
WW02U_:@gK8@V<M[W^IqK_hA2O8T3IaOkK^CkZ^baU6?CU>HqHo01QZ2PNT=\XiV
2PWnF0lJdE]L3`Gb]WjH9qN8W?VGHp:D1]^6pYa[H>8YWhY824A=fQlm\\l@cF:J
@Mh@H84HQZD^PV>4AlIl9>j`QBGmR>F7lC<_0IN=0^50PPe:i\DYElTgOF[<5=C1
q3?;d2]VG59_7cjnZNDBOSiL4[6VcNF@D`4KADm1aoebg]C_FM@XDa]b2l9lWlNC
Hm?\QD;\OG5bN;:Je\E96J;nOYM[gp^_XHI7fcnK`GlQ9plEAXg?LANdgSlVC;_b
LP;>EMN8oQajHFTTcmEmDm=20][4;NT8?fHM2a5^M@k<GjNQW[k79?cNONcR^`S;
jajF?h::P<P9gP;0O;dSRD7^bipH6E<in\k8cadhBZFK<4U46OgST?6HDQ\L\bmL
nL`[Vfig@g4j^BZ=kGYe7R>N\ADJ8R]f4fNo=N2fe9`_93__l[FW_GGG<=UReJk8
8Q6nRg90MqVPno0R\6E^`]j0d=@i^B6T8A]`9k=g<l>7?>6_D72HBOS]2>[oV62\
YeAX`YQ\>]VbCZZLG^IGLSmOQTMKXE\:_9;UC=XX:CAbJHl]6T?_Tm61FGeU]DOm
ilCY<01fIR2RVKoUh@J:ni97PA?RP;Ral3H:oS\BMBM:1>T[CS9:OXYLfHmJa>2@
>\^c9kT`<T]6?O^9CfBPVn=VfpYDNnODq_YC@^P7YoVa[l9]SfO<HP;Tgl9RFP\=
F>7g;2[N:m@SLC6^F6DHGac<JqHjoAg:[Ue<7l1gm=aWlHe1o_jB<\`XO7AM6Gq=
5R2Wd_bTAl]MDLk04C]FSWN4248RfO;f<phZABND=`62R66kdCF9ALScl6g[75B3
Jdol:A]TTf[7AMP5gcIjAH8cl\5lMU?VCk]X@aJ<YOe6<AJ?P[mSWaTCC6^Kj>Yo
?Nc:nfjGQc?;c4Y9UB@@W<>h78UA3HFV[XFBp:8=UZ2\H0^@Zh@@k`4Dfj:?f;oi
NKGGb3l4l@0WBK[QObTJTH>IA=AE@GaHKC4M@KiThN^G83\3e1oNNG<n89>oWON`
5ncID^kBbF06R6STQZJ1j>?aegee5^20J84nMUJqSCX\IAp5E7VbF8d2KMZ\4<<o
fJ[CZOfP^laDO;<1>XqgTiiGZcOnfI8VYc9Zf\N\1]gLEcaOVWPH4MVqQ2S=GbQR
AkH]CD=S:4jAa2V:9:HH:NNO?LJ6n>d3;Cc_aZ>IVcZQ\nK:Xied4k@ROQlB[4YX
qGS9V2I0$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module RAM2S(QB, QBZ, D, W, RD);
   reg flag; // Notifier flag
   output QBZ;
   input D, W, RD;
   output QB;
   supply1 vcc;

   wire d_W, d_D;

//Function Block
`protected
oaOQbSQV5DT^<h=`7mcV^npVXS1;0nG[hQPl>0@CQ^Ekb?_UK_6T1HOGhg[_?0VU
SUdMdDZS422=SKRH8e5_GBfQ5mgGgpo10nfG1ee@Mj`;J<nbc\j`3XS60E=X[BIO
j:eBa`K4g;JUCNC31qUdo2FbpGBKa8:4c;1jZ7R1JVIA`9iZVNW551CO2?C;I[cJ
]Y1g`g`A<`meObLE:[k70JiGRGK]IqZZP\D;:SkiL^TPF1OIW`5iY:A:2ipED@`\
1[nPP2fm>khQRMJe^2_KW_UaH`7<dGCpI\DCombpNSc\GbUQ7BT]AlMd`YCmQ`q9
[6?ndqcLooll=jR8<ORg8C<9V5Z:<dJPkmN:5cMXB:L0G0aPm=UX\_9VAg6S:idK
@DW0;NO]`c4j@lHFPCHhj[QQ?VDZ=X1K4pM5O?ml_9Ec:eThO35Ade87VRNa8\VV
^`K`M=12IEB7Mm<ifTL=8F0Lmf>:=ejNiYFbSMl\d<SXT2X;C]DMIeKT6_jLhhq=
^LPJ19eI7VJ@?6f<TD]\a7>fcNoSOiba[1nIVJL5D?IEEbX4:RE^QRViKDf<m740
@eoQP:9nDk1kE7U_?];Jdj@^<3;SfMc[Bh5G1KT@ZhhqlWVScIoLEVbZ5Eh_I<g`
\iW=n9_PhO^o_09CZ8G;oiK1iF:k<ofkh2iLd8_[I7INUPU9AHmmFZSQQo2XNI_S
d>n^[V0HoSm8geoV;5Wjh5JPh6qLYNebPZFnbEK<Ff<3mG22<10h^1\2Un4IP@mS
@5m=R;4Oaa;m;CH49IdM8CffQDEB@[3_Pl?]=>Pbk4K0Tno_S[aA40:0PoHIcKA]
K5?[CR<3NTMmU@VMlk4ILo8VSJ8G\<IPOXC`iI>T8n7OM5:lI10Jl1<LU_T7_EHj
d@8V<^G@EU49mEWG\CT0G7M=^T=LlLXSBoW^bHpX9f54OpQ6ia8HcSMQEAEo[CnO
_^>mNUVbgKFBT@3bR`BBYZ\@NV9mTd?R;108RN2m@:WYYpTHh=Fbfc:cUZ2mNdKM
4RbO?QcEi^HiXDUPoUpoF]i`]b5I7\Yo<;^[g@OKFijF<1hSg@\cgqEC?;79H_EF
`[WZEl=_Y9dUPEC2_V1M6HC[j6J>4^Ik`?VmTUB[1cW_>RcKWi1a?AV;TNKXi^6F
MbeH6nfU=`l06^eZjFCFOW5U[F7j>9:Pi@KO^]8K@jAcEYk2>2_^p0=@Ea7HXYX]
RIejMmRl;_LnIndoVL:0;6[=g?J7@UdKUH:G_TD^MY^2Gmh=<`G8NNU_19gKKa@\
_PfZ4_]<=[9^ab_e[]GX9oUF=V9>Q8b^cOmKGGi00CknH^4f2EG9N9nqHB;gb<q4
FhD8JC[R`>ma3M<1BKXniaGV_mQ`^<iEBMiqTcJF84I@R2_hJlC[RSRT?X>Da3cL
[E7=`d[]B<]@QYVMkU2SQD?9]Adal\2FN0F?99CQjJ[Qp]5WBUmN$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module RAM3(Q, QZ, D, W, RD);
   reg flag; // Notifier flag
   output QZ;
   input D, W, RD;
   output Q;
   supply1 vcc;

   wire d_W, d_D;

//Function Block
`protected
d1JGRSQd5DT^<lPb3L`1\<ka]ogXAh0^a77phRlE5`0AA4iO;MVJO\UdMSndLlO?
RHcIMQ6[nFXp9F1M3mbU3^jOoFO\kR`6XX6jYZ_j_kT5c?R6kAB>0i6jP;6fjf2L
B5fnFeHhD?;R13m:Rmqg6I?EmqD6496VQRNaF9_QAHEQH6\1j][Y:Em1X9?b\WiI
L7P4_g3mTN:XaYTc5][]j5WGCWDkTmqea;Wi1RKB7F[Z\`UVOASd;7UM>Sq:m]k9
oGPm0c86<XM^JmacMPn5CDX9@7P5Z<pB]YI[]<qCm95LWpmRdh5XaT`4L_PDV:[\
FOWe^3lVE1^dl4>`5_4KmGHDdS;6:OCoc^eMmSo?1j^4=5LL<DdkAdU^D3QQI61j
oXT^PT3mqWJ7lAUd:\jnEF2KafGRdRdF^1b4KOMI;UH^d=X:VNB1H<?RcBSV7\nG
Sa1?HSlYWLTRRQ?F?No^ZkUXV2hQg2T9iW_Tp>GkAa^H@4knENVo=ejO6mMm8lF`
^8_nh]T<i_VOb:eSBmc8b@H^]HYm^3O3<RW0@JlH4QgD`VLLi6C1m?9X0;M4ShEg
m^Z;6O0<VLOcb9dOqZoeJkHd@CI:AH62d=knqHQ89PHfWhB4WlB<mm6T15OfNCfT
8EGUfciT1WT;CM?>M5EkQ[Q2e0c;En`XL]DFA@:Jo9^kHe:a9fPT;5J2CbPXi6P2
fagZcAb[MSm?TTSYXpd_e63cK;aNf>`86QEE>7:@]]ZMnZ]<V^4T8g1SWKdP[9K8
=]VOi?3PNYnb?IH_HldObTbJS31Cj4TJ=PalJ2Xe`YK=PfDDeL2H0QG[]UPXgaQi
TTS@MiNeC;n4SLZh?cjEKE[hE`g=E_^Y]<4idb_WC?D?fKdR?;JaL0TFW@jdPaVF
=TQogQ3Y3`3?Kab2ASdP6[S>2b]35ZIRpgB0oEnqh^=BQkZEBO_U^?N1bT0iWEH5
?HYbTgZJP9e9?aXF^B_SS6`3]HgDCmq[=A\c3ER^<kZ8:nTBIeA`=S:UPoYYTnGN
NP;q5MJPFTCX0JCCn><<N;;m4X34CN2XA:S\?gqLX`l>RFiN>W_\c6B?XOaFZ:oC
U_hD;hP7K9Df=NZ;n\ef35n@lVlU`JYTQVb]k:RK`80TfR]I<9n6L<eJh6HWFFAS
c0866]Yg[`J]bnm5g>1W`Dnbn1FDL;3Cj]NWKq@A16[6oQUg4OVnkT3>G8\ZV@99
Aj_Wfl[CSZSgjCF@_VCKike^SKZaOmWeG80j[Nc3]Cf=bR]P6NcL7U=X;IK:P6@A
Q@>196GG;h1D^`l6if@[o4J0@9m42e??1F4`qO^l<26qk5geGJ_P]D]i;LPdhQ^M
Ui1`Q9fUo[96a]YdpS68ZcBoKKFm]Y^85Hil]3NS_PmKI\e=c87Z<D\\;@lA=f;;
LH7<0`FP@<X?9373?S9:1pac=BfKe$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module RAM3S(Q, QZ, D, W, RD);
   reg flag; // Notifier flag
   output QZ;
   input D, W, RD;
   output Q;
   supply1 vcc;

   wire d_W, d_D;

//Function Block
`protected
kY;HbSQd5DT^<52lnIXIiC<[QK\TMDbhh=d>If?YX\i??F4Iq@_RgF^bD7LY[ckS
Jjm@MNeVg9Rq]gi9jmM5GfjlZ8RYI6>@e_I9JXQ=FK7``HYRkdMh_TRn1=gcUbW6
aWYNPd3PF\JP9QaIU1hq9IFfLmq<V[JjNjbB\19DZ]RL`G=DR>PJHgHB63V5^9c<
M0[m;4<SPZ9<5ISdF`862H9=bKL<2_MqB<Q53K:`7=b:DlYcQA]iRdf51:5q8@1k
?XgD\@X;gfG;l:e[Z:3IFB6mn5mA0>Zp>6iOn\Iqaja_`lp4>Jk7^jgZcoUK9_B:
2]OgKU7nH`O_aZm:UNAf22Ib`;dSH?UBa`?eWcj[b^:QXn0OT34S]hB8O=L`l5d?
BgS?DmI0<qM0k_2@^Ha\cWcfj[1MY`7JmBXM[bCe0K@O3=``<XihG:GP`hg<MhX_
WM=6OWlGn_1_7W_V2e[B?=5^\E`^Re6m1l5=Gpb6KT?U7N3PEUVfG\4o>>=h\W2<
Ie95\i3O:Y;<_H?L8?FV:]5mjER4g^3HjY7lXUmhg8\Q@^nP0Sl>e0dRl@M23`R;
0O_RdaT8:0:1@U=nbq]XDji=X]OOQfmg8F<PiLiV=Uln0b<`U7GlE1fgRW4:W`qV
^189H@<X1g];GMPMa7^LAmiK\0ooX20@cU<[Cm6:HlFhhHTYB^NGVO6Hlfl[oeb\
P^:d;5I:JLkbH??TEKX8:H`CQMOfnd>iE0NWPaHE[3<qd7od:O[EE\8ML;RCYG01
@9j2HBd@j@88fR?M43j5dDfLRJJ]=ENA9KeSFD1o:7gFZ>A36nISk@YF]EPfkOZ9
CJa`m5iiCaA8ZZhQ:`?<PP^Y9k1h38\HR>>nGZg8WY_C`1I^fO8:b>[QG5RD?m>m
lhjn1Sd6^@WIP<iZUmj9?X[[JLNN905mmiN;NO4>:cD<b;EdE[SeVGpa>A1:7pAH
2OWGl\AL9OVGPj;nldALc0<eMTdGd@P_`Gqn3QX\DcU4h[eZD6QMW8DT5gfJ_jhd
IPOG1pD>T=8@FW9i\n0JkDWG\I^FL618^1KIE:A]3CPHRRK`9LY5oo=mMTHO5lB5
n>ch9NX`Bbg895T3V[WE7OXb?nKk3Pf]VU2=j>XPT71VJEF\]`iIj`S>63Ql7Ri[
dK@7q\KNGGjgl8Umn6d2DFLQ_HF4LUXSHCEl?FikOmkZH:i<_7RHRESZTB0i9KmQ
oF0Ro\XcadCCB3mg<bI^lB8=C6VH6E0bFghaSoSe_A;Bh@lJGi1DmeInEJCAL]<a
LYXp`FZiA1qN=bo\;2WkFB^K[W>9KCk6eHeOY\CVBk]WcOed4qbka<5V3>7Dm44Y
5I\TNh_1dPA5\a`dSdK8E_p[eKo1[ggb]JIdZ;7oajP[OEKI`fZ7SMb[5Y@VlWN`
CZG44F9a_Q2gF\4604B\H[\[KB1p]]NDg`X$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module RAM5(QZ0, QZ1, D, W, RD0, RD1);
   reg flag; // Notifier flag
   output QZ0, QZ1;
   input D, W, RD0, RD1;
   supply1 vcc;

   wire d_W, d_D;

//Function Block
`protected
g>V``SQH5DT^<R3HkDL1@n5l^h\:5QQnjhUCUY3\X1I[b<fAgM`khjo4GBKbKoqd
a6RfjHa1:DBSBl[@aHPiom@TV:f5>T\aED4mE=[C<1j]6gK1GB`NnPe\[AATD70B
\kpJ8mJX2^T4WcN?he6D[G1=W`X`@<Cf2dihNFD>CZ3IIMZg2g;7iPFBhOU2?FKT
np@W7fSlpLlda1M@ko^YDAmm4e2BEPdTPX9GKD6_P7a]QmNE2?YUC8VjDN9PacY[
CGk2C2K[in7iq:^^:8GkCcOdjRG5O7_1@D3[SnbqdJJ`_7L@<d>UBlQm\8dQ:oj_
g?U]dHXMgW5TqVPR=]:QSfl0`i^fWX5`8>[D`<M]WlJKW=MB^qVKafZ:_qK2b6CQ
pdL9n3S2NiY^dNaFkVfb?8]9=@S0lg11_T6^Db^@9LJ[]5cZN76=nMg2Zqbkc_c>
1P0oKE=TAohl3IF0S[mlYASGS`jb8]8jUFRXmJ9cf@KQ19EJhIA439K\[didI@Ej
TgU]34fISXg_AoGhRZUS2Bqh>I<FLHidfU2W>aoK219k3W9OS8iocU^;V8n]9e_R
15OoQ=6I2fAe@UN7lNHTEKKdSiN\I`:0Y22=D;^FBU@V=:b1EbaqU49Lj5Ll]UP]
CbW`W@38LFfJ_JQodQ8IYI;h\VSK5@EfJM;dXW=<7^oJ85D9]Z`>W^^m^m<kK;h7
FI@oR2\ki`PC:bc9g@C:ocPYmLja35fA_oq6@mXU2C;0FQL3B[:X`X97]oJhlLY2
2^`mklB1ImKN=KbYDRa_@OI?TXqSnRNN41a2dFk7_j7]4`P^UdRJbPJB2j=d`kk]
eS[oD79^3]<l7M2`n_H=6XM9lG:[WRfaS^Ab;dE[Ie1N@<5ASSZHMB\MWH3\3<L7
dcl4o=9>1pNfE_QHX8f11cF7BWbCA[ZUa?=JCCa9FLgBBM1n_P1ec];6YD2Y5X\K
UBA20n7G=@N3aIi[dbURh_GTkQ:d51F5LTBN7X6LNj]JgE:SIkDnEMEaY537SH;e
G4f:@EL^cG78LDPS=knO?fmGFAXHgLo_dHE177N7>D]\WokdiA_[l4WUFVC2ck\7
;JRV1i7f3=IPl3S7o:JT:R?d4Eqcm<oC`G7:`U8RiE3L99hEliGmQTJIM;Y5Yi<3
ogZB_elI;W[bC1nelHD1kO:^Ag1cOF[]Gk_gVPWSH>8iYcFKO014c>Kc2YSZQfQ6
3j3K2O[Ugo=iT>V`gN5R_5L=Dfee?l`_^\Nc@LXdM[@I?WQ2K5ZUBG2;NgE;Dn5n
5gEJPdJ[?E2N`oRekR9nOXeSoIE<Egl2<2n@OB1RN[fpNK=Y9XVG1_33T4EfHZod
InZ1WENk]\lPb>XY[`>QeKKZVi?1eAL<T7R\N=l[pI`M9dIp^Xe@OjcNEmb89gM:
1R??A9AnkS3Fl?IllF6_5RTqEm6@?:1AZ`Y:OUh5`6[QFedY;<CP:kk`[3a`MMp]
IT@M]l5444N>h2mf>A?Ne_ZJ4WFgXCJ``I8Hc1hGo;b;V5;ogIRI_Xm2eX8BiibF
TTY:V2G6L9cXKngjJ`UmSQ2fnQQ:k@Vk3h?Kjf@7kH5RVJNUkd[Z;A7Q[>b]GpC=
5C@^iZYYmEQGF`bPU9Q\eL_K]G<k]G:I[?FoLHYoSV7P;h;Y\KXnSbgQXC5H:M`l
U\g_CXGgUO\@60BIn@OKMeAamfkZ0P3k^PIEEV^0VjAbGeKAa2mWg[og<@\1p0JL
B7XplMeA9XM@M=Xd3?2Zog4IXXYNdEe27DUa^aIlaoSqC3`h\Em\EQa^Ycl8QRe^
QDIgoG15UljWFZFXf\:5ce[25X^5C3djN932^[R[eZhDCUCcqGO0aE]:=EVHcMe<
\hbkR6ai_8@T^RSg66B]9AL>EZ>`_E>H;Dg;l?@\0W4EVhCqL`6La]b$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.2 --//
`resetall
`timescale 10ps/1ps
`celldefine
module RAM5S(QZ0, QZ1, D, W, RD0, RD1);
   reg flag; // Notifier flag
   output QZ0, QZ1;
   input D, W, RD0, RD1;
   supply1 vcc;

   wire d_W, d_D;

//Function Block
`protected
SY:=1SQV5DT^<i6a=Ncm]o@GBj;I=0;j:M>dD\>;Q]X7OZnM1OnJUA4EWNR5P1S=
ejIkiD0E_ODlpdDJPh2<Q_M4Vn2qcB\0HPU<F=Yk6cNiMok4I]<<Eb?PI9TU7MaS
UGnTfDj7bFmLJ9l>S4qJXFEbDqH6_WMFT9a=bR2[dA<oTS3;32LcH7D5O>HJ1=5G
D;dnc2D0IJPo4QO4HSZ__4=4SE:IAqh3OlK\@:WVPmU>HQ4lTE2fii93qni9LBCE
B2c5Y2A1B7Q^>QcQhK>OM=oiCdZ;Jp5M9?;i=RABenI5V9Y?^THBPTJ=RMca^]DO
==qP^Sb1X]pMO?2DCqC`kO0iIGdNV@D6oo[Sm4JWhdhjIeXUG[3X`GMDBWK9@`kO
hJ=R\47XP?J>VVPIR;3@lILL3mC5>Jm1Io\ISWNf\AegcJqL@D8UFGH<`T^1_CM;
P;7kEWR@cnH6J9SYH]RU\1<cTcn3clHMjB4k@oZFcJ@GjSBCR15kaJTAPTAOaeD2
GFUULhU7J<_pB<jaT_eRdO;^dX5CLbOK;0?`LK@?E5GmLI_W8Bqj8Z[a^m@;0cVj
c?0mH9;BnBC8Tm>j\HAC3jaN1CEaIIbjmG9NU7DFF]^I92E2ImP:UZ1i=T9_\fPo
]21kR9O\0cg`:PKM:inToVJ4_G<6VlX;>qlc=QU5k<RFC174NUB:m79Y0i386YP_
iP:SkecH:4fVVhJPF2`:n?42Y7Fc_X0XT[GSReQcJX80nXk1K189YX61_<kZ1gni
_lK4kYl^4o?\LLm5pMmGc0JI[aIeT^9?fR[4EXY72gC9`dYH0O>]d9agRF5SoXk_
\1]b^`cf?6dEBHRC?Rmg@bPQJPJ]X5_k=_>=:L?l5ed=]W[[iXN;ITX]GNNRkeES
fEMUmg<IiF=ngM6QM\GADe9Y1Q=nEEj[_@S@IDk7BWb9;@YV26N3eHZH^\kRnT:[
NYGACU;EhFH<enBKgMB6h;RGg3PdFqkFcd>5ImPZ]C=KAXGE;KYI\AV<fZ:117lC
d769b2:2gl6?UVMioB=GPe^bmkUOZ2mU=K?D0RAPEgG_7TgQQA?HDcYg8jWaJQhh
Q<6I=6RIjLi8nLeOS:Dg0=\0>KEA[[RX3__XEZTB[mL`k`kQni]F\3cJf5`19cNk
G^dW4M8f>Ne2a`>V_AflnIKjcJ_oJokAfdWB3emURDq>\H>3kqE@O:GUf0@LH?PM
XI5Z3KIOg2d48mnnHZ?Gobe6Bq05YoE`ZKT\8\@@flF1Ti3FV\iZP4HY_<L99h?D
pRXgFU92=>i]e4E0ChTH8ZGag<EE:@kP@`TFloAJV=KVPd\33m\]lH]DQMaS8YNF
e932ikgb^=c_Z1O@nca;h8CVg=BOJllkJ^W:M8o20o9f8lG0>`\6M>=T1YiKNQEp
=nJ@@_N^WRBi178ZK>BQk@`TMW@O=VY\Y7_>UT>l^OW9o;`GkBLd>iJ7n5\9SmO=
kSZ`c:RQ[V0TA=a_Nb<@0?R;gf`:\Z^54cG1cCYkP2C[bM:M@8\UekfI_[CL0Dpo
9Ajf_Vh1]=f8TL_c>Qhn5XJN7T47jTgna7DDnS7TKQh:SVDU2l7NP\^61gDYFIVB
ZbVpVjNb;=p8E9bkR<U5ANGALa[4MGVZ\XC>jeiC3TUPKVIm]8qnfa;0=5g;lH5n
Pb=MkF^j6cGKJ?XhLo36F8GLd\^YaX4134SXVeIe=;8Ree45>`cn\LYq7GQaKYmq
k_<B=<[2c:CmgHELXAH8`;Ti^aJf2bSCX5>P6O0NK]9Zo8j;IWQ@hoUUed`J<b@Q
TKZaC_k\$
`endprotected
endmodule
`endcelldefine
//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module TIE0(O);
  output O;
  supply0 gnd;

  //Function Block
`protected
>LUghSQ:5DT^<=HM`TPYU7daB5O1U=pn\?HiCi0[gFjfB44B5>CO7_;9ib\TJD]`
5cA4B=2mPFPO>PVZcnLEBCipfAX=PSLoi_i\7be\87K1TSGk4JOl6of>JIgkT1\5
5AJ>cBS[8YaqePF<nOpHA>DQFA5ZmBmN94LmE_YH1VgeaLpY5\1Ej=qOJ67a8D$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module TIE1(O);
  output O;
  supply1 vcc;

  //Function Block
`protected
2n1@8SQd5DT^<mjYjUfAd9jUhB0Cd?=USdJIIdP5hfZpINcM`i\AZaS56R=>gHlN
PmZgpHjQW_YW];FPkoN64XlHq^?TnXMqChbB=O\iSj>UML=`K];DN4LI[^YpmW21
3PYpPdamQiZ$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR2H(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
Gi@icSQH5DT^<d[YKU]30HY]5=0hi=0Q]`OF0@J87<f6UAGZWe<f4YM=qe4;SI16
R>C6Y;VkLFT5EVm6T92q<PkV]kRH3c0iGo=E08;pn1;C5QplBJB0VUgMGV9E_GjU
5jF=dXP4Yl`3FU8qR]aJViZqGWF5cnp2n9o1m]RmhKHV\l5]RV3FJ;\W4BUh?2@L
PdBCC2k_;kUE\b2H_VUCVeTa_i>p^OfG?1[K9<85Wf^RaeXbG=af=Z5cmKK:?@dm
ERF6mISJSgT5?6NL2C33DNf[U[je^o1hB>=eE=OnJkZa]Ta2U5jhl\cP@NKFUl=M
KCqob\LWg8XY[m76>WVHGU73oO`HT6J:kbXmbN;n0FKb;?9aFlbk1Zkm@iRPf1Y`
5A=oOM4mnXDcaLAhh>T2Phn4Mlgdb3cZTbRRGCIKQqCCRiaa[BoVX3g[n_=?Cl7C
E8Qe7ET]mb<gF1oY[5iIU_@01dIWOod_Q:F4[jIR=:CA=FL;a5h]XRSd2IK>Vhd7
p7O4?_@AUGO[8JoI5<TE7a=8gPU9O23C=>05\;UA\F=UlXOEF^nGVN99@WR;5nVQ
U7<ha\7MeBTBm8m@8CUb7a_?ehlXPNnC3f>5iW<q2l9;Zg>W<8KiQ?MZQlJ:Rjd1
kX^LAKogRhS6fU166:\1=F0CO3I<1L_B8lB=@QW62IG3j=OCPo=S_a^d6FPO<J_l
0A4j4_o1Z>L@g6qlL^DAT[:Ohj1UXjIC41_^QUJ7hi>DWAm:Ki8@WR\7DpPk<^Ea
dDlkZPG`a]Z]mASB;E@QjB1<4lVUa8Pd<hZBN5BNPAOh>J`ATVERA\2TcGPh:MDb
]hXnNBO65TQR4DE4p_J5W\MpJoNOWnL$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR2HP(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
314RoSQd5DT^<^Va:c5gJNJBalcl6XIECD=_Kk=1B6X10GHN4U^3[EC=j^2;FX6M
WfNEmmTp6K4<\mEenQ=BSX48]mdF^9bAOZ=n^[eBDQ1]WU?hWWpPT=h?>Ca8E=ne
h@71\Pi0jTDUK8LHJBl64`:]=G8cK<o_4nm3b@Ff;Q8IR4Oh=`QqYYX49mq5i4<a
LQcTN>20ndnYA0I@QW@jW^IF8GYp^52CXUHplglfY?p8^?D9_OObAYYmMU5CL=\m
`ThhdD^n:Z7=Z6Z49MWgkBE?cbYH9Ng>KJG^J_;QcRL8_[[PKM?:A]<bGebR9odZ
Di@;O8:G4ZfUY7SWjp?HaokjBk]Q42iLF2W1=QLcabM7LkE@W`jbf[ALY1ok7bIi
\EXYGLe]8_lR43HDHa?V;VEXD8lPjYBUnS12lP@D]NG:FhOoWc0QAGPcp=WP=:ZF
UP]6aoak=4ene72XVHHgmaSCZ3F\R9S]Vj`Kj>Raj`>@KoHOXYeZ7\6fZ=Uk`B93
:4XomJ8N^G;j_bJq>ZHHUj8nI73SLFQDV0K^1D2R1:m16f=fPe88k0Kfg5MAJHEi
9Y7T3Y>kh]bna^gT>4Nf??_ndfDZ5m^gEb3VfQif::F1gj=7hSmli1q7QZ;6=?ol
KDENNB=Wo;<C4TQS[]eERc>S:lhJ>_LWc<E_PX`iJV^Mnaf9ccSISAO79dWEnaAV
AO8>D3IcV9I_b64@9:nCHc>G\3c^Qq9nB;:0?\SY^C6g4bXHm0[0eW7XBGWWC3P9
U?K@@eY\kMi0ECqU@RiB4fV3_HTdW3hmn[DBf=QiihXdhDcR<<ho:f3Oj8GnBTSW
7X9=NRncK2dbIJLUDfkmYL^KaDHVk]>435RNRqPe?V\MpKReS0n@$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR2HS(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
5<EhASQV5DT^<E3]L^OdYLeLqHo1EIo2WO`Q1aS>\oGAWNnUF:0jaS1fT[=b4C^_
6kG7=9WX7pj;GfARdjSiJiC[m?:6PK>I1:THLe`EOK4I\=Klbp5f;B60q:klT24>
G8XJI7AeKoKNLgCDgB<l\E[gcqHNkWmHapHfnJaDpmFhTK23hQc^CTh8b^Fnb7^p
UadGohZb?6]E15o<jm:a4L`H`H_>_`ZRSnib9>BU?2AU557kNB[B6Y^HV_m619_l
U8:GOB1]Pm7^On^?nBT7S4g`Ej=mGMZEe_SFMWq1\o_Zc@QN@oSo158KQg<E4`T4
Se?2R[U8;a?[MW>nAGmQP3<J?IAI1<YOoD4AGaP1^IF45X;`6Ckac6R?bc3Mban2
I06j@[f6VA<JDq4LHCRlj0JXJ=A1dZiQ5B[Kf1:4j=R^0K1ATHR6\lG8NVeRndTT
\>3JLTkc4i9_NW4OF;lZK^bHcc5c18KGDob9pE=Fo70E<`TRnn^BdZ3GI5_LBkBc
nOBnSoA1?dg[;HE<WOOmogSOe11Ne4eTLR5JAE6MGge^]\FEcJPlDoXiYUOl6g:^
973nSkBebjXpBcC6^MNcW>GK=j5XUDUMmI_oPV6_55WGGMDk`PgRA<If\hR;VVf;
VYGUU<7T?hLOB1EmBj>FMVTRJCDBF5U3SMYQ33YTcHWZE2;0@Sp8QOLVWjH6N8:L
]:6D8l@=KgIM;PnaQl52h?7EQ]>^G8i=J1C4=he9fRj8GdKDCTo8397XMT2M\TKN
657?e_VU6pl2OUa2piK<Ja1TlGMYHmT2]ca>II]:?L@1<9Z6]`dHoU]<6iI=40G4
40c4mo_X_aHAq?nQFfd3$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR2HT(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
lY6@iSQ:5DT^<?2:lISX_ADeclXBNVje3FQ1GPpGMeK;=GWR]Lj7m7><8Ok>\[TA
a:chP<4OZjh7;PTWmSk3>Eo7P]:YOSpM5W3jXF2T<]IYWWCpkfblNcpL3o@GM\`?
gb=1;MU<Z]lViG2W0>]PN;OpWo8QNgYq\KD\i`pUXWVQ_O]:e:?hoVY9HSgS^li<
=AE1;WogF9:3CZI1?Q5k>WR=8GT][Bi?4oCQhG6U<ZOBUG^fW@`@9?SC:n<<4^iW
P`[Y;Wa_W_loWpdQQaZJHRTBPWlVV]=4?`MP[4R6bf9HmX]^4c0>RHRM=8676oc9
ZP>mgg8GP:B:b]dBLa[llDh6\N^>:AV5_1j<:i`kPc6Umkeb63A<qH=W]:@0VWE;
8``HNRgl<k>hh`Q^TGERbi=dA3;p6jb]:<HQ<c?D@IPSUC6KWITQ_KL`EWjhN:<A
5DYhSMZ;m6d]NW[8KBXB<ga49]bk6\dP4nHCX>T9`jF?]XgGj^peZdDllGaj@;M9
;^\:49AIo]fTF[iooV9\Mb0EZkYj\JlHZ]RN?<eQbRS\6el\`0iel?6O7DCAM\g\
Hf@>QHdChUVPFL84;VhE1XIQ:qDNM^jKBE69[2;nTeO3\:@E?lSgc48D1f<[YFXc
O5m^3P5o6`ZHfbWYUm04@Y=n1=Da`Pd7LiPNc]59=B:?PXga]nA`b7en17okJi_K
qOn2=CX^FCJ`GKkb0he4>iRi=ekBI?WoO1lL_a]KfW2XeNMH[Q]^XT3:g?BETXoL
2OUhP3<TL>S=XdcIY^TMHK2plU14X5piACij<Xck;hGFSnCQK@gnCTJi<P8Xo6H@
A=W2fe^JXfVd\=UI@:IL6`3XhG<92b`\?HCq3eD4[aT$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
FSO6;SQ:5DT^<K5a[gMN`T]OGYkR0a]6><I7K=55T3BS>YV;ikMpL5eh9D3gAeE9
_BMMJ8XOB5b2`LY<T17oDY8CNNhb[:U;YIcdWTaJUWPdO=@iPhiqmA4g5c[9c4cO
6WWUFboV0CihQjgqg?Y_bDqMD`\<WPEX`JO?T0=`dS<CMFJ@A2WM1loR8AbI3oqR
5Hii_TqZ=`nfGpA2aCOGec=5VE]STH=Q9G_ka]8b1=N7R[PKQW@E:iSY7mCSA]DT
9Lg2<R[C^Sa3ZAADjAE_ZaF5OiA\Xe6[gh@4=DoQ`g0gi2CKTWRX4MBE@VlIO9;@
1?hjp5YjBjS?TceDFYLCQKP178RVa>1Dd;bC4W4;0O^F32NUdfZnOV;cP=Cq3I>]
^E9OLY0W5[8n3iN<caA^<7[Qh:@2cV0=CS0GW>TXXR_LX<RGHe77Do[8U37c3]Yb
\Df0TiV:LQaR4f<\g0n85YjNRc?I\V_V9Th5ROL14I=?@Uh392q\@@ZYH?=PdZ`6
Q7K5Z\3D5S:@C49U4Xg@kdb;RF425dEF7`AI16Xh1jWoH30]g;=\oDa]UVeYYc5I
1A;^H300j?G4o3R`0]81kRi[fIVZ51IdJFB7Pl;6<q5cKLT9J3L_5]i8UDMYJ989
h5nWNK`WgVdL7;U:Wea:791O5c_TLJGkkhahMTk3=c5B9hX?P@=U_iH7;:AHScP8
=ge2KE^d>JnLZN>j1NLoUI>3Dh[\NFjBqH6E<iH\k8hd_>R5J\I=kTlf_oaCAHm=
@IQXYVh2Xc`n77Tc<`C^d`kBO8XnP]dk1HJ2M;4\ao9BUWE7Xg2N=WYp^h^YH9`;
dQjiMFVoE>QJF@Nd=UG>J3H32CFa1@T:df=8P8aCc9INFJUVkTWSU9ohh`:S^3_e
Va3WkiAKR4T]O]meaH^^9=INT02[3BLi7l0^nmFTX3U5\Xm2=@p_fnJCSR027lZe
j>V:mo[@\KhU9N^]WoC8@82jg6a46cJmAU3mfbVEVVUJbW^]Ae8eA[SnN\YZKdbg
o]no6CagT4=O0m`0nS1>XZiSga\C:LG@kZmU\9S00M7oQq63cH94XOJ`34C_g?=i
@]8m^YKn<:eAfU9jT:B_Uc5F;\KJVUP]^fT=PPcICR\Hc``8DcbiP6=G4`lg[S7g
::Nen0[6UXM<M_GEc=S_W9gCbdUgZ>:XPI>BZo8?qjRN8c91QU;VakFZTB]SFIA`
\@;;mn720`RUTY7D0==KgLUEf]WYYfO42Caid8:FCbS8m3ll?17T2eHRbAAF5;Jc
h<dfQ>b`ZF?k7OX;bDoXZJi=eiSKhH2J=d_pKJcOLPC8CG3XDP]Pb]2]A2BCQf=C
M652:RYD5nX`7^W8P7c;`n=YVD_l@g9d;JUVi8ng`Fd]GEef9Zi7f\8EG[3MMSq>
J@bGC9`ihG=6G2PNj5I<Wk>0g<bo;Y?dQOD^n6F@QcnHZE2:HeeGJabQU[`772P8
Xjp?LFC7\@BJ1^f>49P=2IJHm]FXi0_HK7?OQob3jg8[neM0QD8lTGW]nZR\F<I@
<ah4OQQC7T:3LjRO1NGcmi?VK:1IiidLAdEDJa8SiGQW;b\J^;HfQ7kF54oXf5?Q
7qOocjkFX\j<KOY3`4[CniMo?jRo0?B<^IF_\^chUW_=d^5UY>l;mZeXW9UFW\M@
0j4[_^DQG>FT;MSl?<R34CJaTGMh`ROf@ZM5Z78h>VM8jYXX<dFV33eVD2H?p>m0
ddI>QDKPJnBo8P_0N<IagaQlOdTKQc0goKL`PJMJ?fVK:8QDJAAl7;KngYcS[i?m
nofV<[\c\fGI8g_QANUA;?QZ`7LMEWXdhf>WZW[JOl\^g`cRN4i\Ega@PIGpOn3`
cI9>UZoJL^OnkAFAQL<K>9DQkiPq45NLlmB_]f;SMfBW=nV^GOX[0=K6b9BR[0bF
g3_N@nbKDk08SY\2B0S:EC71VE`jF6Qie0Pk\]@\jkML`7LcWUQ^4=h6HfJi22=n
\43Fo]d3:GUn@I?NY3l>=dR>CAq9^SBiibU264SDIGB_JF>:M9ing6VacD1b1fk=
kIT\@4j4?cYddh<CJak`DITP5f732<UXICG7_d\1Lh8oTHBoFk0B5E`11p[DHN[4
p[:SLdQUCTYHBITaLVFT4qL20_@ek$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR3P(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
k[WD^SQH5DT^<H<X5QfPgYb:[XjF6[dV2cPJdI;gA^KJodN__5oIT?iHRbMB77EG
q6[I8TfC63Uj@l_:<XLnYN5jdGf2RQ`el<o]_h:1bokiZB5bkEnoNccSRoE>gGN;
;md^Go0f9p77N[DULEnC7Y\A?encj;d2EYT[ceq[:S^amq]R4TY:\<?kYD?K4VMl
6UId7;]P]3hKm>\n\_c62p9Ga5\FKqE7oHn03H]_CcL?mL\`U_29VN6d::]j\DBV
_Nb1[4UE_3IAi54[HeGbq>3oABXq2fJQ1kS\lm8fP:^GgmfDoP@b`0@BYcmD[7:V
9d3A8H3f3MbHMm:[cb6T3`1ER>P2_Q\6kQ8F<URaOURnP8h38RS:LoPRXEHX>Z7k
AdfieWWEKh8GgYNe`n`2jWqZ:?CW`5]nHPQ6F;WG>D[T2E9gS5;c@<LU9o[gem9:
\]SSj7lJ7K]b]:<P@=[mI9[EhCe[k\ChlQZOlhD4F]=X<8kLGknD\C5G@:l\H2Pb
Mm3_nV\jDkk[3:CJmp9VbT>4D6oSSTO2dbT@9H]:6eG=c?E^HAiS^^57F4^don65
Y]KZm8PUXBhNCJ<B?ShGRV3B5<DYdg`5LKU[oEMA?;]5Q>R9DJb`W\UCFGi;HHac
hY[QP29eVE=hpCe16D21o`Ud`k3ON;_menma@<<FM^Tc?AAgaiZWPVonNfnEkZ]R
JiDDi>L6Q1XbhGW7\j87WL1cWjY]9IPQWQ9mUEWjRj0K\YXmocZ7T37L@SBD7b\N
_3UiL_Kql5g7>j:L8bW4_e<DEo6NmDUY7RZI0La:81]MMf3JlKhaI`J0OZDoJSJT
QfnBTSQ4H6g5ZV`GUO;V5XW<Wafn2EZ]GaqeiSCT\Mk4IfSWB@[5>RC0Gj>NSYN6
NFCV2GDP<PJOm9`6AA7DD<YI_;MWcG[af9oRQl]:Hf^:3FH44]4OSRY\IP8ESYNN
I5ENh6b7^H^SA0[<[XQ3kKcFRa@`@N0V4p`WJFVGW@b25cmUNn?`;AMQOeW3RALA
]OjXnJd?7d2W3cT17<_2RA=Fe:R=lNIC512IVHm0iHnij;b0BN5TdC1U8gl1ZgNc
BO5fQR;?lc7@jL0jZ4_8oo`PTQb7pJWA_OkngS3mU;d@YfGETc;N^L732EL^016N
<PEkDgAVcL4O=m07VZAMOPA;?WRaFcNC9eGC:Hgo[bUChb6O7mm81a7A;_hSIOi7
Uk7B1gSVLL63G:WNP\J4ZL7H0SmqoGQnGUkH]aNQaKY5E?20R3^TA8VDfLk72nEL
GTODB061^QBI4_gdaJ5mfCmk<jA\N70cC2pVGPbMKoSoV4J`gKj7RW=K[fA=SE1X
33Vn==HSPE]@mdn2:o^1kISKa?MFQAZ?60ZoBA[40FSj[UK0S=h5RYbH8;S`S8li
2iOBQ6Q]8:\hRKNk@gln`;@OoQd_WnGn1qY;_RFgReoe>o5iW9bPni<\nAAn8G8B
;=1V5_dOeH@QELk]aGJeiWOFH3[eFj?ce=P2CNgPE7PB:eYRRPPPZSa;3mKQNGOh
qDe396D[eGagHb]\D?<fi9iD[TTL2PKQSmZM;OHm?jn3Ef\8EaMA1eVnHfh^Gj4O
GMGGYaP\NW[nk4Fg9XKlRk5Bo;T5eC1Y7R9BLcfD4jhP8f=UFXm3\nCXXRG`FFDq
a\8bAkU_?O\UUd9jD1PXec[McMYm5]V2mWL8XTl5:l9H57XA=ZjVcjL>\MSC0?SV
?n<gSP28S8APb3KUhle1M_D;8MYkPNkSF74RQ8Y9^M9DKcL911a:EMRQ]ITC3opC
]mAajF<cfT:BUG9[XD6=@Th8do44j5ZeNKU3hg;m3oT\Sf0\AKb692jB<@hEa1nc
jij@NfShNFPdHWSmKh<MSHZfdBAG]mXHl9kl19^T]5=AcT8NhFNdK31:H2[`Zpfl
j:I;P1XMOdag]niX:TUYV368lNc0<Ic>Ja<\D1AT4M?>kMgVVKpn`l9D8R05N=0n
QP0la:W4JXXN6B_RglTI5@8\[XbMQaRf?@4BQmLZUNmADcmP@YI<R3Y=]6Z21bd<
VBKQ@IVP]dYo64?Mkac1l^UJ[4A9Li[7ocS?MjPjBK6deGJ6Jpn9b@io2BC@h?_m
kQA3gV\MS=FQH9YED<eOk4Q5dbGg?ODO_fGAmI]5kIje>E?KSY5J7lYHZBhR[aU<
=aW[A[C=^0;ino37pJ4iD7XpN^Dool>$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR3S(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
2UmB5SQ:5DT^<TdMc`9K3^i8YWW0;E5375el?0AC<]j2nc?n=jmlZN8=X[CSUCY6
98VB<4FgB;\k7n8q<:0lRdIh5@n>nJWqR2CmhCFoNgKbNf@LX4ilD6<pWlBJ4Op\
P>K^M:XCDLgJaki<0J^P\a0@TP:cQV9__XKG13pUOGd8Depc:0=fGqm5J^O5PQi`
7MLce>MO:Pnb2goIDkQ8hCKKAd;@o?[@X=dffa7I<EaBlNUFiIlNoNmfkL@;2OUi
\jcAUAiW^>OS5bm\NC8^mTjKPhX6`[NQ;FP<U@STCG21p4oG_7\gTRC2DI0:aA6Y
P1Z?GkA2@mAL<;3S1mEhXGi:f1a7i\KePT\P\dQkYjWO`UdWV8Zh3pQK9OVb]gcT
6n]_8;lEB^;[OiJl3Z]^IS^Zfl5Oa]D=f]o<;1Da^jo[bZlHEH\MUhQJ1mK12I2g
h3kWFh[T\\Dd_YddkNP]B@?ZJFESgLdNY=aA>YKi:C?`qk[AI;\nlQ_XOZUT^BiL
:o>fIhXh8FgLd167U]>K_\Q=LjmB_ZcIdAGeXC;^8L;[BkG4Hfe^_XEM[WWV58X0
AeJNLSNcH]H@\^6PcjAFHZHT@Lj@e7l1X=2pR3[9l@YHDNZde0SS_fn78N>L3BI[
P7iTY_h[jIi1eAhH?=^RG47V8cX;=]B4LJ`PRVa]FV1n@neVIb38PE7WkC5eIY_4
2D:>?_jFZ6\[BEaRoYBBB]92QXpXZh8EoUPCSRQZ5[T39]gXC@QA2Wf[8X7FhDg0
8Xac;H^mS0GZC:Cfm]X=JUGdklBXn80K[437CeVBjdVKFNTDYq:\4aW4e@Y`NXJh
W80?\EkLL;:H0_L3PnfZgaFNMKbA2NiRF7j:oUe[WP[9594\K0Y]aLI;Q6V04<1m
f>IXGMJ9BelkVLhbI6@GkFKT[F?icm`M9iOg4gI12KQ>qO@ck4\[=Re[24mkSg<F
LDEMFaRb4@e]8jF[E@Oa:Dj:4cG20Rj>:nk82SnnDm1hWbQNJhc1BTkI;8YbaFX4
G3YSFjg3BnmE5VLcD`Oo<h9H=k]<d[[g;UV0`>nqL_PXPUUW:N[G2oah7KR4@R8W
mP6e<?nDd?JdDTVb`Q@LKejC;eDT:Qn21>BhR]SO>?1LgQZF`3`^>aoUi?@dD=_b
nfXURKeFj9cZ;T5cO9dS4HAfLl`RNggmAIqBZ88<j]8PikRQ:f4hF;G<lbKL:1SE
E85[Jq`iUoU1bAW_QE^gMUDPe9@GQK?AkaZJ6?c46kYbeELg0=i2`8KCac0PEhFY
Z@2Wa3b9mS\U[J^E1U4Mle]gBQ<U5INV<19I<gl1=m9?Z=E^;Dl2PRQ:FMh;fm^]
p3G^B3Bc1@o:Sjf4^bcFaSK3ZReEmfh<0ah9fof5:JT5Vim5b>0SbMHA27<A1h=9
7U55bb]M<k8L<l757QW9J9AW?oKqJeY]k7XXZN[8Fd:^<Y>:OV`8b6SZ;I78L_EL
hSTM@32AIdXU700?JGKRlMm?TVH6g^@4P4Khj1o@0\357kG?A8aU@6W[Y7b<fUiQ
9Z:aYY<B=F@3^1<l4fmJB5gZkKp7nk4Fj7mlIZ>`AIhEB8iEaFKfeTS0cF36nA<c
?8FHon[4g@QLKeDdNWW_8liSg2fPRS1Z3IW]S8KiTaeZlIjanY0=eSPcMYS8<>mQ
a8QAVQ0GXcK?KdEEX7S\[H_HSp:bcmncncn=i=7Z2aA=2QdZZ42gBh5K;Ubbg[bC
4UEHF1Sk9K`YN3=7l9M?RW`>UYj?P@CI6BIK7:<[6SHDSJQ[Bm@ggW6HELU<^351
dFV1IlKADA9K03ECMCamJQZ?pXMo;g`3VJ8QHO_La70lX3a[0k1R^[g7>;hRPoI?
do:emIG2\20eHW:<a7C1hAVg41SS]QBX]b_=:[HhP1Q`X8alBE1a9LSU4[fAf798
?^4T1Ph:M4dBh3SVCnJj3]7pLY7;fk48M:EHV`^DbQLm`=]6I=;X1ocSn85O^YPB
CQYGn1=[loaHZh^Iib3]eVJVY4TblH;ZG[iejCHOS4c4IZdCT_k6`Eq3h1<?cp7\
I=VKl$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR3T(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
k\4o1SQd5DT^<Fg]4;QQA2JJ>UlQR3=9qGgOZ_kS]Q6C0>XhVbhFgD]V<W[MFEm[
U\2q6Tj704GO<b>kY\egBdj9^=KqL:go4MqK>7m2N\b<X\D_H9g:;amA6[0H]k3N
7AY9[\98oYpFLB^kQWp=Jh;dA5Hgh\IMEkJoM_S79?K1EbCMO:MAcNNoHdcD<=fZ
=pUIc7``qo^lIWJ=BDVBB:;c66nGM7m>\W33XTMTPnnAQ8;KA>_EN`PBW9Jmd7BU
99QW]:1KgXU8o98VOm7Dd<f8Z\@TDmcGKf3R7HJTZ\C@b>N_og]ENH]LMQAQR>N4
6nB>kbmqAdd93dR0`GbCM>HN1Z3mJ2P:F5DEV3UH\AZLHMC1O;boYF=W6DC25HEo
3Lc;>dIGhYcLX7i??D^6CBkhhahlXIncg5<PFhB4`5^>066AM_gCi\nEmZTe^Y=D
jRh0Y[qFRND]mgI\1F>neSiCA7^OV2=]Q^2W0LOo=JP8LgeVj3Ah?@cGbIUWOAKa
iX@F_RD9fCc4OX1iZIELFCHm3WQ7Pj>LQZl_gY<@fYJdNW@[[n0RSeh38kmBH<SC
Z=nE2q1cf2V@b@fEjEa6EHi>VPe0jb;T3OEAinY1TQYXb9Z;UVc82NU>Y\6>X1V1
PoYWmSai?5m@=LX>F0bSQVWhO^Yg]VQTU4OkBOKH;^[Lae86c`FO9RioaUFB\G`B
83e9q2C__i^=Ij_fR^W7fkM]0mDec6E`@:<fLAW5lf>`OIcnGOTW=e_f@29mCLTg
HYDA]EmLJ7X<S?L2n8E_gFS8>8dUGIGK8Vopf5IoW^Wb:?=MFZSJec\X1jC=hn=Z
LG3QR0@B?IeZdkLHkj5c8LS@^7i]jcCZ62LJ[^<lcd@dK_\d;dl52<kNPF=ginYX
538[Q019[NY;@c7XLcN2:L`@?2>;R<?blYqbJBdk\8cPb5WgI_6?E7PV<Gc[LmYD
]LCYL6MU0cdK?MEb]=fIM36e<GeogAE3>3:Wj?<SgE@Qi0RkXPkhgl0V:n2MLmJl
0o9Ci1GlXN5JHRbFJiFeLnHCEUk=`WmhlqYCJ<c>a7R[T2_mad2AYOj7@Xh6]jeh
k88>5K^9<1GaB\m`in6gVD>gJ=RQaj@dM2=e@aRW9:8CciP?gSWo099Z\2M6QgmX
ZU[3dFW2W`K=E9h9Inkg:VJD?VToW5k^p?7=AA30dX=]86eVnj3@S0b9OGKhT@j[
E2@N;`8DF@L`FOQHC1iIVLQJ=H2Wgpdb;jMn1_Z[HUVJ?f6cQZ4eTN\EmQLf3k?K
<>S5P;TR>HRl2<jUAA[\MU7lZbXWO`SkTi;Ll8<[36RA>>Y4[34Of=^EaZ^T2TFk
K>BCDkV[TI=34CUUaA4KSQjDHX2Cq_M5L9d?3EV51aHY8>^leKBMf^55NLkTRCT<
BNVbXYPJ[9:\YhU9ok9m5EFfM@\Cd6PcheUL12`_Fg653l]VoV>CFYQJbj\p5BmR
JOFhg;hBlk\oU5j3cUH[KgFeS:QnZHFZ<DGRmP:>6G?hO>iljhnAikJa\P[h9ZF@
nD2bbP:QC^0EG6WOKNhW9g0@0ZS;`SRN14N?h=RJ\\>UP<WC;YhC7]5R`kp7<T_H
IiJkcM2D0\RhAC6hH5Y[g<\IS\h4gd3P9XDPEEL^id[4=Zn>G6L[31RSWR:\^PJb
j0L8;[>VCZ:f>`ECo6nng1jcRj9]=I=ljB@;k1HK`7DAJUT5ih6\VbGKGqgh;LZ@
C19fU>7M6K?DT;cJd:X0[eW_UU1i`=8@W>BL^;c_3X;ihbME?X62VGHk9^Bl:0UA
oDDg5]W8NT_1a0W?kIB0[7_\Z:ScDoQM0>Dk=42jXAjjKNQn=6`2nJ_4q56nejhh
obZE0dai5jI?cfY@G?nZQl_?J9lM3Yhd=;GlMi09ggWfQ59dEeU0EGilqIA>RgEQ
W[gk;@Q4XX`:N3`SDScUgkO]\MeV4SD^GW:JJ07TeKhLmSIo[SY7mIWAl[bRTXP>
B4fE553i4AcR5E\cQTcMdFYjoX\fE84KVo0eVGgEPClic<MORA6?e3hqGmDWLQi]
G9=QaG`4JEIJ@NSE6D[bRPNZ8[fjC>KA<LN?be>b3Skm2gooDFQ\\RmA]8kRBS:9
X[6o;ZHd[7FINPHYlei8oiqCi0@EcqX51]Ya0$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR4(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
PH`S2SQV5DT^<YZDEgJ>52>8J6JbiTn_ICV9ZC\^TS9T5Ipl7?@lL4l\aR_>8TJB
X1jjaOQ]c6L8DR]HAeG[eVRnX@mER?a52]L951n9YWTbApbUbN>XBobWAZ]2UW[;
cWOL=>N7_aCj_P9\FLe1\qP2I6b?q?3?4k2B6VQ44?D2C]7iP4c_ULFCLW[fICBm
kXNAYIWCg1^pTke8TbNp<>SZIOqB^if3o@gT2V8B7a5M]<>@c9N<HN^4oNllLfZp
d]bdRmf?PX2`Y0hDQe\Jb5<eVNj<b\ET2\SgI0IMYaG@<IPE];S]ELGZmYIYQae5
i3C?abOV^km]4`SWl4K3Lj;EeN^6>HdKMCMaWkZ;>PJ3C9Y[W?4haD\U>[CP:Ra;
d3cAS7caEE[APWq1ji45CjTb@cN=OSY3S_BIKT9889>P0I2Qg?_eAMLR==3fR9R[
:hJa7dXLmnieY0]6iS1;B[YHE7YKGA`V04B4>cbj8W[;kYT1NNA\8^5l<nh4h?;T
3ZHXHXB4J3SGB`K1iPm?YV@R31_USp0Z^;=3geHL`31=DBFb?C2YBieiNkF`SYFE
FP8K1H`5K@kcV4m;lHm\joZK26fMg\E6_;;A<5Nkg37CUXa:k^jGgPfihk<Rml^B
E\J[A<1gVMhKPj85W_aTe`XPl;5Kc^06Y9V0?94T?@R`q2<Q8hRZV^ILD70TjnDL
o:S5b\RqEH<Re?@NQ164bdMHKEI=fheKF1F[LJHh==39O_TH:WVIG7Y=TemcGkeJ
kUYK2c@FGbnImF:cnN>Q_J6SL7@EAX_lg1F[_VE5Xj^JTS4XHnXD8HObdeED5VYE
fZG`9Wd8EbXfAXI5EM>d`>qJJ@EYdUSe51^lE\=kWmJYkeg]DYH6?6Zi=JHh730O
HJC8_e``N7`d^aOaY`T0j8MMQ>;b:SS81XF6QnS1``JSNG9JDYa8`L6NKbmd]og6
RZoJ5>94k\_e_nRJh`ZKY5RJQfbZ?HUL2<][7pch?3VYNEm=@=7MlafQEc84dGbm
n8?1\fJ`cfe?=fJe^NiGfOa>FOf2lZ@>3CL?ZhT3B872e8E7dcaT9S6nnW7XW;Qm
RnDcW`=?8EcmAlU^ZQF>^Tn3Gg6kT``jC>d]KEc3NCmIC[1NS9=DqccE_TL`\FYV
]dKTRnVXORWCAg77QM\LbD2PP:R[lMIbEe6FUBh`SJg^^6YC7c@OKn0Uhkh_j;d[
>EKo9POV=>hFe37f6kE^6[4;K[GSa^NTdNIA`YgIob1hZY80jXlHBc08`V5i:0gc
>\IqK_<_i4hb^O]H2]LoaP@VeK6<nd1W?Y<o_na0IE5Jmh=LO]m^\ML3l3bIVBc^
?KfGPKC^d5BE]?`]d9f^?4L`5HUl@dHUC\4=^kB\I5PQ?dM0kCP>^?i4AWYnGKbO
FXC\KKa:CMJmNb4DlWpm[?6Q>Pi^4jf`T>gD4A2F4@<1I@WG\1bKb:I7U7CmP3E6
WUR=aB33@V^ho]8NlP=5<OSnmdIh@9e295j4TbKgODh9[ADF7pH0CFifX[17DWiF
Ed3S^h7J3k9VHW>5PCl0^g26BZ_gi;G>FQI5<F>P@Oj;3PP:XW7Da]\TC`7\133k
I>m6PgCQ:CSV;P>HZ6hWT=<eEPHfiC:3^WQ1>INlR^Qil_:A>>HofOmEd1c?VTTC
q1KAI_KHS[c]MR`Pn3:lQ88agAG2AHQ9V9C\baW_WXC34[LXCn^a3ch7MP3KX96@
KXDObTZfJQ_gd5jQ9SO1Z0G=2aGeA4aBkA9X_4CHnbSLY0cScoPeO]l4Sm92AH01
G1DYO^1AR=Om^lXq;OF_h25?EDBk5>TKA`RjTOm;[<4k78[h9fjdbc4<\2_@U0`A
DRmqM9Se^VXSIF;BB5d3k=:eA0j:50N8Gl[OVo6?4U:1JlBEUMBJ`AcTM>Z739Zb
d`DDdA:fN=8o0TSCY5KGJ=gkaPI:L0[P<GKJXS4\]h@CJD>0?EP`Xmm@>59ZI7Cl
O`C_MA4L0E3=GU8N<npLI1o61J:28I]Bii1]3ZHlGR0`[HOC=_7YDQ\j7aG7DWB7
P=;P5C>1DJYW]L]0F0gB_9N0\H>3?:gm[SfZ=ELWg^B>[<1UmhjH00g[U20hHX84
1NW55`0Elk@b0IM4fj]L_n=IfbNnVc985p8Q\_gEI;S9_fg^J?]Y5bh1gQ[P3o^M
nDESJ`41LA\RLW^P@[KQ>mUQ\16I7fI`<QZ@kgYXWZRmFcYdF`jgFQ?fbMaPNBkY
AYVX=ck=A;<3DBjhP\jb;T9_<jC\Wme<OE8@2G]TF@UVBkOgpBeEI<P6:5f;\I\D
FNh57NXdGaBKHA06`cg5R8h\LEW]6NaT:f;4K0W=k57XS\@iE53M4G]V__A3=oCE
anA8lh7VO:BS<K:g9EfOWol;N6:iBl^o4A8jPF8AIOPWY9DA7B33mdKeB@cbA3Ip
MLDX<7@_XAYf1?8mJdo4\:a6jAQ5ZLU1\o]oS1jNcCZ@=fjLN8piiBH7@:\\02O\
A32GXVcA]MAF51aKjo4?D^L]TlU_@>_KdDCaY6gLbUo@g]c[_[2=^ZM5GT7:59XW
OK<`<\PS19155[iUhj_dhKTG\d`n]a5oNl2<gG:Y;SEW?5HKEM@ijT8e2bHT];`S
KpS68Z?SA_c5JLV7m6l66mObW0f]c7994P8eG`Oo<<QSj@\;n0h@N]9RSX[AlT@e
:X7X=Z^mBS>JgVeh3SFTh7]S\f8]4MLiK;]3E;4`IRU54NJcG`Q@BT3;m\F9^jNN
;GSX7U:G8XB[7SnRp?`<V=[RUo75_j@mQU>l=`HRi5VIoAcNCi=b<8=VoH`FYm:A
8Wh[mkM\YnEAmBX]cdEFMNb80XB;I4P<1kii<?Q\IZg5LfDqfF;nJR_bg0D>@MHj
VE7boRQ8@;3af8Sm0OIKOE5h3jcmZ=dFfn5<PFaHEfRL6T4fTHdch^E:?N:\lSYc
;2SMPWEfni7Q15CWmDnm3Eo<2Lj7[aPZT^c2GJd`0n7G@V74>\bj>0>[?mqO?YfI
_V^bJM9AFibPTCoKS6IXZLd`cW\_ZD@DC]goi[afZF;aobYL:C50<U0YOBVR5S`n
][SOH\@O0UYe_a^4R?4kZ\FVK<@C6MbAUjEVnke>P1\TDc<nRB7:=16U<IGO5SJ;
Vj?Y^FMRWqcKhlKNZ7\8jJhB;gib5RP4LFFjGg\fW\<<l;^O[2mJml9CF:GGZI?G
PR9>lM0AoQl[kM>b<4`2hAHIFW>X4PY8G;WjXE[[GN[JCZG:;oJARf[IeJB\Sm8E
M60XEaW1KTc[N:OcFjX1R?h6q\aE2K5b]e08<IeAA_KZaTf\e\38EAV=TYl_ISHB
clnaKbfl^\=dM0[=`0Nc9n02@^X6EYF6?3n[3dHcMgB132Oda]3`_YN;03OP[Ca8
[H>Ci;Qo_d\;h<2Xe4]i:;;[X\XXjf1\jE?^dgoq2<m]Om<YEeEmYJHQ4\liMHM:
5=7FMc7:cLVO@50_Cf>;T8QTFj016Pe\PXVih6]iOn=ACnQBKLXMb3n_Y`2:^gka
K=[m;]hnUWfnl`mOFT]ho6oi7V3a:<inBBM_WM__2n6fQ^0[@]fn8bpUZmSeX4FO
7\i[_RUW=9WX3T=igE>5[2B;@3n6FZ]n2gM\3K]bCTAWY8B@UD;\=:IH07oRCVG9
mA<3Bd@jCnG\6@;WgFVl4KF?o<amA[4eO`SoFDCDkZC^XY3cZ;8loeoU0Cjn85oZ
9AEUCqfj=aUE<BC]\Y`1^CoccLp0W7bL\K03LSg@>A_>cFdCeg4X99CMLh?<fof4
G9nJHm6\dPBYmM\N_DkSHDO?c=E9X\\A7LDThXT3obIZ<gW;=2hd9jKFh:m4`>Ml
2Z:7iBJDQ37DSjGgelJ32_`@Zgm0Xde5n_Z7H`lf7pj0P1M>Fg<27K3k_W3k@lTT
DPiCOeIGOk`AGZnS`UY\iIW^;4m8?c;F0^Q0X]7a7L@Eh91b@aj6jd9<QJ:R>=G6
8SlHUaNhZHf73OES3lF1MQ;K8B9_YC2VgG6M_nR`TR8elKC?8oX9qj3D3M38TMF<
iKPiEeGdI??h^=XCN8G]k34o1PX5_=m\BhcTJ0_0T4om<gno8UQ_DMD:6nDf_L5`
]Bk5JbQjQ^KGlYaq71^2R6SS^=L;=2Q6BhlgAiIkPkJjnd?k07JJg1\GY@`<g<AN
k\3LXSb6IY^6BC4lG2DAWO9P18LT7D^cAhUgC[g63k87Boccif>:7Zd_^W`=Dj]:
5\IK?7BJV3MCL`1:7b4CbOTl6:M:Aiq;h<fnm^9=PS2dlUJImHhL:fgcVEf4Fmij
;\?3cYmGQXc3:U[:;X462;^bmI=_N>i9YUe:TfZY4fo0>9J6_JX9UI3IVEfIH>F4
7HkV@SkT@Vlk_foH_UJVj8JF@@@8R_];dBb44lF1QLNUQqI7[B5^D0B`W@LTe=<0
LiAe28mNZ1TC^YVSe6G`GJ?I6=Wk[b<iVaI?1YL6<<HeO8Em6hGBf5_ddFWXbf]n
8Ag5^d@NZ]nA\3Tf2eL\XIB0=6fR4>iim36SXof@Ml`ANCIb69N]1<c_7kB4pFOP
6aP[[gj6V6HMKacd=f\NK=T`le:^P43p;]=?<]PgWY2dKUb6So6W9O_;AX3Nm@M=
ITRiggI`1BJAgg@XVNb@aRo9Gb]@dHCfMhdlgLJ_@G`h0@H`^5kicWV:LX2H^^3[
omO5Y@U9?_cY@]c986DVl3[ON;2g9A]_;PCBY7`V;7\M?kpGFcjlJc<mZhRJN=`1
]WnaC5heFa53lCBeRXL475doDo=:KZhDA1a?XmnZUJDOOn1nVB8Rna\>b\1Kjc4E
05\YCn_3FGg0YMQa2c7?6TX?J5Q`4ASYiNUnFBNA83NKD=[G3AfoAi2ejW;hnq`C
]H_@?M8M<CIeZNlNNJK<0XkNl;?Z>_P4g3?^eHgS40^RkEF[DjSZ_QMS@GP^_m0V
haT<7`=LWOV>KLW140WZflEN7;[\EaJ8Wg^[YK[?O2`PZ;jVl=WR7^Jc9ME6I1`R
YTTT`5EZil:6pEE^?bTT46P;2`?Gh>JFjX9iFX:J;Cg^4O0OJPd;JTk1mJRoh3CO
XFFJ;:WgkD1?YkOfp]a`FbgR3?lRdh_ATeXTMcIPdZafI<eF<0kE?1V_D4?ma57m
YkT[T?eRX8OKV<GNOfIc5fm]GFZ<50C8T^3;f2Zo`3afI6gnDd^_mHZ\Q1b]d7j0
_n`?j1jmg3497IJP<]gk@j]^Fa=3nh1piP1IgAkJ0c70WF`9\G2Lnn?V?LG::RAW
giMOLIKY^ogg2]1^g]fk?M@cL]Fbe\fcN;8OH]ZXB<Zl52[CQGdmUJd_WL^[M[n@
fCH5Dl5F2ogNoTAO7]W:KJL?WlJAgW9hi\^g4IlFl3f2@Lq;FjmjI6Md\ao3DB<F
86@lcS04R=kh;@AL>79hXIkfWgSM?5i6kj85>`QcU1UK6K`T[Q9J<@A79aTS@hBD
8MS]T[ne8gT\ap;cY?c9ql^ol?^5$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR4P(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
66Hj7SQ:5DT^<g4iAAna`G6jCn<iLE14jZb^7NHM7i^?7RGUXmfaCZJ9ZampYNOD
B6STa6<`==T7pZD1MFn5g;3NYkXh2d1X^J6bZcJG:JoXQEOB11DMnYh\07NG;q5@
0e?6pAEN8>fO@T6YYg1OJX?B;_T=<7J7f_icPH:Ibf=4?Y16bWXp::n5MUipD[A6
:7pbgITY4Onm[EHZO>8h0n3BWh8hDD1o4^PK=OB^iPN?c24^j=ccIgXNg:NR1Y\k
hiSoL:I\VM?3d@44]RGG0X=9][JcDOaWH?jKHkaa]ZX4I3ZAlV:4UXiRn\T\U1oO
gZQbLm5GFkfQM^P9PpN6n\KDLd?]<2h?:4@cJa_V]OFDMpC8]X]nBE`GMh3l\LEj
2\8lWLF3>neo6jDYI;7=BnBIP8RE;LBdn=INC_g[POABHJ`DRHN?]ne8[<`iE3D8
EiBC4kf3>XPH1V7[cO0BoNHS9n=kS>Nae_725Pno@K:<T[CDM^T>KG41[3<Xp1`[
UfkWR@JcjjNcEoD`0J]bfR5U2KEJ;a5fQ8li>E?6VH7:WY<BF`HX7he5CI6g8;mM
@[]SolZZXXL9dkeRb;Y<2R5WgZHZ0Hnf3f_fBHB5DH3eQhI6QY0T=?SM:34fX1m<
:F@MbGUDe?lpFY40>nj>a;PoganYn?kka``D?NmAK`K]S@n;4cah>f1cWV0iX_IZ
_l9F3`AceW09Z3N_5Bjn[WCXZ7GfQ8L8NoLVjNM3AHgI]9bPNJ59K1TZVKhCG`b_
0d>5hj\VR3@\F35o]nKP^<TH=WqK;lcfo=gJ5XjFMTlXJEk6@`McfaVZ4d6BRfgH
6dU?>Z:BYd\_c?6]bF07PqLIOlVm1=W[K3?lO=mHafW;6Q`=GUmWgmB39B5co[Pm
fkIjPQ=JW=CBA0D]kKV;3B>_LG2cLH;cX5@`;UIZM=]@hUD=_VOI2?RD5KOFB[Uj
U3LcXRg6^4YT:@7>9W=fmHL_LAOjn9T[SUUQqV8eU@m_DCEM2:Z7=F8WlRGdbFA1
Km921;;Y\b1X@glHMLFK:lH@]FUKWkdI;Y@ega7iQL1BXnFFl3WnSKMW2PYCOXAD
Rc>1ATMDhVI@`5cPK;U7^g^Il9JITSHkR<VlNV733HT4LTCn3CGq2c5AOG8V]YK7
?NP>EYG5WRdXId5G6QDNnkXKeE`jBV6D0j;[TU]1A77B1XmHjenFYcNFS2gPhI_n
P\_=BXHHYa6mOdIc:7O0eo^E7GffS?h:H]7648Qh1C[Wn78Zg3m22cRE0>OZeoJi
RCqWH9McSdeEc\A7BM=bS?EDNJP56hn>VOm0PBI[<5o7T0EU?DeLdl`\jQe0]jOd
J6JNDD^11GY>]B568gA]SHDij8L^6>c;K`\UR=jmBGEnU7E`;@Xm[=JUi^igg;:l
4aTWDnX<Y?RNn>6P>pGM]^1a<;;^Ll<9WMLO>B?7US=2SMh>k7G2<47lDTF49Da@
:]0^H34PSG`bj1^Ecf76eKic:k\BVL8[9;@O^7fkS9U>FCR2qn6DX`:W_g^NZnRO
o8TMNm2c@^UZF>SdToK5iT1JHM_e;[kOMaeM\;_mOBQ\OA:L0ECPZY\@l\DLMbR^
D=`:J7eoWJU>:IN0lFTcDUkL:2i^DTo\O6QDleU@?]TJR?dUTn?b^Tb;oZ8ln]1p
K`FUW]AOUDkg14d2S22KdF6D9[8`]<RcZocEnKSDin367^AB_hAEV0?6BeQTKo=5
;gTI5kR\I^YO7^J6eBVT:;lW3[:[lYEh>fJ_4]JQGf3ohJOiU:A5X12VhVT7W@0k
KHDjKcP4`ckeV9q[3RRZ9:CO?I3c<5@WJ\bVMO\bda6an2C_aOfjYbNUO4QTjk?m
7oQ[L8RinjHRjlb<7K[MZ>Jk30[BK6YO\8EVe8EFda65`iedE\CKddd40cjcSV?3
Y=F<7b8T=SDZ:a9[WfSFQC8JjQA0=q0U^gdlCE>;12@ZH8_BUS=fWWlh8??BBef[
q0[61oRH7o?_?leoZZCO8SLGQEhRAV6?>4Pgj2U9MS;MkZcU9UnSCDnR5I\PD7]T
fDJmLKOQFMTJXVH@OQc?ZcRk\Dh[QLC`3?l>SD?D60FB1M5DN@nHCgDEKYjNO1b7
d0JUFo;^J29=6ARp:hO=ej15A7WAlHogl9M_4acADR\Y_?Qn^76[0oNgo6lo6dK<
fiBk>7k:lk3DLZ:Fo8FEI@bIVZ`4daPTOeINfGXh=RTI3kEGb0eB?dCJ0S8nfhCP
9fVlh0jXAcOFEl2d:T@Wffd2OF8_eHp4NYKi[mD5Kd4M`3JYdC]MJQ>Sb1h>9[Ug
1o:Y4\ojRME5:DI3Qb7;?GjZi:OK<;[\U?ZBW\?>CeU4BC>o78:CFAQ>b<7CU@7E
l0NJ1d?QFVlgcifShh:CeUU_P`6NGiF4U5>]aH:g7:mFXp1HQY@X?Ph8@\NJPTAe
gbmkA?hENOUcBQZa1\@2g^^^C5HYod^AYlmd[[9V?;F=5QbaDfnA72W0D?Pg2\l2
\bCP>KiE`:PEj_PaH7S3ZIjP]Th2`7beEJf]RA_T\3F3XT1mS=Nj>D5H3_7PpC73
d6D^66GJNnY3?42n5PP0_`6XLiXV46WdS\CJ[0cB=AjfZ97[U>NNd8TU0D7;TDi=
An:Y2]W:UkE0:P6dm_8:Bd6bMHJi4Z1^jC;46l3egD<;PfggjNb5>RN0U7nJhCT>
J`l:F;;JLLnq>;@PKoLZ;fH>hT`Qo\4V80?C7FeL[M6hjJo`i`n>liaU6aL7l[b1
R2J^3>XSak6kgC=_bUA\QhlFPS_B9:n?=V1ZjLHmThqL4FQKc@M8\`VFkH?Fa93D
bGD3U;j3fVe_hio^]Tl9e7RZ3ok]9Ya6cbJQR25nQ;Q8FbBMH3ioUiQ<U@VD50W4
1a;7UU8=8_3K1JZn1TgFj\J[K15OH`aYTfGN4`0[=??LFkIGdVlWXGg^5p;M:?Wl
TJd4M=SCdgB0U]2Nm4f1N4k?Tj9\bYN[P9CK@g8LSMgK>aB]6JS>[I2;T]MRC]DE
:_28nb]bOFoWlCMGNc;1I4i=E4oCBXKno>4JXb26FlbMa3:1\AFL[eKaOo;R2@IT
Q8_W6IS=qg\S>mEZ2Ec\8WV9P70DBSoG_f^BOk]=Y;28UgC_gI^Cb5GT@=OmW8U=
;^bRnMlWTAN1?3MVTTNd?cPdb?`?^X>k9E^MI8882NdIlVhfo;6O`24_beZ^EJGS
0Tk\:;VlagN8S<h?SUI922dq<YOZfQWYgo[7>FRX3j=pPcdLoch@ji1T58V89Ia8
6OW];K`jF<g1CU]VQ]b70a>43kZ>RhJnN9O;Im9J[IiUS9WeQ^Ejmk;T@`[<1Id<
EFPE5KC@4=T]C9RTN6oF::FSgXh3N3[H3T23Gn?ShSdQP9NldPcg4nR8Hhq<@JCN
e`3KU0>i7FBJ3`j5V_G[9;848c6mm6kFI\8dnF5YBlLYCRCCJ`9fbIOWMlf[9ZK\
FkjQ;lCGE?<G3@>XfB[J9WAh`eiJG=m2];UL]UO;aKS1FKT[`d@lFDh5<C8<9DCF
C3XPGO49<qfUX6QJYD97>j0>;dJ^gQmRYIgYA=D7WEa5`=mjmfoDK6H32o<o:AL?
BO6J<Mm5:VjH\Q?m]>_dnD82^1?FZ@4UVh0Y_<cMZlE]J^\72QZ:_]RH1j\o07?M
W\j:l5Rn[EfHj0XAX\RGNg>^pH8EEjJo5UKm6W0Tfhef5Md;ciP:TON^6M3kdIWC
:Ca@_fe[8\PS\J_S9oOWoBKSkg==P_MkLOfL;aO1KOW@cCo^c5P2EFdmk5bS3efj
Z`JSV^E=loV1fN4^eC1R8fb@MH=9d^ODl93OeD>qNM4Yk^dXKUSdl>H3l4DZFc;^
1>`MROX7nnX@6gTael:U3AU<KEPiC=`IQnSgaCBal9lgeFo6^XfKa`hIQm3PKHoo
G>0>S`@4=i;NZWNASn:dnbII7he]JV7YXoUOg86]N9jmD6ce1U8HV5qME0aGmMXV
]8aXngVSC`YkJ^NjNIibAdjm^;Hb:o8pCXMePB^@Z6j2=_L?TP@@cNIXW=m\[e^F
J_Wg:;]FaTO@R]>:nL=4ObVljgVlBk8H9jfd9nBe6l@61@n<DTIYmbXMRhYHHXp_
LSnUMDF>PB2YG>ReRQ3gmMEN^fJJimbdT[k^\][1Zb5LhRhZ;7b>Sc`gH^0;ebJY
AdeJX`NcE_L3@dD^`i54LU_7^fJ_O1iSLHY88B]mb[>=H3be[Nbm]c?6`993fQ__
HOn8Q3D4Q2`D>qdR\YFnCa?nl`=b<<=PHGBCE\C\9[TDD40`HZ;HSLCH;Q?7RJ`H
_a[MD;X@Pi[P:PK]:\GjN7CVelQ4AWo>MWJN6Fa\bZoUNk34eDnYToLnXSY:[JN7
aLIoh\N?mH6>I]dT6m1UfZ[\NRmcpo2NMNkI<cPX0DU26LZmIL\NJ:n4F\VUjnXS
fgSjZoZ7O>\bf8nJkMBiTWC[HpnBI0P5CPGAUJ6NQ6i8ooNIU1j;^MINiAL@C@7?
?87loSWB^QmR48M]X5KI:EZd8Mc824m5]8iRTCT6YDM_n_4@Eo9;LC6@d@>LFQ64
8m@M4?2FFb5K@]oQ=o52ZP\BdBnFm9ln1I1>i5njqGJkik92n\<h<WG3lR9_lFLm
aD;_8hJEJ[1Wa[Q;479TmN81kRj=1dTFB@0I:\P_^7hLT47;R`ONdX;QD:9>nWfH
bC;:89b@bTjccAI\=j:A`XAmcNXlf8j?kWmNCN\QfGKW_T`aHbnOU4[pb81HO32=
<1Y1h4@:POAF9TNlM;C42kGMK8R[;1l=WP`YUKBJQkfkdfeoQ[@O<4Dj`iE4YDCf
Kh_IP__PJOEFMe\@A;kP1TNZLYY^_GooICADm::O6fDJk?8dV`TbWkPbbPc4iWbm
U1@cW2q\@S3h3:M>MhRlDnR4U::5]X>koVO0jPGIjd;gkQ>7DMR0C?@`IaA5c?88
7F:SA1kaW?5YlFP56`4N9T0>WO?X^0eLoOi3HaoDXP?JETV^>OD=j3fGZl@2mPaF
YNohH[m\bd28LABeAbn85qFK5co8CcII=^dRG60_C7H@mZXkULeT:b1@PgKMH7Rl
h=PH0@I4\C`?H_?aCM6d7\Fl=2SVp8^?D9heYbYVK^lM[J[7cjSIi_hJK?abI4F3
ng?MGoJ=XP3>ZGVo\<KSPO]koFhfcIhVmZKlD:jT<bR`Z<1l;hDC]Ch=Vbh@DKD:
HnDTnETOYb\P1`Tonc5?PPho57cER8f6_PH9Zke\4X`p17gSMk@FNFn16G]^i?o6
S[GK<J3fg9ONVDgSe1Q4Mi]VSml`mjC]P5mk?nGUj[dO2_^_E8@4l_NdDhXXTQZH
X0gAOJS6GB`K1MP3?BmdH]cKUGEiVV4o4B5i78o`;kYT1bNE\PFM5D3K6`qZ<AcN
9;Smkb?amdW9`k_4jojVhF_Pf>IYhT7XhQV6j=i;O\LcAbeC;GO2d:B;IngL[2i0
gaJ3eZM76G@]6[]]1nPb9PV^Vq=dFD`Xm`Ta0]\X:AKkWTk0IdlYR0Mcb6j9k\c@
GAcBXq>^LAa=q2oA>enA$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR4S(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
4Y7V6SQH5DT^<hV1LSDRWJ_]j;[I90;h_UA`jfR@IYE`2=]h5naNg6emKiI;nLin
LJhAJe1nlgpd>N?8aRU625WR?U6YlT\290[D]hi=;b<f\Pq5niMgM55E2<3Kk@_Z
:mg]hEOV?YX09OK7YWdM07RZUiVFQKW34;U4Vk\Zjn74ASq9`fQJ:pV6k3GQCDVA
LR\G8Tm`kIRkPH25GOCG2K?kaYAcg?>XZIMoq6c@5mZcpL=TF:G9D1@jDU1d_h`1
Y\JS4U[RioPlPJbhq7SeD]dpSWDo_F5@1NmBHj?=iZaZWVRP5M6eTKTQfTm:Pi>6
BlV\T`LHN@i;e_4>9nANSga?ZQhk]R_2G@Pb?X399eX1iQ\1oMTQKBoNEmAUY:;2
7P]nl_L<f3B4K@j;j?8WhmhHSQ`X3`k1_0XS=PpfGaRWVOjYGI1@ODI13H>@An<^
D6R^jmdQ@;TPg_aaPJjV4PNh\?2Q57a13?4mMjcegj0=]:7C<6;692IO38o21?lf
DhPJ5@aeADIkoG4^B2Ifl7R>\\Q>1nf\8D6B0FffgUcPmS5BTY8C[q_5lF[BTk^L
YXWWi[`5KV\TBL[6PBFV^Sm899YO2LLMhEEHIS]L3ebgm:n]klnmm;Y_`nAXmQ@S
`e2@[\5GRdKi4Fi6mUHU]1L[b\cUVmRoBbdP9^5d@OkI_JhkQGAEBD__:^]l_N=^
BNlDqm7LD[fDXj?_W4k=C64b>:G[0IeAY;\79R8_=kQTl1m6<Iid=<\bQAQ3\9A5
:0QSGR=@0]`2F9XofN_]^;0^L\^dN`eR`>_>d]56M:lGn>WJI7JoZ_>XBoYaE0i8
;P_Zom=;Td<3HQKGo0^qa9NX]=KTRCZ5AU`V2hNA?65fbXiK=e51kFDd7E\0Adf;
ThV9=M0PD91]SIV8Ke@AA]XS<8J2JZJBUN`;]^Pc052JYXKK8AcX:RaO6?7mj\cM
^c6\EaBncAb`16^IH<LSa]:SKA_;\7`AB6q[HHhXL2S9mP6WXHN^;AlRl2^f7eUZ
a4<=>L31e5oTeN1eLK<S@72=\<ogJ3EEJf]`j^?UUnp^P]B:bWT[ZO\A:UaZCYM;
NjfoGK<c[=m3C<1XC`VMdRLo02NLja6\SDL4TOjemJ3AY4Q4MAZ^h=nJHA0]bn0_
HincGKd@@JM@2aa7ne3DGLY6i]ZBjPQ40Nal4DY?n1]^YNL5h;<^7\Zc>p8]<^<5
HlnBWg7VH^Qkm>`Dea:JA@j?\0@>GfG`MWg5\`SmkR8NR4Q3m5`FAD4^0XMbA_8j
PD;Z6kfX_e25GWNL:G`Jh\oX``6d7IJOTf<5RNIj26;4B7]mRnCX1nel1K8bG_B5
hbFNFXi6pG7?=lI0A;RKX]:6eW4c?g6hm@S_N:7:E^dYN[a2Z^3E>lmM91j1=gJP
3ck:e1d\?0lS6?8P>md[Lk4ToTJ\>SCH4mSHg9bA?[?J[:HJ;9ImNge8BJ9RdZIK
@9fA1aZGOGlPJ^\aJ7<W650p^H`lck>_HdEcT^om>UdkjDHII[SRHLQk^n6YNA2B
FkB4n;[Jh2NQ?FZN;BPG>>NMbid@K?WOIP97FKkCdlj87XO_U=B7?1q]:lcGUMC6
MSle78M7Ke`2k]:>0NC9CK@J7EeKKLLaAM4c:n3_Z1ed2CgUITn29^A4dUVP1BZ2
lNGB>=PTbOk?hKYQ0_g?c`ScH];Xc=;mSc5_nFI>_D2?IAjk>n840V[]d0>^lohE
CgGmbp]5WHkM?ADME5C?AWAa:6c?;j7F5dA1^[W?BS4^^EZMNPX8mmOjmR`UOF56
^F5d1ZbkO=bLFN;S;Y2AaPO30;I:PNRFRcBE7\fA6X6A\4A>CO6VZCKfb]c0ZO2V
:W^n=5]k3<BaO_VOd85hpmWgBV7YOK63<AB_jiXjceB2OBfNWF>Wl67^PnG[h6C>
eg;o]11Wf;I?TWXiWCIj?aS94eaFB:kagXbW<TI<@7B:dLf8DOZM8T2P:JDI;WUG
FXK\foiG9<5NAC7SG]Y4bmSW?j:<2FL;UH1qlP\<6\PGiNkX8eoaS>:W6ame0J0c
4iba2Z_mXUN4\?<Q;S=YPGYnmLAiacAR19hn8gWm1`FIP?UlW:5PnEndoJ7_fJKF
3bODCVRHTV0gOgDOB1[S6TK[]I1LhIFM^\HXlgaSiQ^C9fNXggpRlM4^jK1UaWkk
lVE\Uk?KTEXD=ZdGa1gMA3Z^852V;b5AdaHHebNM=aBUP0:5@eQ\T;T<\Ii^4;_9
?IR[:=5<oILQ=2mFBm3JRU_1[DkFCCb_gRjZcNWZ`LDeGfAX9DmRTXSmdKQ=M_Z6
<p;G5dJ8EI10\1mCDi7F<H2Oj;4gZ5X]HNgQYcdS62SP@MWlmio@5AMZhqIbX:7C
TVaLdV80EXK\@B3WZ;TJ9C>iScS]Vlf;D8`OeZJfjh@ZmXIQeOUB>h1M[FQQYmNL
BiOC2Xjh=l2[e<C\m1mJQ>@kSmUoIA^8D;eXT3CO5fD_HKbjm1@ed[HCFPIQa:b]
mQC6jkdapod67GPSnOl7kboSf4>Rd@j9C>4]SRhHF9CoA1Sl:P6KHoCJ:P@[cf49
o2X_n<HC339I?ihOO_ON[032PF\O7VTe424ki`NHC`Ae7dNWdkn7\TdDX<_2lSCg
kmgTXMoeZo9Si`5c>PZJgGlp>m:AWi3[GCKg1ACnI3IWKfhmnXjZjDn^XFoW[fCS
mBO]Q3jMoRDRClEUR4CVeeFn0I\mO45WeS[g>?9MFOTi^FAJ=XjhgXiX;>6?=OLK
O60mAJeEc8ZRnL[m]LSDkVTF>I[A]HCoid^\USp5M0ZYb]od6gDoK8cFTY?4[V]L
;=li<gP2F9>DnWGUbk@C`j]if<85LJP:jojUFF<aXnCdDQpO8in0O:Wf;4cKJh]8
iK8C0<S`IhTlQ\TglP]lKQFfB?g]lnO`nhVm3_bDX67Q;WLAW<Sko16L_E:e?61\
cKC0_lLdK7n]8pLhL>;Wmi0^<21J]M3h>m\7CDeO10liH82^2WHoS3BodD`g>02j
I>4MNScRm3>gV79n0jG;H5RG>CT?JFnR?A=jb3^DDM;?V_eA5f\oOeVgn@Wi>2J6
f7heYf`fEebTMm<\FK?RMEkBpjI@P[^MMV?16E72NHoOce;TSW;=iEU3]Amch18i
[90M?QglbMcMPNKn16G]^h:oTd[G?P[a_\GAKgS_B8oncWS4XW;;7c`cINMN1]Rc
X4SE19H4UNAN<UDOI5k;VFeInj[;Jm8_U\BF8bcpK9cLKZKM2lVi=MI\eBij8>[P
G?fcd3=_ek3J>M6Nd77AAmej\K:nXTBnc?[K;QM66gAiG182<091fNR7bF=\5Sf3
b?dJ;i?h\Mk7mCQ3LP:n?He@UHPD_ncc?ZHXkJF:KgYABkG7Kaf]D6pg=H2MXfMk
;2e33[_ecn=J4j6PNZ9H7]6<HOFRi_;Ohj]::`Q8K9BEL1e0OM^6jki5WR9W`]KY
K_=YO1h60Sj`Iok=TJb^LXKjeg5L3_@jXFRHIeJQBb7jUOb0hnAcjl\PY<0:R6D=
1q=UIIX^n7;h>Eom@dc\YZ[0^3?fcWnm=FEG@a`mRXM2ZCaJ953<<_mKUmL^19?D
7@14RN6=IQ;e9RBImZoJC`jQE<SLEa6SgahmHV9Q]2`cJaHBJY7HkVZ1JOTaiHVD
0IS\MmME5SkWq`0G6nc8d:ekHP\cF^cE[Da5NYKI<9B]^]lJOn<=2cX`AK;E4n:U
6BIil\m<EDihUS5d4>?:me;kE?KUY\c1eHZPUAKH8XH\f4:fESjXU3:_b0d;ANP[
eOl<cAT8kkcCZ`5mn_dWLa5Zc\Qp6J0bah?OUQMGPfZFjX__d2ICIi`JkhYZEbSC
5D@U:OC13G;Tn9aeoiA6=KoNZ?o9T`lg6_MF@Ql`oXAQD9T:BV?2NijOR?ncm3Ka
;JA=NPKkl9I=Fo1<`AoH\k2QSaDF6`aMccQZX\SH@_q^I?lDL]2Xh9L`XmBB2da4
_lRj2WWf[fWmeh:m^aom1M9D]JdG<D1e?eXWdEoQMfNl@G`B9YW_`i7UHNV`2HcF
^I1?ob;G>>6jLbK>^Oc>gnQVhh4iXKR09X0;YkZ4[`2A1;mikQUTgp1kAm7KBc28
:F69jkNXcE6X>fpDQPRNom;R]a>Cfi\V7C\eeo>D74=<M3Nd=0Bl60no8mlSVoh=
;TNf2anW\of>dFX;=PVGN^\Xm3]FL?G9Fj4`dBh>\qk`]R^aZdM]QoOBGF[>TLd:
ElBl5d6^BjbcdZ[GbT_gkg;]K4g9hhl<5CROJUOTSYZ9eoVUaWO9QGP1XW_P[`Aa
19:ll?hZPWA7YFRWYMK;kDPf=ON5?dmjM>@QkR]QX6kTm`<^OQ@ahfFRqXnd=\46
Vog@`NKj8>O7c_e^;10D<RPe?6F5DFMfmaZOohBOenX?7AGNPEJ:HITMa2jZNcLi
6lE:kkSEL^n2GZ;0>L0M:HnJ?C\>9jd967K649ZH7g\l<UkH\RlWI5Yg\X@7B4Ti
eV_5E1<p^mfZ]D0G76;4o[hLjaE@^DPO3=ZWYYQK?l=5Ghc>Oc@oSDTSdg1eE10H
;PXNediG6cfa8B9koJW`F@2dZVX;_?h_V=NEf>4emKD5i\?i:OaoAb8Ac>LE5JB=
eQVoD^CG^jEGHe`PQAge7nqmKiDL`e`k5;UYI\AVef^TROI^C9869V2XleEj\`94
@n]9g>IA=<iol[^RX3_6_EjSZ]WMa2@NA=CMEW_<nP\i[1`[CkPG_2g>hFY]EY]5
3E5Oll0>8KL_o\GkaBT`M?mm>h[2QO?;^nR;Kpm2GJdV22Z[Beb=FFLMUVUgD53]
Y^YgK8ca47X<4_KjKD_kFODPZ_FjOl`X`CaT<a[K>=_?fK4e?QA]EgHO9Xl:3W_]
5@AcT8NgFZd`X9?QRXHQATC:Kk9NJ5hm[P>H03m=h<MSHZ;<[SKJq69^2Ci;8eA0
Y;GdD5oFP4IoU@?ZWlX\lT>7:Nbdj`f<\O9nn@gY1aUk?K5XmQoonG[Q``2cSFC9
f]hVNm07K6QCML?8N^]lao3TmGeaAj=Y8gS18=Wgf`4k]QlJ;WnAU6@\fiZ<hUOE
6MipJ1VMH[JNJGXmoSp==O8Ho4>4ZC8mA:;SF7bO7BMHko;1EFL2A=B?I:Q9]=V8
6:`k38\XZE<AFcQNa5do=SELXPWb[kd;f[B4EE^0hA^Zkhf8k8LgafQ\H<[U4XYj
f91gC3ialiA8H;^_4Mk=f4T^B5AkQi7iKqe2@A;[_ikC31\5djNi^3@8U3QfKmTE
jW[N;VSIXVDAa^K77@SC:7EI=iN4Hnk1E:RMgEG5[<W@OmK=VnPbb2ZfB7EfP<RY
cSOINkZ07TYLo6d44bN60H:<0DOd:_VQGleJOA:P<_jX\Na^po8nTEK5I@gh@edS
<Ed^YeVc0]ejoE[SFYkJTAol=o0WW^h]XFE5I0\aO4bHD<KlXjlca`8DcbiP6=G4
`lL[F7g::^8he4?pcWU0U@p<\]d;kg$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XNR4T(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
lD<R\SQV5DT^<d21F93>glT:X4Nq]6miP2GIVYT\3ZS\dgHjAbfgPfC`9kc27Vh=
II_V>>VD0aYGQnV6j>ESkg`jqC11\CGfgPIe<fmWaqGNfR;=p:8]jP5:C7>TYEc^
jKDDhXZ32g]2_\U>ZPGLhIaIKI`Q1WQpfL1fPE`qF3o:EmqSXQQMn;0SohTimG?9
a0NgJN5>KJZlWF_;0WRRYEA_E9o1U_MGO=\9iU4LBMnZ::>UF8hZ6^?M`4j;8GlO
aT\]_Z@UK>2U>aV=bGl\kG?]6ZI=>IVD1K`?JH0iM]`Yl=PS\ABoM6<36VUo`qWB
8RU0ZNleR^J7KX4F@Y`Z==E;G3`k9=Vd_Z:g:^<aKD;Q1F2CaJbgHild60Y5MbGc
5bKH5G6_[FV_Wnhhh;b?^Q3;F01^[D?UBdijgCCT3ZU0O4HdnM32n0MKMj\FR`Wc
>cn:2lYMRW;XqJo\S<?aM`fEGiA?eA]F7`Ib_i^59n]Yk=8gRh\Ch^IkSgT<G<fE
>3C12ZR1JblOJ3gj6fQ0YClX4Z40jK432_6J40^`9NVa9kcP8aU8?C5km@>hL<hS
_<`;RFRGgLXhZJX5^PJM^>?j1@Iqm\]2c3PG89Rih<nR?Nq13M`]Hm7gK^DaoLBE
CD7cUJ4YX>RXY3j\_E54`mBm<90K>\oZ6B[]iFJ<1^1A7mehjEjP?@fck:dn4Pa`
jIim`AS_X`Cd^lTNG`2_Oc7HG2S86<8?;=YYThQ]FiGDKj^1j:jC1W1f>7inDqNc
EcX6mSQMc6h>[d369g^CP5OH\k2b6H7hD8R<E>?:D5H]A`D`=86R@jbl2jXRH6@m
C?0dLeaaVHQPPkSOnKb7OGWH7LEkRcXAnj1Nh9FalJd8]c^M14Gc:61B?3`\1MNm
bSNTj0cYllhAqX90<JM2m>l;D4_QJWI\Ohe]]e>j@EjNZVXVK7JNm73e1?_@1oY3
Sg7YZbEa898AC1]g735`KTMDn<\j2L=Oi\\c:M>Qdk99lYH`=LI^bUEPhW@?A\WD
S=llfJ]lBY\BdX]FEYm9gWl9i[Op^<ZUXY@B6fF;im3b_\CFjAG5Rg_@flAWjjmU
OP30M3bR76SA`765d4k9RLm\[cN18bX@QT_T[D5QkP6ic\hFY8UGhg7kU21g;m[`
ajEBF:P0^8Ngk:]?Jf`Il]\JkgRe^gPbAk=L]L@dkhpATd>G\O9n1aLXIlE3>f?N
jYe6:n;QPDZUR3hGEJOo2b\PkR<B6N>qbDMccU_HY;nBOFZe34DejZl8B4@emKXM
6WKDdDQaVdLfWK>bXnhbT^3ZB[738:Q5N@6aLWCcIOVl24NSA4kEdl`bm4ik`k3>
\8c_P4VB7dL0PZVg;PmA4VIf]iBYmoZ?b0AaN3XAn5LdabqO]aW5laj>GNKbU8_g
15e5SQ8MFko?Do>?@:nHgnhDDBWfS\\UY7b?DiRlbc?eB7_9g?TaM7`\5W`<3SkY
1Llo1MhB[ca<YqB?JioA;:d;fX?oHo]LZOSJlOFZ>k]Hc6EQiheP=3^`7A\kOmXU
Q2NF3\H9a]]WI1NY6a1Saja5dci85OJc2G_1Ko\ZTWBYJZI]6Jk8BTjm9@dHX3R=
6LXciG1[VBe;LYBlHET50iBjEM84pD`Fi>RRUmA=T<jDYb;fGZBP5GeJ3]PO[Gnm
=Yg7U9GHn^cRHZ]G1<FnlW<cFN]Ub<m@kV4Sm4[M3\cgLheFKQ^?6deS:JCP][B>
M0hJNh8DFg_=iGBmVZ?]<c4iLFXUlD<LaK]g^D\5lTTq^Lk8O8TElIO6c8ogPZ_G
P1><0K2B;TLdT6LL:I^kk?Pfk<1R]nnAToMHLg5[c3:heGjD@ed0e?ZA_6_97O0L
_b:WBKZBFP83o4JWX>_6Tl[UlfEKmPc?Rika\BaF0E3[^gFXS\BBX`n`hSqZge2V
D0N3Fc=Mf9jVnqM88jB3YBfH_\o9Y_Abg:e_XE7oa>Do@0o?ddUhcg<j9C[`Hj=;
14h>CZS9ne<jIT72K1O4Jmh?ajX^0[\17Y>H=6bo2>Q3QhjNOP5:VBNK02UFBIQK
nNOV6]1IYP13;OM[bdWIgQmLR;0>p6gPB<XH8PPP[791>45Y4609E_D;iY3DIF^Z
5BB\cOHPJOglDK_beKY<5T55>mK<cOj>Hgaf3Oa0=LkenlBhBG4\S7D;5?71k>Dc
AU=BK?l2JO00bG4@Ub6\8M>1V@Y5^6SR=PeJL:[RKX6qmUK>YMZhYj7_1cMTWTnT
TYSPBboSLMTQ0V;]2ROn_Xc]d38i<kK\I^XP<HC4_NGULcoUJ4?FkMo>0R:BLe74
4fNE<bnSFoDnGA4>=CL^9\c_fKEO]=aeAo^SX6X[7n1Pm:Y2=DjA<S1:ZmqY]FD=
nCom2g:QN38<F5@gK[@^OmjB^WQ1A0^fT^E[WY:hSfLaD<9;eoIXHN42;Oi:obHm
PfdoOJa1YUfl2n81PikcOgDB3ZgF089:l<dCBV;9Q^OTPR?V9aKkm^P7[WkY3S>U
Y[kl4`6f[pKC4f_J<1?^=>CD^2MESSV;[HJZ`R@l0B55BVd43=BcH]9B4c1YH^JT
07mCC^:YOHk[mdVE3[[hKL[G?B^\mFdOYALZO381LkY0L18lL5cLkYjhf\;YoAEK
`nPV26l`K<Kl\RC21@SFS[F6qX\amgjHi6JVaJkF:gDFOR^9UIcGh;7f0<Yh87T]
9@6_eo3O>?VG6gKYhj?NiF7Om_LJ=^<M::V8TmOoOolXH8VfNK3AIZ<p]cUHbDXn
^8?F?3;W=n2ITeq>3iFH5Cf2YiM5aMX351M@c3a[;68`GQ?DDd:<=jO@K\Pn<O]O
cHH3[`UMK:h<UlBf`_E>:8WFf=hN26c:djO2JGXe;UXW9nlQJVYCf^XRZ9oD1V_H
Dg`_JZN8ia5gCe1>`Qo:DRPf4JTI=p^a66@aa1?3>7cM_YKJkdaV4cSV0CW]Cm_9
n_6ZT0jP8Ti[LR[7QFgZ=[MU?m]R]E66BDWECGMa8b0<jCoV[``fF;RV@>^oiTEJ
]m7co<k9=hPOW6TGY9id>A4:YV<^BT^6ELRmnm_lL4lBqEF5W4^H5K\FR=4=XGlT
P7ZRfBA3^2Jfh3V[KA<HB24NXWUfJZAId?Eon3O3BJG:2[8nXoCegeAAKEK4BSOA
nPBlf5A3PFgbN\D3c5OoZ\Z;8B<5NL\cf\5mcG5ac0:jAE8A4:@Ind^YRXMpX[lQ
D4O5aUj;hZjan<dfKIKkKol\\e;E]m<EnZehf>eTJF?YJ]:0SXdhhndY?KQAIh]P
Q7FJRgkY^H3mkfKLhAH?ioKGWnEnMoBT2C54F6OVmeo3`]3GbDE]B\h6DBD<Xh\=
<QQKlCM2KXpBMSlIGMn\U=DSP0;:l^o44ONiSS:Q51U5?e`AU=XF3RGSSdoQQ<SG
5\RE>NfHh>4n=Wc[CaVPZUPTPCZdMMZP0n>SSHFG;3TL;\P:P:ZBb[TTZWJBQO<E
@hR?ehJADm>B=5b`mR6XmIX@4p_22[c=RC1>HO1ZWhUVYXjinnWWk@AG@[ObGF:j
]ej\1^S78L8De5eC5O]>:CJ;[>_L\>IIUmmPhBmOX8nMAm=>FJ=WH0J72lFTfY>S
H<oUIi6A4cfn][o9^OK^VNHlCl_LW3LJhbQ39>3]p5cAUHAmgZe_IB7=oKQ2kGl[
k;4nmDO3Nm<VCIZUPRT75mFMVoWAWIP\8a`Q4`NnUk^UF1eX2e4`?]3PkKm5V6eH
f44n_??J5Kd`BYOe;6JgiTCQ>XTXXd:<d`JGHULB65^^n?[ole>24RbphOc2\Ak?
i?NMK]dLIc0]fXkVd9E\KYN8Th:MO]i;7UeRWMjHIRC\YINFmf4hZCLkZWBaj_cg
KW;VW9fPb:oS4SeL<9O\oMJ_L^]`9LIHdafkl@d^__6Qcl<=jcFV]JRahW@bHFUX
Pcg]b1qN[;\6e?T=UB<X03\5[D`1igO]g\Z7eJB6KHl;R2Sb65YF@0khEliVHq?g
di=RE<7XPUJ>VVPMRPL@lIJA_XXhmcaGaQdLX3J1`CUI?;MoGM>_SfiJSoPe78`D
k4KPmfUU3P\Y`A9`MT<ZM?1LW4g7pjdX`GZB1c406b=F]n<K5B]IZS8Pl_FV:V:I
\;LO5j[\SE7maSdZOJa?9O]^6V<3bUlh=dch2l]^bZ3D\2XjaSSB3X8ejO8@P1mC
4k`[DMUo=>4<UOXcKZ;HS\fS=Y5`lj]bl@dZCOUf:66qLL01j[P`J^3KeL[a1=O<
cZ8OjBRki=IW;UfCZEDfZYZEKO^Z9OlI:U=LU6i0EZH[HKEhVg?l>7l3_83h\_7d
Af1ATBfiWogJPHVZ?[<jf@ZJEMA^G[FJ1Vo3]HdFdCIfLKT26nUi[a<J:ip06AB8
fiinS8`5@8U>faJ2_VgkTg7]S]blVCS6=6cA99_QBU1E>b=J^J?dWWo6C_]>lo\7
6\Pj[@^1LN6[1ckdo\R9Td3TeWQR<cWT6n`\oQ1D70]aScghf9]0^gLj]DA0l_`d
HNLZDRNbWpRHbXdS5JDSIAERL\dFEDh^6MSlNIDUPpU3eKABg8PGH;S4HK4XDWQ7
U8nRKd[>_MAIT@PFC8H[3=Tln1BXLYmcZVRcDUW4H738WmGW@Male`A`HE?QPci`
b9fRKPLOCoh2N?Nh7YXM306PCJA=@94g[671EaXQX2UHXRLCTGmM]JJCp?dIgfRZ
QHjPkbaNckB<YFXMkMVjCK0Sh2YGYl^WRjcbP38mh1SbjCIDl;QTElo;]gm_]dWb
N5KHSF\LNlOn0N5c>>V7NgaDo6IlCKdCNe^l89lLhPo@RXWj<o<AY[C?S?aPgR8\
GSlB\]Wp=L6C\Id<QcTDD]I4nN:AEM8UX>L^A?B_jo529?lA6YI>ogI2>_TLZlgV
A9kMfB_9n<1A@ER`VR<cY5n;PN^X=V^J_>A4WT?jL0n\n0_fMimVMh^1l6UCW2]I
ELm4@7jn=<n@?9kbKloAZepeS[o4UGNLahARP]>CeCD]bNIKGJKnn5hDDT=HT?0Z
Mk4oodA>;YRF3XXclD>BZBT]NB9IbjI][Ai?V=_93VBUF97bGUnRVZC5EnRcAI5b
mkG7^MfC<TL=kaQjh>Xm=O]eNh_UWC<o;EaMipMm9H21hKI?>ad6RI?L3XimKQNN
Glm;QFH]i]cjZDDL>j9`1l^g5Rdl\ciL;l@nGjPa^4<<3Aof1;`l21;jKUoGlUNN
<<Gc8WkK@:oO8[TFZD;dB<4:@^G^n\^G572EjcM^Wb0j5Fo2fA1nqL?J]efWTX@[
Wld@kO2`B8?Ql7N_]>k[ITmO<k10JaVBH?bb6]XY<=MDj]i\HTh@8ARSO[YLFZQD
>eBU]]QkPB:Pn]j?Xh`qW7m<;\]\6;PC`Dq1K0791pO6DeLXV$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR2H(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
6:ll7SQH5DT^<WT:NMn7o@I0fhXAOb0lmOHnf3Qep8jmm`AjfHeJiPPVMj^L:n1B
?G6MES?PqgS02_`HGf0:H8g7kMM5]9LIoAb^_mkU1gLa;_9`T\8SE0YqCk>;0cq6
`lNkP\=LAOT56OcUb3J7S@DCM9a`8G_p^Y\F6aaq9G2GPF`ZWhUJ<S<IIOo6I1=B
IA^B8]oLR@qONbjJ:pSRbhZQC<4[JF9@_a?8IVLZh6CFnl2L@5QRce\ce`P3KXF3
@CBaRi_BH4[<187jidSJDm0H>[?<BbkE`K>\;80CbNb?TkC4@4bQRP?Bp0N:UN67
`SLgkVikSfK8j>[HbJmVZhJG\`<M8_X@_^@8O9oY>TdDHR3\CcTR3U9nC0eX4d9I
eZ\=XjdQBcP8<moTKHFYh>FG[O`MC_Pq<<I8eYM<K^8bGHD`JlR_WV`MI0EE_E08
RRF7F9;B9]bBoig2K<5K8ReW2iJdQPlQ<^T4nol4[5h11OA\W5KDCnqk12_1h5mi
@4ASH]=OPKn4MkXlPb4dCLf9?a1;i7bC;_85FVcMZRdJ<2h`>kIR5GWk6NKYMlGQ
ET3K2\^mBW[125?@hKCkjLfgFleQmqaOIOY2OAeQUG_RTHba7>;YYcJ<9IlX\4n;
]cgV=anSOC4mG9`SnEFPlYO;j?V>_ca?KgJSV@XjkL]U^j\a<CSUJ9TIb^gf\4?0
aFX6pPD@`Q\nJ:M=Q@WSfWV]k4:>Qn[gfLj03>Q26>ZI8aOnTaNV9lN49Q^<n=7f
JH^AeP\[n<S>KnH=K8M33248ZE]p9GP`K=pjV0n<\X$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR2HP(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
=E_T@SQ:5DT^<_>DYaCQ`VBUoHLoGcWgacLcK`3m[L7F8K8`o;IBe6qc^6TT;aPl
`Q`cB5lnAU]eUXI>kHXQ4ET_NRW6_FafPTLKWh\WLk9mEg59:LB2<pa3jobk0`WD
0mc0fk]K`Na7[S85g^0N03a<BUZXm53[MBO4PZ@8p2UPS``qLfL3FdFoh22\1e`T
4]1L]TG1H7Qkm7mlpXj2hL^eqYYdR^HqE28JSXTn71n[Z@JF237Sdf_GmOPRnm7J
`j5SB;_NIlm9ccdBVi2gDOXIljXa>><XEA>7=N@aWnP3OAWDA7Xkhk0Ygo2kY`7N
d:K]jdpZ]RY_3hGf]ZmD1KGd>HMOhd7IIEn99\[og7W9LRGUJFLjkdhW^nBKT9:B
`]GVF\EZ[E;Q6]In6_GiB99KnHOgh@XWiRge>\hlOLmiBqD:0=gALZLBMnHO3@jR
G;7=b`205enN>OA[Je;6cIXd:34N:KI^U<;5Pm2df=d^_TD4SQX[]jGFF^:d8W@G
3HbJqJXlj2h;3NmfH2LRN@odC5V3lbaH;74Ue3JJ9K9I_dZ[GUBm>CZR25knM>lG
OCV`QJR0fN6@HXYIC9[1b^OfXdVETI1m7V_UjXCJF81pPD:BZJZnIfjT1n_0:;hR
aKRe1477nk6<kVSe`5R:fl>1]NDJg\;bAeAKL3IO`0TjPW5i^`84JKMXNZGT^WUK
:_eFBGRfU36LjdNPI?q?>BGk^0J>9A@ljC;p:95LOOYk7Cd1U2CdBeE1L6IDU;?k
8QBa245ZCZ37]FHi?QLa=gD]I1oJ\jSM?P`@:_Z^G^R:kVMDCNDk_hAbkWq3SQ[n
gqT_A=JZf$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR2HS(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
6gIE8SQV5DT^<Y1Ri`R>YG1BIfb`A_m??Q]1lbV6:<6=86^@\5VC08:;5EATC\AF
HO^`qj`Mg:<0gM>WOZY>KQd]>ea?;b3be]Iga^C91SM<5P>mEE\G]l1p4iS@W]j@
DW3h5kbK``bXaIbZQfM[k=9L46U6R07q]@kA``qB4;SR?2IibmE2Um0aL;YDR[Ad
WbmPm:Lq0`L8R2Kpi8kk2^qTe\Xc4mP<gZk4f]:>GQ@<hEHZAa]dLJ]nV2N:3A?3
`3FBY^8S1==0=aZFBSEoWYRT^dU?BhVI^4OhIEVE`O;QBK5a8Fh_BJ?PZXc7hqC@
V><@`9U@=W5W7XPf`a6Ok2`E7YbLZ:F?FD>08i5o9C:Y8=>m]LZY5h:X4SmZGACA
E:l5eflYbOmN<8<n`f9nYDWPiS\2Z@>lfhOBq4?YLa^@neeka2XVGhgQBS5l[:A`
RIeZR2KmcZaP;>@bC5I7jYZ:jMN>aAQBNJG;o4BXQ]N=I;DVL]4Yj5ZMUhWqDO[H
1=n>VLVELG7<c64End6Eei5bLnh_4ohK8d`@nnb9@S1@miD7k^CX6jI1;MdSDAhl
QcW1c5X586ei>d8X]J\f1LPWI:h3ZKGXkCqcF6Am>iVealHd<=SSgLC3TKIW@Pg\
_b_pP;K^lW9EcJ9NQ4HlnLZjRBf6_F^V<:kEI_OGY=ZgEo0M4C?2T4k4Bnk_VMC@
jD53PD>MY?mZY5TnMIb9G2BYBG9R_:YbgnkC2KEV?bq6iK>J^ZVd\UQiCmnkaQgY
UHo?6oJ6AN8EC<8<f8612?Eg[4nc4?U1W\12Pk^dgJQ6]7V_PDP:;KDl2c9@K7;7
^pVlJCKQp_e>EU\2$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR2HT(O, I1, I2);
   output O;
   input I1, I2;

//Function Block
`protected
VTO@USQH5DT^<h=`7m?minpP15cFP\bOhm<eg4f@aXXh<CNFgON@HBGY7Y7M]CB8
?MEbS[CQm=9n>9YG:o3g3[i7`a>^2q6>mOo1\VLD:Ck7Ph32e_PM]1HHPf:i^gol
1TW>6Ph=WZ21qiPV:4Op=;OYnN8]B^2]ZkI6Kk]A;\2E5Geh1I=eq5;Wfb@Zqn28
`?>p>`J^Mc>40X@Mb6A0e21m]D7WA7Jd:jgX`nBGe?G?WZkA2@ZJ<fG;^a=ADN\H
UYhe>X:Qkmc2FMij`3YVMT\?fa23@PFQSPgfX5<SkmpdRKnk=O4ZgO<hMY0T50FE
>QVV1`Ho\C8G^hUo4CpZoLNZ=`3EblTndg4B8][;iFj`^[5=dW:G4CniNo=VHW]o
_7FPNj?^oGI=4J53S\PZPVn9^EDDVUe;\hom?]M_S[\:??b0OW0Io33>7qNl0D?`
FC>C:Yg8eCHL9n_=JJie98;>dGb_>]=]XkV`=9]`PJNSIYg]Jb2m8ZYiWZNniM[A
c[;71EPj1ORX^?ICqYR_X4<B\i>HO3nlb4]KjA@P\5W?LjEl4UdgElVKY8@NQVk>
j[ZP7;g7_Q8?0`_@aYUaJTfMiM<>6U^\F=F;cL\mlBe9HO\lGOLP^1np\SkM`Mn:
]I?G2BbdFZC81mm`<GE22V324D6305TE9PWMaf3A`1^oh?1HlcjVH1@N\5RDb9U^
AfecK@`EXHA9U07NdIUjdi3\0_^jIhpJ_PlBX38CZ8oAlZ5UXcjP00n1jaLJ7oGa
?F9DH0h;\o:G3c0\0^:4:b^^CA7@BEQJ85^1[?]FHM8Ug[iEb`O00qSX?ACoqbYP
>9LIh?1D_GO^RRakQpJ8\kR^8$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
AjJhLSQ:5DT^<jEifP`=YL@W0HggAh0^E7`qHMVbn_kGI6^`gmn`;XiHKIC^?66G
N4ffHP]8E2BEIdh<K7cRZb5cO7P_AoVFHI8qX@Mj5FCKT0k5PQjBDgP0n`@9p2hL
PNcp03K7GQ98mk]aKN_[lB4j6o?nam6?GnPP]goLG>Rp3FM_[F<qMMDd8LpOUn53
<b:5H9nPUfPA@P6@=1JP=jIEQ0ZB3McRiWmZ5BQA@X>^842RZdDOS1gR`DXpSXD<
FY`[j_AL`BPVehWUFKLRni_]J=oe6bh>E50ISO>RPHifQ1FL:PIVQkTSk6]6SP\n
2`9@QWWikmQ05l=eG5^RdieoUC?nZb3V;2hRkNQB6ZolVYd81mqXlelMi?QQ^ieb
Vof@RM6:BDiihLAfL2n\=:cj\S7<MKHk67QVK2glO=J=GX]lD97XUnCS`<RdA]Bg
;b@i]38:=FCNVXN?YV0:=`3idO^2R9X;XN8fJ>m:[pE:G8CU9c5SEWm98c[Fb>C3
l9LX\m^f[EAk^bj]o:hkO7BDJS8m;<D8D_BC4^8W]8EV@4B<X6\HNPSEikVj[8X:
aEbShhB9fcokYb?CbiGYNjZh@IC<UC>2pj5Bh4:e80l:2aSM<97U]GfNU]FZ^Q99
Z>3ZPXZ;V;YDgbTmI383j4bA:JY]nXW74jOLZ:`_SN8N>iP_KlnGgI=>jk:MY[KH
4X3BMeTdkQLRSD2FK?>6kbIp1F7`?DhF\UBH8hk4ibG7@id@nORNTaToOX@30h=X
=MM`_7FgcjOVUB8\XZPL[6Cg1OF28l[_^I:E=^hhJF6gcNqY@;Q>?dGc7d^D9FcQ
@XRSJbDdc:2;mRX1XK09]Y;[Z_AeGAOn0FJ9Zb;=1jQHYWJe1Y=`gU7>VeZ7>HSl
XUcIgL^;0P:LT97=nc_D]cdXT4PKmd;lkLkKd<Jf1pR>TcjbX6h[YF@45`Z8me]P
K@TgEajAbQm<]6]gnY2eDZb1Mm6Km7_ji?2lX5b\gd3783\kMWl<IJmI1l9G:eP;
?k9e9=4JdoLe?g`bi_lNW[T1[?1eaVVngOJgqdU;6R;_^=2BoVbD;`^_[Oa2K5AJ
N3QWCeEPqTojR7KGl=bl`b<IeWdGXN?VYBiHBfhK;eYck5U_fWl:Am\_7I:4h_lh
nl0W[FlTT@IZP4S<aZMZ688>iQHbQNVQVGXcK?Gd?EZSoWk;?2mOg7RO4AbGAoC?
X24q08DO@[9Q4YaJB>l^SUDlEJ_Y0>H]U:jI`XbMnPFWlMR\EI8Hi@PG;2_c1e\Q
5j3MQ_:0C12l?<eH8A2G]TF@aD_10d?=jgFQ?Z?7`PknkYAYV6=Jka9EiPZ[k=pW
XM?2EQPSfH[N@TWVO2CN>ib]?2g:ioHd9n2N33^\2E_RNDV;b><^=`Gg;7ZUU9P8
<_1knjTT0ENagVQ;=^`HiY`G_q:8@6Ao2A6oPoHCcaV_:PBEBBfR_52b5VEE2mhm
mVk:aX<]j7lP`>2XBWC>S;^bfh@53:B^U=IkhA9[WNEP6=aXo8gR9l3WkVbi[EA;
8[I;a64FZ]:7lnk=F3GT;EQ]pg:oJHQRW9SVkBhPe\E8J028SMAE;_N9oZXJQX:B
35`2GK=olK[lVB4mIH7L6bZ@<M[::7[ASi8g[5Q10oFeBoaJ^SA;>L]\[HRRP1K;
K3cIDNGGeYGR0FWTZ3eDGlBp:f@d=PenRo_X6<iaGQMEP?39=\]FAEDUnTcEbLbX
dbP0gBPH[Z25C@P5QSN?]PnI62XjFA>F6Zb8YIm<?9_Y<eU:^\fh;H2Q^4lTEPmO
lok_cI\kh6lfBf:W9`ROTOp;iTiL]M3LGL\9C4>GOS7cmcPDCBoL9l[i:EfTR7bS
[Vda1V>\UE\fClhhiNEc?i\b6cNg2eWPmRjlYF13OlR<1K8KDAC7NIHEn?SQRBRC
lakG??]Km]RcS`o^CqQJ7]k1LijW1dM;2_KfN?W_oQFY@RGKV8TXIY1\7FOHLKf9
n7S:]fHk861kV4E^C_FR8h30l44G4k[lC4>WXHmEgV;SqD3G_`:pPF=A`]on76MD
F`D4mWMFOCQqW`]3nFe$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR3P(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
D81^gSQ:5DT^<8La]68U@0HTQkk^XBDJhO44elWBX\i??O56q\JlB=5\kYaFQi6P
Mk[2bmVCV8MTLH?I[F^XCK_M3A9WRYXGoa^K]eV`Fj2pI<HnHgJ:U;lV\6=3JU=4
?O6dVn_=[BcMO63ag[E[Y@FEA07D=h7TPdplH_V9mqcdNK3>TSHP=N;^:EAgUgGa
0S_mTA9F1;eMmo0hnpMhEMZZ>pJOBQ6Qp`B]`L=A9`1OQj`Na0178XgJeKP<\`Y?
i@>2_W5:1N]V5VckVJ9gE>Q3S:2ncClC6N<eUfQEU6kXJS@V3K[;W:M<E:G:GK_L
ED?H]V::mgXE5_@l<QWJHLa4jQ6pk]<F=[;Jh_gS8O6e[l=Cm:4KEUM0^>hkY<Zo
IJDpbmk[SXAI1_go[Kf18Gjh0OaD:AO`Z6__?[YH`X3l78J]\Lih6\BSGZ0Q6^][
Qak?[=8QE=b[`GooWHcDPKd4aHooi5f7Bh^=7K84GXYc7O71H_M1^FFXc_oWAkql
J3cJa@93YUToBmXR9o<m<JfmhaFJOhM67S^9\A=JWCW@e`L:e@X192FmAXZN58:;
;XW5AY2dJBh`S@Q:?A^og\1m=mK]<W88UF2L\6=9AHRI2YK5JHJ:RAih>pgVU;m:
dX49>lK8`W:^QQVe;RK7a7;C_E\U2T\1BX=GCP:o:_N3nIX2OQhn^J>0UN0L6]k9
7NlhI`HL?F=EPfIPSeI7g[PlcT2J1NdE<KjUkNf=2mC0=Cg^l]JaDRH@pWJ7lALd
_\HD_F2KalGRkNFFd1bfZOMWkGH^h=X=VgBHS<?RcBK63\PG[a1?HgXYWGTRVQ?F
?NoQZ9J`^X:0\2T9i^U;b56p7ZSNj[Oo]GfPDePiYD@Yf:;F`BR5IVK_>GSdF66a
Wdi\;>3`_YKZMT]gTM6oaW1n[?VkVLT>>Tb\aTTYhUkKmJ>U0B2J3o?enA6kMPP_
nHiYO2<cT[bXkINiKF`=8mqEF_bO6f`ZeCWNLaFo7NoVk:A8GBW;;iMY;_:H4C=K
ii\757M][Enon3=aYGbIZN4fi@=qZEL:E_;JK3:4Wa1JG_?QkRW;L8`IoI^1NJDd
H^A0A?_^VTL^MHli7Yc1Ibd8_^Qi8iMLB<:l6DZ_8VI2SB<K^Dib\8ZoRDb7RbY1
gCle9eCAkAjleH=Wn75R22S51mpQZa]E54McjAlif42\455^XUO3d4@J\Dk@B`Hg
eBkO]a2oek<i3]4Eb9=gNEdB]dhhN?dF>lE\WP9NaBZ6`UHYb>n[dG01:bNKG6F1
CV^lYIGnkFI63k738A?d;^:2BqFTn6`NDm?ODd4dlCUaV@B[]e2h8T;3F:X8@g;0
NYQ`gbX;iaMd4hI35Cab7I[D3:_mb^QZPmflRS76le?U><gPQOQY2hTmLIj:4aY0
j7g7an;GQe4nLDT\5eMapMSYG_g:84bQWA@P\ef?ejFJPFdHONVKY2S`jCOOl7jX
HeZ;gH4=E_gMMNjb0`oRfln6<^4W\cjo[6d2l1b=1fGPW_op\:h9o`j_6YA1ULj4
n<8X6lfYXaLV_`dmHYGMKcSW2S>h0D^9ZA=MF`JokDA5ji>ATT4PGRBE=Om67AM;
763km2OFkae^Yk;]23MWHoEE6=MEOUIl]?WXkl>AhBS?Smq37XD@2\W@FCNmF2<>
4lk]1\5D`709U[IAl>eHYUH>:^4`CeP\N_QV7JnUZ0PT1Z3WU?7ZT35L\0E^kM4\
kcbAjQ2D`a9?S[^OohZmNe8AU;^;KOja\?6mM4oZd:^Gmp5G3@BRG3kc9mInFM5o
@Wd\bbJHYN@P;PEHSV\Y:WAcRdeok_a]chBWGjJgkXlSHX8C]=5Rb0_1W:JZFJFI
O<NaIU;H4:VW3N[hC^bhRYfUDI;2[^8JC?j^T:UGNRc7q[BeFiak=GiGLWlcQ0hJ
e<2>=EI=Fa?`m@@Q<9lKYMe2`cVS\KDDia>IN_6jBnM?>gIgBFjAMQ\TjQ8DK:_^
4dfO>1I?;=mJ:Co1?UWV4[?2VO04nAV@>2=Pj7=CHC1p[FLbgOnd^1Q=0K5MmT1>
_;B3d3L3O6;C7JkC^Rf41J1^Anhp>24dj;n]FU@oFUa5_bjlo]^@l4I`T=WdM>`F
_a;JlcQR<d:dTD>Nbf7;1hQNVkX2QJ0V;l;SXM>M`i\TZK9^b:?>`BiiekpSTXGL
6p@5NDYbh$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR3S(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
6>A4TSQV5DT^<\Pak_;<Thj?kOMd40WDnF:XRY_;9KbWP<R60jP;Ejo4GB6>Kop7
;ACk\dmF]>EGXZ5hSeAq2QM7gQGVVSTK6[R1k@G8oiBbDj`CP0:XidbHlLThGJQO
Y0fUQghMq]bLOD=pVOBGkILA<PbZhK<E<<A0lP^4aMHF;JM]h00KLgTp:I>aMU8p
C9hCU2eRE>W:?YgLED^DOb9U4OHkk2^3[1S6aJLoTZQ4:ih;E=[Ld1ghL\FRp4^F
47Xpc_bWB\5ADh7lM;2;FD`C[:>W\AEGdQ7E\kk4Bm6k[J;cJi2Hb[hmMf6@:8]4
FOJHc3dW@aH>V^dQ9dZMN\nPDF7^AA6Y7fRi8k3TREKLRGc;gWO=`1O94=qjE[]V
Pi\R_6UBD:aLL<^L]Z\]6nQ5:`IaKLaG78gK2D@5_DPGXoXWIJ?k]W]Q;H]jAI=S
b`3e0Jd@BOO=69n32Zh[7D;?3UjAK>a7N\8J_>N:MeKEjkJohp\[RMK^XR51Z4el
7iNP2P4Oi]Wm]2FTNnLToVWLEWc[DXJT:nmBEoil<hj^42SMLN\G7W[ObbA7e=61
9YQOMa?Y71cmoYbiB=NTADPAFi;C1<Pj1OaXLh?mp[IBEdEj8\1^\RjHRS455WWZ
b7XB?]341>kNIHmPA;@<;MBDk4>_ODlE\`k6DMlhpX0?`mKjAPXlIQga?S5aVbke
>TPgCDf`cK:cm:\P:iY3C4=?>CcAM9kI93V7SmdO]X1EQ=f2bU=iBSc4N>e\2mnI
XD<UL\Lo5G:hT23X;K1YVlh>LIZHM?npBh6;:kdDUMCCiG7ik?ABXiXWAEIhZKLc
MK?lS\IKc_AfNT>WA9O02:J_FNChE[6CBaMUeJhJl]4ORSd>3;g2^1qP8dij;WV?
EB8g>3?WVSRlljcJW[<:3<h^MC1gYbFG8IfK8@]?24CK1<h3:kHD?5<K07;4XkTD
2f320XY4Ve1O9[_fkYcNDMNF2o5XY8fh1COQGG:QYTI4[;46`qgOWL50b;GV1Y>d
57oUPcH49mnQ6SXLi[09aNS1HoWgVM[mN<WYHQILEk03mCjlRLFm;lije[iUjlDP
<2ZkMj0BA2^g?=^]=Id1_VnmY\kJ;aH;C[l0XF`3PNP4p1O7UVdCZ<VRm9F=ZYXU
SodR[:5GLF37S5]K]7\>`ie2GH8dHT9;KZbCfd2e:hboXnU3kLQ=:AKDML<o1^99
:[:>08JU@jRWgVKPdl<YTo2K;>8YP^>\>?SZ`@iqmg2mT?JAbanPFWN6l??WHXXA
L>074XbTHCpKQZ5T3C6OY:\CbTh\nlf=JQQJB9MRGa9VS`WECdnJ6f48?0H7KBE7
S9Qc>h5faKmT=HAJ_573C7eTFG]7?PZ@B]9hKng<X881R1NUCd`1LHGJMnnVS\0B
nNHP<p95VaO51d54JhGbiDAROh?GlA[l6hEgl<6Z37XCooO5a71BLIWc?L2@TQn\
nGK2]=MYGETOA:j:dNY2nnGfQPaRiKN2pIM^>dd=69:<jgH6hmP9S1?W:<]ZjK[S
8?6[0R@C4^I:4Ofjfn;PP=VSidlUJmkH_g:fg2?_i@G=_\X@g6OPn6Ee79]VK5WL
_ZG2WC<1DRjbZfjmPC[Q>b[FhG>AX?3q2RENHfd0fSfIc\kngkL_BZc]ZL`Q]fcg
Vk`5liGYj>R\JM3PWJkMWZ0fRIPfUn:cPUon29aW8eeJX39Idj:;cROLiLYCCeU1
9]=;`G3cm_SODGPU3L4oaVXoF00Z:=q`[?OXWJX2a^5GIj`c55GH7D`b;On7]1=`
OE=G3@NhUV_I3MB45LdWBX=LZCmnmfBP=`7ln>>HQT=@Y9k9Q\k[O11D;jLA:iEU
7XYnZf\`EQ<J^k7A;[GI`[[h@6LikpBoDH^ZfZ;LBKTQ0W5DjWK]DGH4482@nRLG
0Ti\IpG`F`VoRHI54Z`;[nUnTn=>2lgJV^=I0AI^@ldhCm8nPiL050l@Q14\<UO;
l]IJ619WjH[dHm>487MKR7=`l6_9OeMJU5l=H99PU9CdH6DA1W0SC?SmUABCHXe@
dhTJqnhCVc:\MShN]B?X:QKjB\jE=6;UD8A6NDMdG89OK0LTlYF`eC9THC]g5Z=i
m3Dh0;K5CkmdM9;hMJ]V[I:2dcROkE9W\U`pPN=X:`phZQ;UFY$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR3T(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protected
168leSQd5DT^<6HbE\4<]2G@\^dP;Fki2^X[R07cdj2^3O2=@b4bUJ6FG0AOPYHe
<D>=iD0E_ZD>pbonlXmX0FPBn?M3q9eYhF[31`m`^Jh0Rg<9DBZVHYJ9ceBS=c>k
LfCDmVcRhjQ[S_Ml2V<>8KGQCT_DOIKCm@1npTOlo2Tqe:=a[E2lX[An_co][c2g
^?SAFQHE<bQLVi:Sl7hq^XP@:NUqQA8]<^p=Noga3R@TZ[\C\E?XibF2^YMM@hqh
RLonLn86cmSmO_3[ffaLZ9UlmJAcdFjScNDdAfHW\L4<F2HHjGO:_FI91b;DOMZN
GHC7X4``1Afe739:R?]_J3d5m]iWOkZWdiS_Z_FObHd6[NOSlRO@FA[7USWLkpVK
T0CRHMCn12=\Ch5LF7IAiIE9JAO@me^k]A`;f?LlFN\:K=?Z^kkjmNSZQ_fG9[;]
cYlhVSJB`mHSTbl2BI3AmQM9UTd]_f8lM640k8=eNBB_4SNMldo744agK6P[q<h2
dO1C;h[N;UG14\]@9^EJ8?FPoDLLKY7<<CCBJgi:ah5OlBQ>ckm<aYkI@g^BmS]2
?ST=b1ka`S4L=BV5N`gCe5F1SbMbaOXcf0oQn3>:KZ;Pf<QOX6B<k<\dC;nqdYMO
7\E7MmYO=C_Y7N;]I>XDVo<:^T>[ebSXlB9=K0U63V8kANT0h3Oc2hGCe^lC1Vbc
916G<>UjC0[d5NGoc<DjEo2gHEQh9llE2b?cl53Z;j1kL_W^lRNl0oJ>e^qV]Eo8
F<D>32K<:@VmRcI4h5dDGLa8mO1YGKc=?I9\\i[Y[nfc<J_j5c^4RRS=Y9LT]@3=
3T2UjYM4Vc7PR_LX3cQC>6:[aq32GBIoQ=LdI:hM2I>1L9F2f;DW5c2VD;OmcNZ7
G_^kK4>`TJahVLV^S8^]5\W=>OGEo[KG4o[0TJ>3Nn_Y_>_1;eVW]QG@96U8fdUd
HNGE?m1\=caHMV;2Ed[<783Xq=MX[`=B0YY_<91K5c:TGCPFHBn6e>hY;@eMod7e
Po?MBSC?G?2aTJ\QYY;YX>iiWlA1UYbH@nebODeYM6l@@DKkEXnlM^OdOa4JILYA
7EEGVXFd6b2DPFUmBLNI_j=pW=1J1?`HAI7k1[c@Wa1939cJ1TFinCE<_T5?2:S9
K82P;<5>ld6OahVMe^hEaU[ZU>D?3KBPI027Fd_[E;0^X`iJ_T0D_oh5QC[30k@X
mFJlhnjijd0TAmJgAFGZ68p<_4mjV^JfSTaDJ5X\9J_LGomeNA04=6gBSIDjMEk\
j`K=c38:KMbBSGob]1Qc7Ca[=^KqiglX15c\<\0hdOWbCTl;4L7`oHQP>f@9N0o>
GI@31K8=G:2mm^4HWJL^3[D]Em:^HF65_:R1ejElC^b8\3886N=b0H`6CgZgDd^D
eedh<MXEFCJf_V724^hL[JloGVq0:LZjJK43f8TgERDb:T3Hm8;P3OKDZ]=d=G6j
Ri42fHA4\0ZT8Cci=aXJR[`igmOVBM7<MB0LOKTM29K5_fni@dm[=CBV2q3g@[k@
U3@FPKCGH32Bgdd[IH82l[0[ofHPn;jbOLNINVPBYS1l0=BMS8ZT0hnnWHhHYWoU
SWAnc8XOGE^8La_ZCP42U1lbLXC[3;b^2\BGc`=N22NjC\D[Tf0?WY]2pUT?F=\k
_FIMA?_O<\RDc1g>81AhPi\C?mDSi]=Q?0c9Ak68IC\FXWaN3T@:]lYcW1dU=jOP
PVgkSeTECS4dlfP98UAcJ]Yj_7_c]ie5EPZLcNWE7nP:=DOhJ]HlW2<q;3K^mZ:d
m@;6JeV4Id9E5OhO4aP6aZN4>C`\L1?c4bBQbW1LEYABS^hf]2FVbDG4DB2e1XlU
2lJ5Nf;hM<BJ@a?b8a3`eO^@<Pm]MjXS;FN>imYoCEVlAJf2]bnmN=plm4KG4]Dc
`;O1U1RN:FeoR`^C5H3PX]5oPaUUagUn54kIFM>89e=b0h08@G47V4gJ;5:QYBSn
i^g9Ec?PbejFao2I55Yo2dRbOdPJ]?Z__ed93l71R;1B\>XBHMG`Pq]4S8@eiJl4
>6BDdkJL8CK`f@PIA^]ifg5WNZYa4k26;2LHCo_ZY><ZjREXj\9TSFJX_SNXX?Cj
7_kjOZ=AX2]o4^IdlPPhpK`XmA1pN;@X6h6$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR4(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
]k=9;SQH5DT^<=8bOYVP`7dIB5^V5=qV6DBOCG6^\g<WATbPZoUMP9lT?gTVQPa_
DbFBX=5E6HiVeShS[8MN2WcpA;UYL=Y>_A4MSL^<DSVMlehBW3YEXTcGHgLG>S:O
W[;b^XV>Db@JS<UgPZn?0ZUXNh=1H@UUp>h<J@>p\Va@X74gXKPbB@YFn^]0B]MS
Z[YO4=0?]WeK5>6L]S[CWCp4C?Xl\Vp=GG@O1qf@ji1jEQ`2bB@e`LKg@7PNl<GB
X<6ODQVfP;7PTd=TgCE?6:B<iLHCJHjg]FQ<jV]R:]I^F2SD=P;mT[93]3mma^?B
EG2U6GlajIU@EjPN\VYA\L2@Ul`3=57hUk93\[fRbi=:2[IAIa37p21g<eMoDaaS
a16==`:L>FXB0l?CigMe^58Pk=D8>Q\BR9L9>9DELN4laf_5FlAYK?4Y6hicZAH3
>QMn<^NDSXMlcj?Ra[J9KYTJM:=@omLOBQ]gD\\iIkMR<m@DOf^N524PR@L<HgC@
N`epVV>_ON86NVTAFL1_okX7d9E;ZnMb8I4pm4FQaBP3bj;FnO;X\^kKWShTo[mB
]fXFRVoN9nAl8QODRe141d=S7Nkj?VDF`70PFWE2jii;gg<Tb4c2W`nk<Y?RJ[\Z
a8Na]7HDiiHlc6>h;K`\UC=bmBGEnU7E`;@XmW=aU94JK7FE_AqDWhiASaUU_^cC
gQ\EjHg_Pn?kWhO;h_VQ9_7e>9OJ:;=C>3L_D_LNhdYAmo4>co_81DXHmm1b6<GZ
NF4g:j1>?gnLWRMa4E@JP`D>>AP3PGg_5K<WFY?k>Cd3f9e5k]gD1k?c]d_@?PdC
@qjMZ;@i_7?6C]m5`InOI_X`3NU[SQ3AH:US5i;MHXYc=LGH5JV@`i?6@jBhMU2X
Fo8mL;7WEfk8k43U03iim:SAlW4[W2OdF2l6Qjchcj<Q:^NahD]ON9onZ9GZ>kCE
5Ojm:;nMn<]_A`h:qecgAE]]:1L47nCNPB8:XlFTMN8;=YMVFF6a]BoI]<6P>Lme
YL<jU]JYhX;HaLGMH2bMOOmR1SX4Z2?olYM5I?iYOk8\?LXSF_[`FEn?AfCoTdkM
5Q7R6RTS7U9dKBoCoebKR[mTRKSOZf?qET6h_8ollSCk[SSkGAN>P`:68E<STU33
jo6L`jOf0aQJ2??WkVgkQo2kh\ofg6YJoYk3`T\BjkC\REVTRXBSKU`WaE?j5W:c
Z^EO?3;cTIOj24lQij117W>6o:ZX:kdPEY5hOn=KX8UCXaqnk<ULO34oEC:`Q9NX
G=cDHVNmWFo\heTWknbNA`]3B1OEeFkkf5mRE0CbgGjMZ0<EMakJj:3LZ\i>9jG>
kQa9LTdVWVcF3Ej5Y9BX?A@=8@kK2O?d0JcD8CdeLj\9d[cnM>]`YM?KeCA;9qX3
ZTKi=2Gano\8T95Ncj[XP=CoLL8m@Q?9BJLK?5P0WFdYb<@mR5Kgdj:KJN?jIY9;
lZ[hMLQ<a=:b2\2IVUDU?2f484=3qS==]TTbSDd>oWdRb4Q:QZ@\Gp?15AA_b9jh
3ZZaeo;^dg=m5^0KM7ZWXLJeA>62HQjje>OlnMHjRg3blD<m^^A6Bmc^Ec2jeRC;
<a_0XJHCnM3dDm>KM\\FR`Wi>cnH_56`jmC_7EhUh;b1bU=;FQ1^[D?^B\iTEJ:X
5jDlqPTP8NTUkdX\TVGA\63=XH[3g0SQl[K9?Hk>BOCl_a]CnTSP=o1\VG32fPZV
7OV;RI9e1Mg`KLPP6@iKH?CgQn]hXbS`fh<\e0JnDj]d>j_?^c3L2icB]KS;Z<8O
WXlUKPnOfoZ_Ko_8UhDp_ceh_oJ\Nb<;mhM`C\<G=KCQ>@2DoS\l8Go@a5\UZa4F
RcLm34ggEV0=XlNOUb:NW4Z:Oci_Z4kfjM@[dC=KhJ7cH@@5cANN<icaS1MUVo<h
V5c^74RcA`C<MB2CfK2F_4VbmnYoUC8K71pc3RG`P4D2HdH?jN3NX0eE2_FF<5hK
O``gPJ\b9F_bb;HC`T5FU;[fdMT80NDP[GHTR]LA:C8bPo<L6QLJX`:EH[oM<gRC
CdTRj;a=U?_^V=2\?Qnn_\RRNU_nU6AMlRocYPjXVPYU]@hVWqEQdeo:ag6O3ZmC
XidQoBYcR9V\abfTkg9=AGBkbJV1hAIg7biOd0_MAeXF@RA>K2I=Pll>]VBD9G@;
U58iT>WHE1O\abeoH7?NS=MO\ffjhAH_dWJehB`:O4YcefQdm2E:Njf]lUdOHJ>X
q5f`V5KQdL9gj9b><]\WKF;iGJ8J\Fl;1G7F\lSB5FH^8PZ2f<EFl3Imb:Zb:AUL
QQCblK\?d:>Z33AeEk\S]a1K6Q8NH8UPF?88iM>?BRS^Nb20C;6j]nV>7]S7dHAc
_535KPaDfK_DO]Jp?f;cWCjD^T<1GEV:ii\cJKCqQ0P>JOD=W`I9<Ra00^<`dSZ9
cInNG[f>BUlJM:Vh7fOK6oWCFBQFUZNX`JGOUN`joWK_;_ji5kafo^:l=AiQ[_dc
HIn>5913YM1VB;[20TN^n1j;4f@EMbSP<?KD\Sd0QWEDeZejE<H;Jgqoe\4fEa@:
]@JOXFnYbo5]F]Ug?5[GnRWLdI1MRX@Kih>eX]_H6GPdc]<L@Je5`>Q?@4iIH=;9
_YgT06I3id6OGYZb?]o\]B:<^dNnN:A?0<R2`VA^d2AVa:okF;WGQ^\o@<aCBL6H
GZ]XKqSE;OJgEUK1F;YZPLogWK4kO?^c:aaZ9c3K66@9eg68YTfnYW\CJK0hGaRa
Q_67R_UgR0CjgShE1gA\Qbllh^MnN\GS3KFYpFaRWC4QQa3dJi4H160Ph@8h_I4=
5bhASOI902:ViXKnTNQE;M[SIH5bPUPFd\hUKaoeU2cWVKa\[YceQaihEjC=LP4P
8QF@Ln4fjm9Z``SOEh6ah28G2la]TTl][I__aFo>P[UE0E]O>>?qGPQXUL>ObIc4
0g3E2jB\NiZ`]@bYY[1M^<L\FGQ[h7K\pa`>mN[fSmQiePg]Jj^Q2jY@A9K`930G
eRD`D^TXF[o^`oEHIhehkg]_dlPi0S67=8n@o_>XQje`XkFe\@SlT3PUkmKhYX]^
7BgXICU85nmmX7QA97ei@RFWeA8h54SaKanUm]Y[CJ1HjnCqM\^eE52bE2UJmI_o
YK6YC470TMHW`PERk52@<Ej1;>ennl_YZ4G0;aJf:<:>RQall8F[oBmP5G@h1UhE
^J\2^6ZNk2HRJgam<TTC<EYOUSfniFb>:G3h_VZ1;^>?FOiBL^h<h`SR[`p?oFI\
j_;g1WYT0>N6A8C3=mb2PZ2M2R]88hYHW6lU]6fM?X=dTR6EJbBS836o;WXlXR\3
1ZGYb5ghBV\ZjaV`WlJkPSH0TF_^k6A:eBNenk6TOFQ;2LLDYG5[SceM3Q9?XW>l
[mG3YMC:npWf;TUe0iAhO;[Ka_3hb;XA_G>J@WV\Ya@9>2\AEY?LlZ2D9fB_mlKj
Z_[aMZ<:9IZ\0We6L2F=oeh^:K64IBNfdOlJED^B0fhON0iC]2EQHEdUd9EG6=5I
e9OAWCmf3jW\i_3YY1[_fhHCp[\UP7b:IBI5QMQMN9AN>jJ_Jd`EnXH<5<[Q]XOb
<dBMZmeN;^KIm[<K^:2==C\HcJK3E0jHDJfo@j>bT5TnX0LU1I`=A6]W9^VCanV=
DoUc7BORQP51=lL=YEa87ABc:[KVQJQ2lT]SEGXpZG>jQNY<\4mmiL1Ie\@K]b84
^R3V80VFMH1dVTJAW8E^4kbGnTVO[SL65hHG@CkG`GWJK]37]GH@@e<KWSh[6MLQ
LJamnooWQ3Z7LTe5[g^C_;eFa=_Cdh:>i9jVM<]SGlFdPK;YQMp3_CbLi24<39af
m5GLW>`_UbJ^_O6L65`A:_kEUTWDig1<lb548;m`T3XG@UDTX?@iQlYSf8Z>jIRA
OY\n7g`:HmW^_e]a^ld^_g3O2l]Cb5185hoY>N<b=9>3X>BRPSF3Qjl95>C>I30^
dqGJ`JS=RIdEkY^Q=8LGg?3_Fk8Na4CneB1Ff7Gi0l3B6\Q2=X;O;449^m@WQS2C
G5Tg2oMPXH6YZS30>J5MNW7:ACkYJ;Phq3\LED1n3UmS?]WM`KjLM49;jfLQ16LM
NW@PgEBMHM673UWl0YHL9DQk:1EmfTof^5WK=C7:eTNF]T:k[[WfSFQC8NLG0DK<
XOX8[VQW1jd<^5`iedm\JKddd402jcSV?3Y=F<3T0bAF2@ApIX\DPGNi[V^Od]aC
SiU5bJ\hILXdN3O7BH2CKMQ52PlR7;LnM343l@E;PFT8HfD]oN0qiXVfWV^7D2H3
bH0aK@kAd=UK`gT=WhcA;@;T6gFIQ6Tme^C:OeB<3b]\D`cEGWZE2AU[_ES29[B[
2b`Hl:o85\knNgn_gA[\PWkh>jGmd6_Wl1Sb<mlhC0`G53ke7KkfiZ6`DJMd;_^2
;7qO^oaZe_2`gdVL6S`FbcQZa8e<4gMNM?K]_Gb_ijRkRa@]?^o::YZQnOh>WA4<
>CiG8Cn`DNA<RE9OBU<5o2g\A^WK4a@W^g3Cn_HY>kiK=aj`d;GUISX>V:3g@EH8
[R8Od4K@_nCXjLniYqhZNdGddD_i;5Q<?<gZ;b4TK5FH3OiL?fK65n\?cRM>B6Fk
8S1]`4en;UYHQa5j_@9_C?7DJ5nU_3dBQ22efSK9BPRH5C@STH]M]e_NWX?>Jm0^
G]YWWF6jJY:eKhMD:_h<FAkimhoFZ\jcq9<:6QiO9cG^:6FH=LkAZ;<C?YGgo8V2
pm0?IjnO_a_6<IFF;Zjka<J:Xj2MPDMcoalKZJaL\4AhV;=K2V5B044=<i6FilGB
iQeQOaHE7FoNVfOC0L^mQnJ7WM2gP3g8gb_3>XCT\?>BQPfUhg^DR27`6[9I:KR6
jm0b0T@Of<6\f2=q8UnAV_4Bg3^3m0W2jJ9`n0Z1`aWD5HmcWe\EMfYg`N^mgZjX
mM5O_?`DT1o>kmKoZeFA_QPB>7ja\SLal0?AECGNKa8AX8m:^;3P29XOKElWahWm
Z7TJh208HBRkZK]h8RH][6i=B:MA5cq8lF>BND6=ehoQ`[UAmOnEa8SWUn6Sga0=
d<=OIF<INVkeoWf`\ePXVQ33=YZmE=F:]DMcWbV;D>EFj8G0m9^1GKR3UVP`KdZ5
5>`fG4GJDio<]Do^Nco<Mj`M_NeeYO883bHncMM[2]TMMp[ClRP1RP83f2>5333a
p^:PY:KdZl9fV_2W8dh\Dh9=KID3M99@_O2B=M=obGKjl6@Ag;?RhQN;Vh1OAQ4j
?6H2oD;aEROk=;?5FRTG\D[FhiDAL2NJ5G`kZeE_5l@@H>5@U9a_9O0c>]G8?dlc
C^hc_[JI=HF:c=dq1<_R:b8ig8<P1KS91cdg@@VYTd>l@SJbKT9:fM<_PLBdV;:E
PgUJOl0ojc=P2MVWK<18b0kjfUco^Gh?h<C@eaI2>?IbA<q4F5aR`q8F]JT_V$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR4P(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
8=e?gSQd5DT^<2g`j9`:6H<<2W0H7>AkV[J;IdP5LfZqSVlmXoid\Z982@M3Ic@`
FWo8X`hYRGDICeo[N4hTJbT4nc9Oa3Y]5:X6qf;P8Mh9>W[k6n[_=eQTID4Id`Hc
m8iQT3L[7VHMeOU797fJV]3J?T_\he1\m2NGE<G\q\Jfh_MqWlncNLWh24aMRY2=
jQdkEYdU_bU36R=fbiGFG?6PMDE0ooq`@62Y6\pcHRS2_oDO\>dn_SPbdq991I64
q;<=Bic6NMYUh_>PFD46@kW9JW>dhLTM8]I[>^8F0\R6YnR`ZdSm;1[lVc=Z5mbE
L_AeWk_DfDk__hb52_j;6gTMNL>9DJ5L0anG[2K4[6ng^hg8SHj[7eC=U7l`KASJ
Q;AAjchHAJ<l@_kq`0G6nijA:mY7P\cFX^Eb\X55YKQcYBlaklJ:n<ADcXk4K;E4
n0UABQil\m<E3ihNh5di>?:me;kE?KUY\Y1:HZPUAKH8XH\f4^fESjXU3:_b0d;A
Na[KOl<cAT8kkcCZ`5mn_dWLa5ncnXpG?GG5cHmEJV@XI5P_0`[oBeGa9aF8`e?J
\]34cdf_7X@QgdmUdnR5DaF7C4_]GhBAQf:odL0NMgIl;U4l0mBZAU7h9PiZSiWZ
9a==P4oS4SiK=V?OOD[ZIjA:AOE_5fJGQ[Pg=NDhi>dL0qWNUB9EoDn1:?6T77L0
3n4e6LAF@;L@]VaTdb_HY<PC2ZDjQoM2R3[K0KeAAKGH9N@aU4IEIacc52Q:0h8K
81A>^`0F@;^Q[hkET:NG5=Og0>3iI_AbRO9Snl98kWK^14WaHBcf;gif=liNp:O2
=K0Nj]2Jnkg:k=Cm;NYG3>2If27CRDP^NPU;G\<@WOk1C=jL5Kj9\E:hIl:<PZKi
V2;C;FZWW_kVdVlH\62HXg2Ii;F0c4A6:dT`d^YQ9<:6dC27M<PDd3_6cLdb>:KL
8=gJ^\gojH1pO^D>m=m\T41JmKf;CPhZHUoUW=ATni\9_H5cflHhL:MOk`dSU5S<
VABSqN2R><=iKA:d@f;Q;OmeF[M6LNJb_ISZngY`GJ[0B^TY^RDYe2gfJaWC?[8F
>_5B2^MoF6ET@I[`mKl\ihHM5N<?[:JbKdWIETW4<:mD3YGE<G2\Q>c_m]H_c;F:
b6TMANML^>cebRWU^idp?PHG`nH[lPWVk\m2O8:l=TEH1hKjBn0cMA7ZhQcS`WX1
8dhgI4m6fFdLU65DU3b`ZK;;k^kiZ2]f2Vk4ZEUcH0oNdh9:Fe7`n8D6Hcm;UEi9
M@O_Ue_?KPL=nBid`6[V?KB8BmcanimBcYqA<>c><?5TGc4XBh\C3mcWe]IjcE4X
<UCfYoo>];K9LP5DN`ERn\8C66=En?dWhDAmmHVjdLKi07dM^L`@SghTVC[Cc6En
IF?BZ[B7`TKQNN_Ea=N32i<k5iX6a9Oj<@6AmkjfYfG\KoA`Kp7nn@OgNZG[:23f
6[_]i6b;NY97LLDk>UNQK7f9QKLUBY07hPdnPf\MR<mDZkjC1bP^BRZ2?TSfcc>m
cmd2`8F2;Wf8KRUApE@9oJcV@GBG9M[IaH\V_<>\hQG>hBg2[f8oGXMJ\omYXBXb
jD]G287ik_Lb[]37kYHB;^Nb\JA>5d0`DF;fc>9]haGHaY;58?LUH_>mnk<^Mm^R
:j?76\R^NOh:`g<O@Ee<1]@Zd_IUZG8q^o<lU_2>`m\PJ_TTKBgG7B]HIiA5dhK9
Tbd]9=7@Ae1M<?L3o@`kJlIQ]mO]lZ@m83[ea`6Zm[\j3DaflB\^c_:aAiMFT_mM
=4UHJ7MW8c1GTJlWf@1ogJjE?a1n_QV<^FVdEE:8\@R\c`p1C_JJKGBQY5SIXVnB
YCPV97gkc57HCnioceLeDR_^`7IQ^]><dDUYim?ZNfQAd^0[<HAT^Eo7>NZR;BNL
SfQ>L;`dc2^M<GDID4<_ZPBUE2L:`\om[mAOkkdUWQJGQl[1<`YRcbn5CQ95`qPk
ZoG1<hg539E^jDgE\WL0bJcFECl]7N=PXihITA=4Y]a\nXYR;nY8[6jW=pgmU?YD
<@;;kMjXC;WRoUjRRjjF7_l11<HR5E_fJIm`^MZ2njOac@akB76fKM_5Tj[C2>i4
8De=FoW=ZTdC2LJ2Db\FKMb@EI=KV9E;J7nUj2\b:C^hYDInV8h4GDUSUlgd[cBn
AKAKRj:EpRP^<>M0WajdK<\jXk2=RP<26TcMYoScC1Dd:_T=@5\J1EdiZ`imJgTN
MnROoI8MVM2c[4?aX?7fgGf3k;<d@^kG^IcMYaY8jGj9T=EVe<o:<aBXNQig?a8?
]R0lACRE0R14\TmglWNlXRMqIR\SaPE?\G;_U<R2e[AJ4R`5m992M<aF^?K`dmWT
Mh:7cYW@Z>nDEPMF<ge:K_:]4Qj`>0SBDM;H4>\C3<`<9<1^T9F4ngM^?mCBZ_Fb
]igglA9c\`899Ca9nfFA=K`UI9eMC:gOCL7OYdpIhgES;b@S7R?lbeYIX=k\=;Ni
NIIgU`T5T5m00klh9ER\fCTb]EcY>31XcZ1:LQ14XHX6IadV2O71FTfinD7YDd2i
N9[WnaiHXUCYBb2^c[?Adb3Y]No2miJb_OI;>jUIaoVa]^PXl:937pg1j6K7]Rkj
5VAncVm\9fCUQ4M9\ZMUVAHZZ5K9>o=:?=2DoHBdqm8=Ce6TbU<^R\k5oF:AYZf`
oPU`PMQGV^0S4Bg8?5?4R`_@TY=hh_MdABYHb>ko_?f_mB;m2gC@VDm`F@4XFe5C
bJUWc>\PlE\MliP5Kk027V\Jg[;MDA;8U975273kAmf9=[CDiY4hc=\qc@OnJSg0
2A5Wg3d2fXIGJ=?0chhO<2>L;\B@n<8\gID\5I8NJmYCfHI5@XW=DG_X@kOFkEM@
lSg2@D:5H:]NB\1Q9H1kZ[qG?R^G9T9nDYFO2L:WAobXV]75^he8l=<PdCGjn]ck
]K4HTMg=emdNM_;Kd>YK2J\B15HocjV3Kk]c?gTd]TBNVVWE^SEDc\GdFB;`BM_\
8Knnen>;LYY[;@DRiaWF:7HG1?nlA67FX:Q1QqLR1Hm;?Bb=4Ned\b4Hgg4PF`77
c3oBdlc@^[8S:cGcD4RWPU;lX2oLe@3I>`mKABlSO1`;UE[9\^H@:?J4=a]Y1RX7
O3VF76>GegooR=>57Va?[FUfb@C8`PO81;`NOILS^>ZQ5\^l_LWXpFNP>920J[>a
]`4O4FOj^NLKLWL^Q2S6D2LaPNSZ7UUChZCLG=lQ16Q8HklcYYJXeI`O7<N>_1hO
Pl=STdGnAGU6?bL;h:o@kdJ`l^6OXJ]CJlI5=1e@3^6EKSA4@Y>:kF`8:]kM5gDK
^0Dqi<]:TPUHYc@<;]Nd;nN;@\fjE5TE1`FHH]@A?[[5fd4bTT>kKm[S7oMMN;k6
6;6Fam]>^0O?D45E9H32Ca[`\P0Xk5PbmnZA\jC<<j_O=iW0@E8@8N7R@jcbg1nE
Vbb>imS3fHhi^k0P5]pFT^3XXj9^LW@]5:h\8S_PL6YKYTLV0lGQ0mM]m=fPnKan
WMCMgjUZf`]@IjU4\23:PVK>H;N4eMj8YfCek4QlWC\2YBNoUEA^`VDI^b:SW6eX
9V>:oSo<\NdRj0fe9^AFPQ_b4E]k1OYhepc77NAVVe3C2<S9H9Y6N<M[KA;]@YUA
NVmAALbIGa1JX>b0H]3eMa[W8fIRkhJBn\:@WHC^[BA7lKCB==<L18Fe?ZM]8Dfa
giN<7MamcVHS;`o=E9AD8=<Dm>?^_753C2c@0VS6Pj?l2l@IpcA@j@\7QZM?T_dj
W?OOiBEjnLhNgLT\A<]`NhboKIKN9LCNU8]8S9NRD<QqhMe_dKKeYQ44l^TJP:MM
GQT;b?Bbnnaibl_?nCaC:l;XFZG7Y>UI=cATFV\6nDT:=W2DP^TE\[nmPmfbN^4C
L0Ak??_PKT7WEVXZH=bbG>Uda8AOOn5CRfW:^HlEJ?;RhWbf@8SeB>DldbpADGJP
3dkcmVeIo]fZ_[PE@ZK[M5BdZk\UfjaQOXeNCg?6]Age[NfF\TeRN@QXl=7iM;al
`mShOY]VhLMPFL84;Vh9MYUEhWeH??R;3RBjc7QUOCU[^WTW`M@e>Pnl7^>AM\g\
Hf@C:FbkdqY;HSDT8ehFAHbDFDTKIJ6hg1=CR?Igc<ejNI0M<a@TS^KeInPB[aG7
LGdO8h33kmg2ab_MC3V^5TUS;SYFC2JaUb8SWB?WqGMP8MeCV1oV[3]QAL?0DYo=
chf@HIMinjmSZOGDoiW0V`ai3:KBMlofg_2W8d_\W:9=Pom>M62U]iZZ@VW2fX76
6Df7Mo[W9AB2UW3TjZe1daZl_QK2ZTF=7n]S33i][GKf1h7m`jN?RX6p>C8]d>3]
Ofn4mUHlZBflkncEg=cWLlBYC^jaa=o7COLjiC06M3YogZJmMdW4O[WmhARc2=AO
<G[2nd3m1V50JBehP=Q=bn6RUXoL[L^_]aR5G>Ffn`f=3^_SOeAC05F_>=M[VeD1
3jE:>Wp`;1\fbK<=n28OY^:]Q@Z=eCRVB85N:gf5@gagMIF0geaF9GFG8WI:8Kh<
NO8QRh81JUZf]L^61RHKF2AOejAj?OmZBS6V\@m<=GRPdVAeh0101Q:ghm1^n3V1
12A03;a`mNhmYB6^heZX5p2C__iF6;jCfJ^W7fPG]^gDek6E]@R<nTAW5lf>4Woc
LiOTW=e;;o2Cm7LTgHoZANfmL[7X<S?L2n8E_gF:8W8dUG3E=oei55O]JgYOB=BC
\5YU?T7gXfD@2F=b_P]5\P2_;FX_@_CV6ZL1p=g<]gQoBV@QT0<mlLVPi9IF7o26
TaDAKbccP^6:?8HNG2bQ4d2II^\8_9S98ffRY;cbGRMjFOob`0o0e3KdIoLWVg2o
anEF@R]:Qik7C<2HX=TVE1`H\S4^=B7]1K^8B=EeK5Gl^DI]Nm;pFI;mJ8:i]]\a
Pk2W]S:J<6?[ffA04X9CJM4Y<eR]92@;mTSS>kZ[fV?elkh_eN\1d=7b?6Q`UCKX
R;ViRDCLlIk6XfA_T7PAh_^UkkSB3FNI\X24Q5fk4JP]3@E<1JI7F]FX_[[k`CBY
2opc`jJX=\kA@e`>`opD^Bjn69l@Z]1;iFjA^[FKQH2D4SKGN<kBAmNOnjUPQNAB
No@1`PDd1>o?4`C9=JS1bl_jjc=];OSVSkK:??b0OW0b4I^>88lYd__]GGh<9gQj
;`lM\fX1SUEZ1?NK^8jDVUe;\hodKDJP`q39\]j?Ol=C_L<oSU:PMoJC@T4<Rnoj
VT5<COZQM^D`]h=E3MH6FJPeMAFG;0@i4We;2<0_J9EUQWC2gL@A\2JUWiK<G5?l
2DiB@F_>`^]mEbg?Aai6O83bhSB=0VE48:3D1YQ6Z2[af<CRq0LL5Vd;72fZW2\1
YW90h364HRZj:eG6l`MUcLG6ON\M>d3d4bn;Fj2^eIO0Q37GkQ37J3ko_Cj2TB9@
N4;\0=QBnUm0RLmqNT>YBGpJn=@0IG$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR4S(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
P]NgVSQd5DT^<CdY^FV<<hkVa5FCG757Ff1ECU3H73m6ARl_We<f40F=qQV<cUO4
Rj8UXnMpdL:YnJIE@1m:WPmXDG^C4JQ6[AAY[@@mfPIIC3D9;`H7haa34:bN7D6X
GW1q9A`jD=pMOEfibLTI`fkk6@o\je=aJ\YfemH?eGfjBNgX^cVnjE`3Wpcj_k?Z
`p@^HLEXqNkh9]8^VZ8Yo`7Kf1YI737Na:g\hWeT797kI=\A1E2P<Hn?SQliR\_l
`]Go`?;6[IgmYE\Nm1^jTe=4682OiB4?;IgY]cF5nE36>l2X89[bV]6b[Z1^jb]C
_cA:h1nkSNg@aS^8WfREdAPpmf2VOBV1fc7T[\;H:adAi=9KMKoiJXO\[ed[kHUQ
\e<^lJ0KDH7e0R@8:OSVThk?FkLBT@U@he?8H9LfPamD>U1A[K7k9`>J3\OPTD\g
6lk1XF3fVJnek7VZF@6n\b=Jmk@?@l0OQJGlXQq_HXll4Ka9KhQQdS;0I_=h5o2J
\klA25G6C9cKCA04<If<E6DF@?\5XK8liSaZ8JKknVU?VedoAjibfNQfJLRJCbjL
\P<@l32OlhD4Hg6g<GMLGknD\C5G@:l\H2PbMm3_nV\jDkk[32PeSqll4g6SeO\h
`kN:dcW4mVNR7a>^NJY0kf[_m0flYmDjR7]oF9j>5k^AU;JGLGjiL:Z56DFDG1Ho
1aBcBi1]EDIB=T>^<5Y89b9TmaXG76KlT?]JM5MBL2M2Aac9WONEUDl5@3@kKgi=
0LM>q6ko2`M>KU@54o<>9N\[>`ZW]miO[XnM@Cd<0U`Hf:=K2?N_MUDonXTD]62p
5Ud=jLC5a=gWV_J`8^::L2ll[7G[B5[h7nf00LJJGW]\Z^oQ]AZkJFYOe6<A\5Pj
PSWAMSaoPBUQ^PJWmlF3>lQhi7J8KPHGZ7K1]QXHGl2aYV19hAgiCeAXZA[CC5ji
5S>CTPYeR5Bc8BpO@`P2iUIDNIaZj;m^WN`0L@dTkTA342[Q1F\cmK23MMomKIH5
gK_:]8VmISJd7T:3^TbNMgTd=B`Z[:\^YH8BW^:<k49T@Yg<aQYl5IMlC06_5GIo
Z`YmnCDcP7N7i;]O^OK5fDb?b`8Z>qBkP6dO?N@4]_BFL<]=;A2iBiY6<EOY7X1H
`AF[OAG>7^QWKP@i;cT;AX\NI2C5:>`]Fi?GoBZomR63JR9[U8UPL_662UEbV2N[
nYm:iOm96?[EZf<3dMa=?b?1aDH=LhB]K_fM:`Ld@AR2ql1C\5Q90XEfXGIRcMC;
7fg;nTa6N7hdD3?7G=8k3CPMNJ;Y=9Ej>nK:T6T77LK3O9e6MP4c7[73ISdTJAO:
g85MnXa;J4idiM4@L0jOik6PnQ7L:GF1DSf9igNWnU<fOleD\3Y@<GQW7gCq46HW
WE9Re>;I^f3R=mSfobLB8iJ=>V?:m5MFn7\GDGX[O2\b4_H@MiZo7olnXQm=;[^d
gHXR;<^o8_@mc>:IT:9TjbZVG_qn?PB=MTGHWK4Ola=gRdi]7L:ZEOCZjV3mohSQ
6VDKhWk=kU<\a\2be1gI@m5JO358f>\M?\;Sh[bhaZhWHn0PZ[ESEk=G^]eOe@=>
X7[IZ8DdmN0i2mj0dC0`:oR<l<OnfO`U0>9GZ0WI=q[L[f0maOh\R0GJUAS2[<B>
9Q7K49WG9`lS\B@SWama\Uf;j:]Eh[RAP;;ZB_ocab8F7=Hn_NUcG_^g`XW_0M>e
F\\K1WHjN9fjn@^iiPFkQd[IM[D4GGj>F7>4>2e_Y2[FYfeb@IMW?SWBpm:5dPXh
^7\H?RH9YV7<SU\hn8D6=\M`P<SG;IhMfV[ST375;jmTeNahRkJk8d^R?a7lNOBi
9mXT63VCl:f?8V4cTYD6g?lT90eMe]_i`0jOVHXTP_k_71P3oLeR:479`m7hBFPh
W5?HUiLqAZCiiS5Vjg4J6[C@9Ejc<KcQ?ejcESRO_1;[q:klTQMS`cSJ_05fO;X[
F1C7lG5foOiXL86;O><AUlT>N;Xb@;Bl^k14ChN7e;mQ@O?h5lfa08_>05YUj`cj
VQN:_i50i]@aa=1iKkIe548T\kQFkO9Lm8FnO?00DjPhN:?nhdJe7`:_8FnqSmQ9
hSAM8Ij;HUc=HGnB4791@XIUFAc1Rbf14Al1Pc1XdeUQ6J>kg?@gUk43=biaA<UW
Vjc1RX`8\FmV>67JA2Vf>XYNiYZ3P`10H9[?2PeK>7[5N_FhJ1jgO:cNX83DS<SO
m2QOL0k@VEp3;X7X7dMl91_ncAZdHYLmAElk1dRl5h8RcdVe7?RmV;d3>\8Qbl\X
6ORPj33Gbm8]^QdM>[[CE]k4=dZW5WMUY<3018V@9lSee7:MD]k2la=2S`oST;[a
`iln3nA@G<o3^gBI_Y1[Dg53]pgh62iiN_Z?fP\EhJFj=N>aOReIT1kOA46P`d6T
EkfnQQB`Qd:9AA`nil>V`4360OOW\h2kg;R_oO?Y5SX^7=4TieEICiaSQ8^b2OZQ
S\I0M]HnJ?C?>5jd967KAb9ZH7gWl[UlYk80j19bpCe8:SLggG\FYC:U>E?X:93J
[cYD6N?D7K5^eFi[<1K0kl0PXlRY^\AWcY2TVFQ^BjL=?k4C[cKG=d0d_leXJ?MF
SPYD6^9]FZH=Xjll5jP87moTKH_YJ>\M5a<K;5\EXCLd?lBFKX@beQdqkOV]C_CH
2M<iH^iWBl<Z]4J5Ld>S2\<:E1W5X`0g`_QMMjg794\:LCWGSV^7<[]lU0RibTAW
8:0oEIK[f19i02TbBSBB?9pJCS2D=5MKIW\VE4iX?X^;dmKc1K81hpP:gn2eDWZX
J8LFjL2;2hDU700OKS\A<KY<m=cKOdl=XXY>mM?SV<do_JhmQ3o<UFAC^Q03_P5=
TKRcRUf03WoZ;GNOKO<XfE]_><Co0^6=@i;D`amSACl_ib20S@@WGoPC1Go`i:Ne
RN^1p6HCSo01dm8_O[YQ^X_L1TE7=_;fN]@f[6e?MjU6W8\k3?44CS2n:NPU3ZXQ
7^W0b?L2j<]1G\`GXZ_P4YB;\SU?4jfHR\g\K6dZ`KRN_^]@emFiB_`WGf?_CTT;
JJWWHhUPkik4B@BpF2_nL<nD@^170e@Mf^N@k4`N8?4S62L:ebVoUF0XaH`KW=2U
=BAdLYgVXk@V55=k]Hm^5\bA3D1chkAdbKnO<TbI8>W\8EVn]LXWFFoW^S=ZL3DN
AQA][BBZdZM;TKimAi]9g4h7ecp6IYcYcnRD2o8<==g?6X5=mM5XRKb?bpOBZOPT
;7]NTgQ[6a98c3mIkDH;9oLAoneihaYMZX_d6gX;Ui`1=6bTAFB`BZH_6H=XEcC4
:Kb8EVfF?;P8;;Jb9W_;SGGLfme_;?mPIe_@48JLELaIE=f;_@kdi\6_`=OX3eFd
EXdc8ohjpOK:OF9i6U:NX`JGO;8`?1WK_fF:FTk?[9M1`8d`;3^5B8U4OfWbWEjI
7N5@\W9@QBoWLi4Q`VXmQU9AdJ8POGk^V^F:oU<G9X4CHDe51^fgM^B__H2fSO[H
AL:<U7dW0OoT^6cM\BbUST?q0NiBPWcDb7DHK12`^_PDKhP]NfVbYZN6<A=B?ESL
I?S<=JWKe`?o[P]oKPPWnZ\CUP2PL57I;mS7de0UJjE6NYjOdCoTUCJOeG_>6n^b
XNX3lm_43733QGXj5;mUYZ=Nm;PL?GfNg9qAD54QC8OU_NK\9@n9`06[n1gh]PTB
\`KinFYEDm8K9Hh3]QAi70k]d6Ee5cioUOAc0ND]ko18lAE^hc_[JI=4Cf2g?=ER
hGgDk>DND0\2NJ5GnkZeE_5l@@H>5@U9>_9O>SR`3M>72pD83Rlakej2eToF^HF9
^:1UQQGL8BdL3H567]=dOfUI^GN?;9hhVC29@P\\<JA]a3THQm=S^lSR\fBU89`S
c?A=FOPLQ1kddN>nd<MK17=A<9\17HHh2CD=BC9bnL`dbYDHid80TaBD]Rcbq[Pf
T2:mQ5mT6jgNhFY<XbA12GGGJ2Im7JI:F3E1hbYM21:6FQ5[YV68RJ7VDPC6^@7=
c@T5G>M?5<aM<Z_4eOmE<fJSjI=qod@Wb>U?:<Kab;=Y?0JcKjg=n4mYXBGbBbLl
W8cAGgV1a;ialEh>KELkfRb;GU23N0dF>BBZ<XY0ajMQUb[90d0Sk4mYSU3V@H9\
mY231Q>dLem7dRU:WO`0lNZO1Tf\oVdWJ`m1hQfVOkqL;9doPVQLF2k6hWIbbjn0
fJnD3Wla3VdKS33kmoEE\L@>SUMKeOGYZ1ZgB0QB@<PNQbI?=WEmUCVdj0GcYORM
0b^S3obZ1I=aW6kEanY4;G?U`WIe1:od:O]>SgEB1eKL1hG>KL?N3FR]DpRP]<\T
Xf8CageFRZJ[9`DCY?@F]AJR=J?YMJEBMKcISg4UIUZ`:^eA@mL3[_9k7kOmqdQY
0>Za>LNYce>RL<FgnAoD3FQd@<m3a8k5d:j_?\7TedOg>??:`]W3>haJ`A:>2c6<
h?BhZdjV6[C^WckSQH3@dAQd`CZiK>UIIXB;@h4Ho5;CVb50DkH;Gej]nb]b3ded
kZS`g\15@ioq_\=14Pa?K33ijnPMbQS_2G8P]4M;KO`D[oB^OEG96f\Ao6cgCUA@
6m?R4fPX]6RfHVMNiYnAX?:B]iVZ?_:[a[Na74R^:M]RgmIlGC1Tbnk27_?\bEEQ
Id\PhBFWQXlF_b\jTdkNnXjC;2pShWYFa63jJUPQOjCOcOo3HWcZM_SLV\0]d<MU
E`[H:9d<QNdN1n]SCHOH4eXQl0\TG<MIM0@DKPnfj=fjeKhQn=61M=oi553gTk<1
AReD?FcD8;V_DaTWcCPM03@_\Z:S^D4Q[_4gUDn5mpm]k<fNlR:LBShU]jA7[:79
WDYoSW^P<1ekaC8WT5Z\?TG^O5`L3fgM\ITm?iOWY?<UI71n?R`]KE@5G73=lL<D
R3BoTiP]:WUECm@YXAZAjH\HcOCFnLcZZ:Og8dXWRMm7ZVDWePXD=^m1p2SZ<5nl
9b`T_ffkAB\JDKh^]lil<C\<ER?NGLWkYeDf[LT[9BA5BC>ef\0Wc:Ufi_hLi6Sc
1QVUQSB]5KHFRnnd0liMl20j?:<UCOEAS<Rf=HBZgLBKlcn3C_^JY[akO2:g_>jG
;McT0\mqkZE2:QSf18@a<oioh=KgS5iM9Z6l0JbD`WW8[Ta>IB\NQ>4hWINhZN^W
TQJVgHJ5H5Y:h5;=[H[lS_;<LPX\^\ZB3Z\l=2`kb]_P4[UE1oOiTfk0ScC_k8=h
9h``fn;<kkVUAn0`XgOEKjpk[]H@o=igo^BnE32GIL=]KAdfKNM\\]3^cId[8RC=
44\R>@miiYVCm\1S7JLK0_n?jQGQ[ZMYg]DUPZ]oRP[1gG:[]JXKepImPDKeqnfL
P?ZbIO<5nP6ile^6fO2DphQ_5Zn^$
`endprotected
endmodule
`endcelldefine


//-- FTC standard cell revision 1.1 --//
`resetall
`timescale 10ps/1ps
`celldefine
module XOR4T(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;

//Function Block
`protected
fNnkVSQV5DT^<ZCXKl>=]CJ@Y[ndb1lQCbT\i;lbfGY[jfRk8X>kAXCZgJDG336@
WfNEI3epRgbMh9j9Y5B^KFB?5CEYTFMqj:mfAOZ>i12``BR=5ULfBBhh2mj1bVWm
cNlUndA=i4<>phFCED=pD649KB_QAE1;<]3a[aZn`H5Vca:1m1>9E>3lBYObP6Y=
ZWqX_gQZf\qnBP^YmqkgJZVo`FeK`Cc8iO96Vd]E5iO3G_`08kVHH<b47hkM[5]7
o79OjIS<0f0;gGMnGCL]6;OcRChhBWbHLIFmMU=53<C3GYDhO:cm66P:Z[]J[AiO
]PJdRL94UA7W?cT;PYk<c9B^WhWo<O<cp13QD3TZgNRPbXlT?Do=9HCfNU9Q35^j
]UR[WmZ@afFV4Nk:D>4ST`MN2IZeZiAEV\T^Z>:^[\UhQU[<9^I5D<GkdI9Q3=:n
^NN5Xfk;FMShQES;]gMPKfU<a@a??4foS1YXZo_A^=L3a2iqc@]kI\4daRdJ1e:c
DQZ4N0JV6HV]I8YD`MD;10oUG;PXidW:[>ceBNjcjTDao?m:Hf]^OEGS5\HRd611
aQWmge_T>H8]YO[oF34PXB4IF<a1;_dkM\c;SnUAQaTXj>0Qcfhkm4a^?;2bElpj
RN8cZhTUG]DbC\DOP5ji4<N^OJLA;_OkcNIfXgB=k42G_ab8TYZYCZE:j;`o:EPK
RbIjPVL]5SQXN6aV^l>UT]6ZO[EEYKnkfhG6@QB[jW9Lb_joW[JY2<e]3dH2ceOj
HOS;m@AS7:ZU=p9TNX2YVTG0HS7C102:?d:Q7kHFaHhNjiUdc5;=IX<G:4kNO4lF
^VIho[J4PV9WKjQEoiHFkG`B7`3g>NGL8UIlNfbF3[@obPMX:\cg^<ib80nELeJj
AgM7B\QSF:hjYc9FkHg4DS[:5EYQqOYR9^Y1FaWISi@EjmgX1P@Q<P9V6P[55`:Y
ocfNn4hS8Oi`oYX[eWl2ZR`m\q47iR_fQ;_d3ShkO7JeJ^?4BVLCXmlZ3>Ph560l
1EhhelZ95G_@KUad7\C3l9TX\m6InGT^Mn^P[LREilMCWb0j5FRC7g[lPI;4KUoo
]UENelGc8WkB@]oO8[TFZD;dB<4f@fGJGHcCSJkOpi:gmc8V]WfRA;_\LTQK5gGn
jZoJ>lT9G`=;:4HJL9?oV=@_Fa:;]l4UYKQ1mHZD<SO73DN[21mBT^5W;_OYDlOV
WOoKVbF:@P=\@0lb0609ZV]g0R`=EfDA0?8Z_<^GjiO[mN7QVOVFD_`qlWT;RR^\
gmKBMKE@3F9do=Y1k3h?l2mDF^2IElA>04cF\F9Ff`UP>R\FWoH=^IV9HgL\Uc90
Lf[S0WD=5NSi2<ENF3h]7K`E8b<]eS15cIGUYe:T_=oLGZ3lnB5VYFi5lYl6QMIH
DZT0Xhpl_3JGKKQ[j3jCiY9>3lAOnVGZbTT:6Afe[KTHON<_J[k54Yk\=mheF=]<
6k3`eKa6ND0=2Vi@gkWa<dcnBmo:W3ZN22X>0qj4UmDnF_fL6[X]LA10H4F`?Ug4
i]kBl[3QT5P;k]FLPNhK3=7aWNoal6A@K5c6CkH<>mE=D^CUcFgV8b;;AYldG@34
i]e9cUlV^RHLha=Jcc@M=X]oWeZlBf2blJ>E1njT^TcGW7aB;g@opYP<Y;RIO9fM
:FPK`ZODDUOakL]_?j@YdmEb71J=U@7B=RTFb?`S=`SM^aohAK?X_Wjj><[YEeDS
?mPY1[jQ^99?WE]Jch1`0NjY<k@5_62\KS]AD[`?K^3lSePiIHJGeYkH:fiK6S]e
<7oq0RfejOV3XYPUllkM\dfmE@KXQZ2dhOH3SU4>VEWOU25bWMX:BaKlMT:3CC8f
7fN9JgbDi4k7GI59akDfd1<O5L?<]ZH?LNFena7jHK?PB?^oCJn3c3RneM`H`=\6
fB>f0g8GocleM^caVkq\DiSa8]WiFo:9AioD=qdPgUNl<@60IJWDH@3V?Hc8ROGS
T?86KSLC[KBFnR8?B5D=b`9=G:l@7AaC\D3bDBQ=`85mhAZUVm2[;TI]>mVdoa1S
XURRAjc20B<SWHil9g]8MQ37bXMmT\@7R_]ZK;d08A=UYnNLL<Yiq93hjH>1HEZb
:gJMj_19aaikOZhN4i@O?ISVJ<OlADQ7Q^BmBTNP`T4ODNQjG0cE79UWIg@OFZPd
_Te\T<272ni>BhhXDCdYkBndhCZja[EU1b0F[d0nn6EKH4doY4DR09Koa>MU:g^T
lm:pcgcDMk6GFGYgLN[m9bFRc0[1lmCDhMZUY\IC9>=;jS<cbWh>0VPVLejInG`:
SX1If0[;XT^dLgELji\9n\I5:==Q=mbW75VRlaj3m<WYNE:DYIE>^VM@WBM40O=U
9j=@c<WaK?KoL_Ffk6pM`m>RTH5I?]bPb[j[UF=MG:FMXREaWXdk`4WZEWN_VNU[
Dh6;\@?_ANnbZ2CQeTnPeoFn8jWe1Rin]=H]dfAfeRoWXR1N3kZ2:0bUCA1@<TJE
jCcK<WM=To>GcMJiULhMBQ>LKG_cUPXICq6We09OUQ87kEePjEDHAJ2aW[?Id@5Z
:DB;Y:LAmOmofRdVaW<jUanbBkiZFmCcl[U;MYEBGUI86F5a51CHCQb6n]hIL7L^
?;?KRFUIcdN6QSQjlIl\B@aRaY:PII11Y76;^mB@nfD[mgk^pOVBAnlmn4LkcnEl
oClKeaBhBYSnoF4^MBVFa?hF2PD6NHUTjS=UTW:NO8`m2KGFUhR^Vh[[PYhMRBk8
[bleQ?4X\4;BCH>qS_[>Lh2iNl@:NHR2RT:aPPL56CMZo;B[`dX^F;jnOfO_0I<k
J>qHZSN0ho7D9o`C>C2GE^<=O`neHhA>eEca;5C:VDGo2T0UQ>WE4HJn7WUZ?<Th
Oo6kneCZ=7GT3X40lZSnKbQ7QQ6nHAf;Q:eEDjEY=[Zj`Y@acmbbYE;?lYb0SDS0
oVlHn:g27UE80BI[6pF[<Y<Whbb>R7MLf1044g^XMA0ObNBAE:\oWW[`hcgFRgi\
@R^M?AAg1YD1Ui0f9lVBE[@G7_0_P9Lc7lb40LOUTcUOM;nK9;iid@V@7QEc>a4W
8;_<9H<g^\<37l^OWNFBijO>2l2>:UilpE<_J17Z@2AQ4>K_Da@lJ:^EVaRAH1YP
`kQ]b<MYQ?H:JPA0b6Q3P726X12?EnD49KIjo8gKkIDb:IgDQ6X48_[_obR\SmOO
6E9iUWSJLR3^JLf_0=R;Tl<C3XYBmDJ>6EILV>`6XL29@@DqLMLXVBPiEi3P6@ln
_8dRjBdb6aFC`MgFP@Z[<LZ12WfnMgf=?UZ8k>n;:hMAH]TioUYc^REGY1XDJ4V6
\FWOheO1CaRBJYT49UlKZ`LWfL2I`DFn[L8N:dAG3^RA=@m9LUi7b_?X]V@d81p\
A<N<<6M1oXOg^D2eeU>A2?RW^2W=^di;f^Z=DXI_LZ4f_AbZ1YmhMhk=AMbPZ:o:
R[W1:>NdCX8NO35g_m90ineE^C`_NDMPWPiWSKiJAjDA3YPXc86m5SbEjioUeO_\
RnO?RlTaJ3lTIq>m0ddbATDAPOnBo8k60?GIagaQ=dZT>?c0goKLOPFMcifVK:8f
`?AOl7;Kng2fS@3?mkofV<[\c\fGI8g6QANUA;?Q=d7LMEWbdJf>WZW[R<l\^g`X
RD42Od[Be2FPeE>?RJ\Y`LA@YN5aqe0[HCTm`_IBCgm:O83FPXH\LK_NXDlEBb[E
1K\6>=ULRKSCFCWk9?l:;?hjIHkaMi2?>Oi=:<`B;>o=\jhcgfQ2GU_nUBjD799;
`RR1Db1ADK3^Kf[B^DZJ<07B`ZT;Ve28HFASJ?5:\Ibp[hO0mgk4P35mQ3EDmg[k
k1h4G^==c\4Z<JG3>V\=_a8B;5><W9FkYi[4@cGVE]e6YVk?h;7<CMN>V0ckFXK4
dKD6J^=Y956R7Pk1]JSfmTTSX^YSXX3V1MVh8YBVJ834[V]XT326]5WjElpK<B7M
YLNHN`ZA0cEDo46Z6LP2?fk24_]Ij42M8TnPd:n2lT76^c<BEMB5S_<MW0WC3=o3
ckQadK5jNjVK?I9Gd2aY3KBQ2q^=h^^X9662Fk9HaBETnj?mTZR@@J4<:HgPFa^@
4qh;33JjG83:8H_@n`JF99MYYOEa\OJA_X]g2HRZa4T4O`Cm_Q@Bo^>i;H7L?61K
HlFEbR51L?9JiXh8N^PLZ3HZ?BPa\AmEa7SFO]n9bAl`OS[Z3_PI<5\cl^LHKh]N
7@hEiRkNRZX]PV[>phY@cN8GoEXI_0?9F_1TUGSDTlS]k]i9LLjR3Ye=GlUd=^6k
JWni3Co7faN1LmoXb?I9NJC:nmSkY;RPR?a91H^ABQSnn2G3;44;gQ]<B89C5JlL
@?kI<3DAKRH0XobSBhU59WLM:6fSOoiqW@Q;=TDN<5\ZlFDi2P8efgYN=`O:kfkV
CB8O\odjhoZ41VFk]]i6D^ki3OZkOl@4NL^[23o4gC3m1ZbhZ^M\e>D55`Gh9lBb
`>kVEd8dGW[DEcT8<h>VOn1>8;T0LSOHWlZ9[4gSmQ]496pS2i_QX2OB;6P@2PKG
WO`Q^h8_??T?Q`kcPI6:n^fGBpnf8;VY;ZB]F3gg?14FnY9LdHmkaN[g0>[S`L1H
]?Ndm2`L@c5bYOg<?lO_;;gDFIf]V1`39J5\aJmnk@HFkdG^X5Kk<OQ?65M^O\6^
ac@Ig6Jk;Nl5aMComi5fCFL9H3n]k9OPhJOL>YKapPmO^E4HSUZ9h6a`bZ7N7I;W
fgJKZD^?6SIBPLQ:Y7EGhV3`f5AX2OL=1gFnJinB41o0g^dZ=\;FPnc?GB7CXM\i
ZhJS84>EEXH^hMhKLQOGE]b?h2OZ@HeMLJ0<jZdfMPoNA_910K:8=VJqT`C8aeEm
f=H0GKFUHdjilUkSde9J<JFaMD@@5AeHJ3AfP4ekB2e=G[BT2PlGIh9HZki=N8]N
;CZnli4PcYcMbMBD:e^9]1Go2_DdaX4HbDGT2WRijB9_@A90l^88FKQ1T4@RM`2Z
hFd7[hqMCG^keTAkg1Ec@d8fdc2<An5kF>ma;EA^9@GmWM2:NWc\^k:5O9fTemI3
cHiMnl8A]oj8b^k??]Y:W>L_W1jd4<jLFUTKQ2Vo6:<iB;mH1_5:T:h<cVE5l9>j
9^o84cFMHFoaQJTa:;[g>q1<SHBdP\GmG@Sc1g@15bWOG\?0]LKBAjfoMU[Rf6hT
Tl`loL>a<7Ni`AcUC\N9BYcX7anWHnJR:Fc`LGYdVKoNe4f0@LH\RUn6;;3_ieCD
\dRkH57I=ekScf:TmnnPe`1XnH3:CoE41ePmqYMbT?3knDn9hn:3W\OhDh[k=^F:
gM\@ATAWed]W<NTFIi5iU5Vd4aC1JYL3dHH@NZGIY:[C=gB^5mTnOEHV_^1`CIjO
]EQpMeNld^pieY59KY$
`endprotected
endmodule
`endcelldefine



// END_OF_CELL

///////////////////////////////////////////////
// Cell Name : dffrsb_udp
// Cell Type : Primitive
// Revised on: 11/02 2001
// Version   : 1.5
///////////////////////////////////////////////

primitive   dffrsb_udp(q, d, ck, rb, sb, flag);
   output q;
   input d, ck, rb, sb, flag;
   reg q;


`protected
hLV\1SQV5DT^<LNYL^OdYRegqa2A3mSHFL7]4c<CI2AW\ThKhEYeNj@=HL[hFZ6P
q@a4LgF]mbM40[0QYSVaZQO:8KKn8knK7JQ8M>k]<C9\ghibS>m5^\LBXpW93En4
p67dAoBlq81O_Hg4><Y4?f^\E_DW;b?=4Uf1GlB9NGQqAYTgnh;gZQOIQ9PAgERe
\D7M^[c^NFV:Ddp9[QTJ1iX>eO^4<G?ER2n?Pe_iX\>?Tl^MKQ^OD`ocgIUFKk63
e[mnO=KqCfOdBK2PMUlWa^LIHg7?j1d^o14jhTp`1Y_E^]EdgD9ICT\ngZT6W>V[
PIW\Jp@1ZYCdG?F>[6K5f>Fd9PUVoVLVC3`^q]bVHUFNm::W=71B0I>=7d:hO:DU
l6JqN[37[IeJnZ2o>:UHM1P3<4_LdS=\57q2O3o4hk8<bKdZfM@9N:`V0Tb?B1FI
5qJ\HJi[MdA\YK31OALAkZBY<74CUeBRQL59q]Na^SlKTF?OGYZfVY`O?=X3?<Ae
Z<Phc^1qj?`;hfF=?:NT[=D6l1N2C7^l=D5A46:fA_MH;a3H=QNl<>`?6]^]H]Oa
<jn27IpQELin8kRI=Lo9An\@A9Ue=h`HKG;8^qXjYE0?i7ZX3=>diOnd:ASW?dKV
]k[Eq62?g4FEfW;1m6LG1acJ;QKVPUH840Xp3?CO]O497Vdm9RO39k67K2^0YV7O
GBpAHFfo3;OT;EbCnaijWSKK?eL_Ya3AAqnZo547LM9?j26E:PLdE<5i=gQD5qj1
d=co1`Dn33Ph5@Iak7b4TYJ:311Mq8:10b^?_Y?c31kfTZ;D?AdUZ?Vo;H6n:J2q
neY1F7ZE;;QM\D@EeZ61NdbHoTokT[nXeGpeUQ85@7@oa5nK?YLB6?PEb=h>kW>C
X1^:?p924T9>2JUbfJRR]^;a0D<LF<<`_eTDD=`H;_Zfm91S_Dq4bXOQYU>I8J?:
YN0igLG33d1e4Y62E[HAOpZ5aFFfC7>46iH\1gWmne7mfm[UD[5Dpld;cL4Lk<\:
H3E=j>[giZj>=g9Sc6lqmc:Qcnk5QOUk;;UF1`B3Nd`bE9369PpPHoSN]0ZVfFoN
Ho:nH>lMc@fHX=opGi\Rb]XB;FfQLUgK254J=mO:OAXThJpGO>OWSl?kjf5`\J0g
hWJ6J[WYfcYfLNEZ8pJPbn_UpDG;bP<h<8E<Rj]127;FOFU`6^9K_\_Cnn<pGUH?
>AKUd3KccjH42cQnC=F=Y[1h<nk\SnpGhOlV`gMJ@6hd[Ng8[9;A^Sg@3Z>9iqDB
n5NJ3HA37W=0@]6WE4Racn47L_LSQM9KqL9lCFRkaQk^mmCc7B5]6dB`n0=PVN0b
_HNR:_PbV_EpGcfDL`9aiBZ\AXcgdFY5A`0Y1UognDZn86pWRJ[mYO;H8STPgc<L
1F1_6_<fGMJ:aPMaaq2D9n:YSm=4[SOP><0G<o3n9RBdDdV>Kd7cp^;lXliJWa<f
ZfFLAnb^ZR51Rnna5eWqh_5@XbT$
`endprotected
endprimitive
///////////////////////////////////////////////
// Cell Name : dffsb_pri
// Cell Type : Primitive
// Revised on: Fri May 6 17:03:26 1998
///////////////////////////////////////////////
module dffsb_pri (out,d,sb,clk);
 output out;
 input d,clk,sb;

`protected
S`aGLSQd5DT^<mYh0j`?[AeJTd^1hVje3Fn]SPq4XK8Z]YRFTKV=ngcgNkCQ9RH>
H\cKJ?I9:Q?M5H;6Y@eplf14XHVm5U<WTDl>ACmSInAPY7p]L4D7?pBahe;iSKZR
h6Vc>B?hd0K;K202WDLmqE4P:I;PZL1OV=ge5bi:gH_1YbMEKJ:J84@hE1GeCY?L
gH0A5q\Wcck[G7m\71_36RVG1e5eeamVmkjBgB:eN<WdSPp\eM_B9T32B=]PVc=@
mn<9NK7oeMI:f<PU=\jU6]JF19Hp_0XYPcPnkWN2X\H\:D:;KM@K8X0gIJTJl`qE
MVgj7jB;9]9f@75jgmckfP\;n?oLm\38=kY7FOkDOR0q394Z:[16mf`ggO[U\[7j
1ScUMB`\;5<7kKZIn9hidW7D0Jq<PdjeRVRTWS__<4BCUFNn<E=Q;nIh>^8fH6k:
14?$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : dlhrb_udp
// Cell Type : Primitive
// Version   : 1.1
// Date      : 10/02 2001
// Reason    :
//      1.1  : Initial.
///////////////////////////////////////////////

primitive   dlhrb_udp (q, d, ck, rb, flag);

   output q;
   reg q;
   input d, ck, rb, flag;

`protected
BO66NSQV5DT^<JHhBNlTD\1IR`;b2Z8CAfIT5KfBX1B]>YV;Qk6p3J3mCi`^dP0_
ZL6JFJJkPSiA3UCW=WOCiI:6q1m35AK<j5=<?M=:5[@c4C`ECpEgBfkRqf38jA`V
qND8jXVU@>7FI<\_J0:YCE:AMDnjA7;Tp>I3OG2jF`DIRdFfmnH;`5jkAIaGqeUN
YUkHOWNJ_BA3=>=on1?oWKR\WhN4qNDXUj=k9:Eg8?3T4djkEb]OYDo@=:e;pmf>
];fAKSUHZ29R^ZQ0[YG?Z6JGM7`AqeNoB`mhdn26aHY0YW:SkFPh0CaW525Jqo<0
NJGCU\9Db:eBWVjTeo=6glDKjo?^pBB;2A_T]bXXbdEmedVPLW>^79BG]=HM_JW;
Yhhhj9^Ph2dWLbGOa[D4i4aG[7Iq6lg[B6=^EG66A>T]_9o=;@a2^YkWTIcqNF9?
:BGChXV@?d2631TC9b2`WXZX38DpJYR_5A7JSa=`MM^T@XgE[dAF_3V]eQ;qhZQd
oGD<dfK26HF@XRPi^:SW<3IP1aOd44bZdBBD5eli^bgqRIi;Xlq`C\HSW`AkZPm4
OGUlAjJP`>1\]m5C<gqRA;85]kT8o<9ed7:YZTYlLA;0e6<G_WqnCC`E_]P@S4LR
_MK5fj]=;2N0>7pSh8Y]h_F7U5]SclY1[Z>h;]ne<MWhaCqSH14S>jS7a6kWEPXa
SmIFZ^[\In3[g9p@V6O;6:eIecYP8N7IGJHb0j:Bj8=jY]qf18089A4oabbAKfmE
XSY?okcTX7Sf`7q21lFd:ddmk2D;i01>Sj]8i]mWBGqe?R9c5=j1EJW[>=G`Dqg;
GXA:@c0hI`o`<:JbBkjP[^oiXqOV2BOIXD?F69QGfkI\V3Rn@J_[dqPRcK28H=je
a^:oFi;IXLX5KD?M6][hbq\]@h\Z3k]_cG^mU:8@@LBoKlDKP:9h@qP@bZXVJlHJ
a1Ojh7o>5BTY3?b0NpESc]1fj$
`endprotected
endprimitive

///////////////////////////////////////////////
// Cell Name : dlhrsb_udp
// Cell Type : Primitive
// Version   : 1.1
// Date      : 10/02 2001
// Reason    :
//      1.1  : Initial.
///////////////////////////////////////////////

primitive dlhrsb_udp (q, d, ck, rb, sb, flag);
   output q;
   reg q;
   input d, ck, rb, sb, flag;

`protected
;ST[^SQH5DT^<K6iU@bb]1[_G[93a:EQ]V>3SY^PAl0h;bcf_1l9MhniRbMB7BQD
qiHM4nK>0glDmK0f?\b@K4@H<ZVXKjAIeOGe?nYAdKXci5Q@V7Gan[6WF3MQdccH
b9?pO0B3h47XQX0492SGjQX7YGpHO]UFbqOF6AhF<qgg@5TA`[JmN\Y]f@R2HC>O
gK<GmJNK^5c4qfZZRV;309;VNmNO>gZhZ];`VgKAGKeFa[>WC\SVQ97pFm1YIGL@
98M9Sm_aC1^]`P2TUgT<U1qe:CnNLZDGc;ME1>693oC_Fc=JECTXoh`hTqYnRhLk
o\EHTNWIc7hHfa6gC5f032L5l^Tep1C4PMdIEgGP7O\2MZLGhdb[6G21=onC42Bp
M70:W1OOZR[WfOAWTKETAU282o5ANRbASHl9Tj>l@=Xb0G]7q]IXMfo]8a4:2<n;
Q@ISH]JM:[oQQ1185[5pN]KhBF3n6H:g7DIMgB<NHFU`WYo?AHhgdVqNOkNmMJ41
iBGo@l_iS\[o<IBi\687f2Oboq=PPQPoSbD4[iX>S]ahBn04;`Cb;:OjFiS<qo[O
c8NXK\@oGk<M>BQVeO^P4cK8`\gSRgPnj7RPli8jgbh4OV21AoLb=O>Z^5<JK4mB
qm@h0\NZ80`R9M\d2KU:2Hl[O[Zm:H=l2GnqiE@N`TqFBi=oSC06a[K6M\ThkA@I
imgTX]G?aS30XqZ?jZClo3\H[3>71=5Y4Ug5eSS^i32nb^1Yqg]6@2nW]DaTTTB:
I^_MBFT`_1C`O^]a__6qO:mnM`kS95^Vd[3nLRQm73fHZk`2n3aZQMqYA`o[`Mja
JSmnKJ@n3;=LWo6og7iokpn?FEkeh\VH7lTTT^9S`Vo0gQlIk:GPq<niH25XR>91
3k_^onCHOlHeJgX[?:Q<^OCp[BQVBS9FI:hUZ[SZZB`]RZGl990VL5]7P_Yb4^1C
LMbIjTQRjL<Y\RJTDoWn9ApXT;35M6fggn64JiIX2X6Lf_@8C\eT[QR1^pVE<;HF
dU[960CmUcaYA@eYLTA0]^]NV6Z?p\6gh7Plc?^D2ML7^9OVhM6o^aHY30GAkm=q
6HS^kE@;[jjaK7mSo3PDbMJj>^\5e41^KBqmohDho8EQ]NNRYWl70DMEWDZ7Gl<`
YpgK^H6AUg;6MiX6H6m4IWUmj;^3gK1npAX>MHhE2ZCNO0o1n;^JCmRHQEFEWU1M
l7>qOR0hPWQ2?TZGZ>0NPaMfCl83p>G[[H]mNE4`_\Z7WbA8?1L9Z\KdjdDqO>1c
[bgG1^VjG[1=6n5I@WJS=]2Pj0:i7kpHEo^NBJWF]SP6W`GZ5[C4_g38VinOOa_>
mqCoED4jdk\=`@[>5TV00eUKTV:bD4EEHIa`pB\_Hj96hDd>TLTTHcdT>Y?TZOdM
Am>J_YcpjoIT<@Od2TQn1\djN48]BV^?BEGBUGoBiiphHTcYHS2E[R4f[g^3TkT^
L]3Ce0`2_qaRjC9o9;eiE]:YcTW7LJ[2=i<bT\6Sp33liQ`2R\f0h2O1=QJWU3PM
:KJ5hlc1@jLmFTg?k=E\:Y<HgPO1\NO6c4X:q\ZRPJ:LHRTTanZ<lR8oJIV=X_`I
N@Y_jbap6h;3gikCUfKlBaaKGI^CGoM3b24kOWpGll2UnK9X9X7;EFL:Ng6=I:K7
7fJ1<fNe^q2>[Hi>RIXK1KTFHP7<SQ]O575Y6kiN@44DpgPLQD8p8@6\Hk4DNGl`
VPm64B=F7QCX_k:GTcp3fELh`<$
`endprotected
endprimitive
///////////////////////////////////////////////
// Cell Name : dlhsb_udp
// Cell Type : Primitive
// Version   : 1.1
// Date      : 10/02 2001
// Reason    :
//      1.1  : Initial.
///////////////////////////////////////////////

primitive   dlhsb_udp (q, d, ck, sb, flag);

   output q;
   reg q;
   input d, ck, sb, flag;
`protected
eI5YkSQH5DT^<:g:1TQi]5=5@^WcAbSUd1hT[PAaoR18oj4_5K@Ncm8daQa^gDY;
n0NDleFZB;\kHDWpahlUF[D\H7P[h[0[MjoHc2plm5nXmm7j@gNeeJJ3?AVNi=;T
HXedgDl3?QBXZcIJ37=XIjoXdQQnoJp5RJanDqRkSJ3FDq:OZ3R8PXlcAG1`JaS;
0:KRcc[`0K8g1qGH@b]ioVC<8lQ>Elh<A0Q=4;WMhpV[dCOol5\HWc^oA5G=Q?hO
[TZHeYB;UpO<5S_oTlR8_k8BIV;f@:6V2RYPS2_k3qa[;k\MV85fX^4n`q?3Z^iN
3lB]Xh^2Q:B:I615cG_9flhbLpIT2E>e>KGTZ2^if51mCkR5G3ankK=:Cpd_B9Hh
Bnm3j3>aDZO=ZQZbfGDaLK?]GqB^nJhUXI[87VTSO3ZSITkmaA9:N1E0UpTFW1N3
A:hn];bfKQ;ga>NM93QV?Q`dkqbW@K<\>C48=0C5H_[P^k<Fj]Y1J1Q8bq`oDI0G
aU;j`Ec:LVWTGSLgG4NEV\felpK;9_0Qn\C4X<d3=Z^m=kFAUJTf9NKOXq@ZkkPI
0nUL[anngEDWo]7;o7Jj<h23PVQQ7eNKPYR]GL67SKql:Ki`BYe3E6K;T<Gl8UPe
Cg=9mCqCGfe>`qf5\N^ZBh1P7hVmoVAmm8DR4bMYIOP8Gqc5d]gbNBJ8`khWOWNm
^VmR23]bkiKU3qbi2DRenFOY8j>i`m52iIh0DH9gTbIj2qh1e>8:Nd6NnBXg2^PM
SgDYA>4g\2d^DqKVE7PZAMTH_JH?T9j7N3ORkkk_Ap=iMM3BoG@XM7A7mADbci[o
\:KAVqlBZ\iLG94O`W5Im0hQUVj0>faEGp[d[Rb:?E_LXJk4mpfmiieGEC@\Gg^[
=k?mi4YRg2XjnQEdhpJ[6cK\S>1G]TP]mGM?9A1]@`8c]AXL[qbVDQ@UlU6>@cMh
JV=_1jNRY8d`_pg7@K_9l$
`endprotected
endprimitive
///////////////////////////////////////////////
// Cell Name : jkffrsb_udp
// Cell Type : Primitive
// Version   : 1.3
// Date      : 11/02 2001
// Reason    :
//      1.3  : modify protection method.
//      1.2  : Deal with unknown ck.
//      1.1  : Initial.
///////////////////////////////////////////////

primitive   jkffrsb_udp (q, j, k, ck, rb, sb, flag);

// JK FLIP FLOP, WITH RB/SB /STANDARD DRIVE
   output q;
   reg q;
   input j,k,ck,rb,sb,flag;


`protected
k[dk[SQV5DT^<\ca]1CQ@UMZ>UlQR@a9qP9S1Y7KHmZRK6M^0IRiH@g96gTnP3\k
Ggfm]0n_;00PjLo]aDHb@R55ob8@7h]iAFB;l6d42pEi^9[Cg=9H@ej91W1WQaNV
F0@al4Y@HN6io9KOeK?Zi2af<qWV?mb?pZ<InciQqa]H=>D2aY]L@:i@]mE?8]NO
[Yg0GMgWfq@W7fSlpjn:KN^qimjMN@7SX]k91QgL>gT]mSUO[F`WGJL]p[cVC7?<
8n3kU]QCaDT[DZ>Q9ZIC>44o0qLA8CcUHLD:RG]jNfmO6?JFh1M4[27GLCqGR`FB
JdOEJDbefkKgL6CEO@H=Dg4OYm1oN]GWUQDZRI5IMFd3IpAZKhl6`9cF0JOmllK0
UO4cRS5ahkoH\UpMSe5DdH\hSA=]hij6ecjKZ@ZUB6e=Qb>pF4B66dL6l<HNn2jB
>X4DRQAh8L;0i70FpXO>b==h^KNaNbded4K8PJ8N?P0WGCXokpjeLA_7CMO60cg>
`b7iJX2j`3TLj1IDH;qDGQfgfON6lI^TZ8<2cAjDk]DHlX8^gf4p:5Yf9h5]cRW<
ZU`?5U3MAJ;IbalJdV`[qb8ha1:AF\HfWdOQ2X_\7_BO[c;MMKRkYOhqa3W=;NCj
PjFKK>X<?_meLfSL2cZoeaFAqQ0JFVKpKl2]_KqB7>PA:8V5c6SI]<\nbV=l_\QM
AAp18L261qn76iXgQ;Fdkgd3?d3\i6PRd9=VmIGJV201b[pD51BHYba0>dePFd;l
?S\MPaIYP_BK8BO7>W@ql\ei?^C@;=i<03PW_>[Yg?Mogg>7FWk3V75`p]S^K61V
L=O1J4Zea?NT29Jbd9[UXE:ocDL^Nq6X6O[Jln@0XgXgXel>:[9>Oj[bFR70=4DG
Q_:fn^oMHTTGdf_m@Rm<pR]2_J^7]7FO;1UbNdm0bVK;@@2J<F=8h<AfIqjlD2N:
NTNZVFD\bNk:B^[g33;6\IPG^OO1fHp4^Ji^l7ijchAPbnj\?dg5<BGGdh^gXZKq
J5nR3KNL]LjeT<OEm<8Z8@Q4`emDo0Kjp\9XhcanXKkNW37jP<:AU]5ooLDD7]<Z
CCH;0YkBk:e2MO7UY3K;WWGFAD3\f<lQHT7:mqNbV8_lq^nZd[I8n5jg\?6hIH2E
@2Y=b[I51@G7fp=o_m7[VL9STO:WZ6YPjQ1f>bLW>0J13kqPeEkE6J0HQ:60?WJE
HGmSS`F]id7edPepJ^mZ@AIjK8bYLJq8157j9c`e`ao6V6;kPP45P7;n3SKahT1p
X6fJ`Ip5L9Fe`?GKS>eO7a=[W]O0[Se3<ZCU4hNqSOn9;I>dUA5CK<B;i]P[g<nM
KDgU@`iOq0TGPfZk\_\<3mi=hCWU=1KE?eghlDWA<EI@kpcinEFlq?SJlQQkH4[:
eU`FJHRdh8Pb=BGgjHnJ0;N5ZpnANTV^Ud6XT9\o\NSSMJeP6j^9[6na2Wk3?np6
LeH8U?HNfheFU[N9eM7W`DIdN2EdomfS>gJqMDJZZeiHa<gQAEOlDM>9lQDPh?k=
pP2=fn@@AF1?\`5N:X5PW_]G4@jXXUd5`\JE`qlQF9SIgm@jhVeK]jFUZZc=^;L;
U=D<N[4LC@pUjCU=1\2o]GK2jL97aCYYa1Q?_n[giA:YkUHpOWB9W]CjD8>g<fMZ
NM<5m9Ek58M?8o`hp3C[BaBl$
`endprotected
endprimitive
///////////////////////////////////////////////
// Cell Name : mux2_udp
// Cell Type : Primitive
// Revised on: Wed Feb 26 17:03:31 1992
///////////////////////////////////////////////
primitive   mux2_udp (q, a, b, sl);
   output q;
   input a, b, sl;
   // FUNCTION : TWO TO ONE MULTIPLEXER
`protected
I2NTCSQH5DT^<7Xbf[Ek52af83g?FTm1GNcDEC\^TSDTlIpR3OncAU7OVUd[U<Ea
<YOc1cHF<?6I9HCUdUKGeoXc>`mP_Wc6Wq80I4\=99eGFU<fgW2PmKi8PGIHBQCA
=hoLkO`G8eT_]95S0`34PVW]j:K>NB@mpDP_X8Lqdi<0<g:p7h6M``q0Ol]\dH[k
[n?P\:lZD]CqADS953U;ZfYV`Z2aQfZVp1R0jX3WOak0`I67K`FbXp\d3?<Ck[LG
P_CHj@UKU3qQFD@5R8@U8@5OXGN1_e[p7SJXP:9=<gInca2f2R8kiMlO]kW;F8Bk
b_B93;VqoY^;2?o2O??Vo_OWYb`Kqb\>D^@E$
`endprotected
endprimitive


///////////////////////////////////////////////
// Cell Name : mux3_udp
// Cell Type : Primitive
// Revised on: Wed Feb 26 17:03:31 1992
///////////////////////////////////////////////
primitive   mux3_udp (Y, D0, D1, D2, S0, S1);
   input D0, D1, D2, S0, S1;
   output Y;
   // FUNCTION : THREE TO ONE MULTIPLEXER WITH 2 SELECT CONTROLS
`protected
X<RbHSQH5DT^<Pa1mX`lhLMeU9IiH;13;ebdNIoX4g^Fd]=9\of=CZJ9fomp7gX_
jNZWmE`Om5dEJh<eqRH0@:2dJ:D<PGAh6O\CSqHV_OkRqihSEE:2p`TmbAPqhYX?
NoXe?n?JH^bdflMV?\g=C>q9E58S3d]fnIPj7[CJ:V5k2dOVHp0QA`M\55]:C8hn
k@moKbTI3Eg?qb=TmR6_QWhS?Y`P49__e\=BnL4jOVi`15l6@Cg?enf@CV=5mXmp
===2k2@4dV9>Z8H\eA3:jd@M_4p;B83>L2m:6VmmV=BgfENoOF<OmqE5[hWlHESD
WBY1]@=Yk<U]cn6`p?\PEG_X`I\Wk@GX>``I>?DcX>6p:2WC=N[PmPX=M;_mUGl5
=o_[CkpNV8gRf8Rej693e]EUWG727T=TTq4XkJefX4U\]WQID`@ZBWOQI_H=HED6
=mEXBZ=nTU>]NHLA]aZMWJ`l<80aq87D<loR_iA:U^2FMK3HX<BB:ZapdHTDe<6j
KTWZ6D^1<D9bJ;`Md>qJFaKMeblEGc8<lJ8UEf[>YEIZaq@\R6;egC_3\NhgGXjH
6j6[^X4Gp]CK?Rh`@>emQB=5BHafV=O<Wl1qmXC1?iJ$
`endprotected
endprimitive


///////////////////////////////////////////////
// Cell Name : mux4_udp
// Cell Type : Primitive
// Revised on: Wed Feb 26 17:03:35 1992
///////////////////////////////////////////////
primitive   mux4_udp (y, d0, d1, d2, d3, s0, s1);
   input d0, d1, d2, d3, s0, s1;
   output y;
   // FUNCTION : FOUR TO ONE MULTIPLEXER WITH 2 SELECT CONTROLS
`protected
:>9@oSQV5DT^<Q^K559UnJ[RLD@TlHV46=BcdBS\KRhZDCYHZnl^:OD<ni9A[?fL
`JhaJe;fogqI]n@W\m5GM6Mh8eG8o<7R8VlJl\k:QV7lJ7<mdNGIDdRaI@jWXBDZ
j?:qDMOM;ZG3<_]1MNE=_lFmDFoBK7q=J7=:?qSRjP^m:pUgCHI?qQOkIJ[:OUDF
Q6RKHJP`_QmKHhOg<pgl?30o78eAIY_W]_CiQh>a5SXB]aqE_T_Ojn?j@KKnGNXJ
]l8:dc3;ckSqnE2VbRl@ZF;10HHi3mKA?4@WFYa]]I2N\b0;I?X<pm]hD868?UDm
<Y2<mTi4b1cmHg`eWqAEed6<=3U4012b\hQXS`j5cGmaamqMRSS3jf[VM8LO6NF3
I31X_^>RQPcpe5MHWPRih88R;]f7RYWlM0^@EQU3pbR]@L[O7V`Qemn_38l?kGfC
jF;i[pB6ZB]@=MRZCT;EmkQaA][oOQ[VFd:P@WqjRNn8LXj5@d\L^mM[3nPOWFA1
N\UpW`kBFcCehk_TAbkXJ<S\kTjF:\9kq9?<gI@3jZ<DiK35`K<oLE_m4mk>Dq^C
Z_013TZnVkoCS38Q6k6d[XK1;]q]\]<eSImC5?l<\mK_UKKl;B5o4fHp6\O]iBef
n<??kI\bG9C\L3MUJK0>qWCJmB32<\[DTJ=]YWP01L?dINnmVpm@mIjWH<_dOI^Z
E6g45:[bMTL_UnqfAe^ZVD:D6h>Di\SeXK1GRQEY7V\OE[V<dU^oXeM]\3GQ[cR:
DM3^U7dP<0]46pJN80@ZD_W=gGO3ElV`6<A]m2gMhSpJoEi<QMKCDa1i4@@K15We
1`:36cZp:A^cZJi$
`endprotected
endprimitive


///////////////////////////////////////////////
// Cell Name : pulldown_IO
// Cell Type : Primitive
// Version   : 1.3
// Revised on: 8/20 '02
///////////////////////////////////////////////
module  pulldown_IO (io, i, e);

  input i, e;
  inout io;

`protected
=B<j2SQ:5DT^<3jH2a3gglT:69<qKZU8X5QP^k;?T9<AA>Q1Yc^MXiPXqJnUbi07
Y?C?:CR\bD7M>IIbo:=<>Fi\\qd<<ZmJqVJW=][`agUh3K7:[7FgXNkDUj``qA<W
=`@9:YoRNj=qEGGjjio?e9cIW0_6qH9K8R\PakfC_hcX4Qi_BdAI9VhVqd[\TYDe
q<F1JL=GlQfB>[40Qegi4`hK^pLQ7kAfYkgMReG]_L0oJqb^\gUhhE3DN[E@K3DR
3o[g_pY5kjCcD>pjjh5e7FFRL2BnP5W5NL3H`ollo22>4pPl=:CDiaq[b8>S50U@
a<Q3LiqF36:b2MM\]iOCNm0ciF@132Fq<ElW6FogW[STRMTT8TU?S^LZ6=mK^FaN
L9qcNa3H9ja1aYkOjkTc``el9pA^IF[TV\<OWgih5b5gQpm?D;h5TB_8jBZBB3_]
2PP:qO1VSPF_inW^N_6=]>eKQ?jJ3jfZA`K^pBUOiEYn8>J;eYZii\\VG5fkmT4F
84jNhcbOCCFddpc<^Tai?>_b;3m;6DN\LioHPL`h<P_2Y\q>fR=kEF[Scdj@N[W3
T>Q3b?Bog6WWRXi_1F4BVBaPHEOX4pWnaliX@`P;Oj?A90:9LmYaHB]HVR27b>dG
OIebRWKZ^9AThqJ_AZPUA5Z9n:Vbh7hmpb1mh:n\C5_?7OIoIi8[846LbkQe_l7W
CJ^fGMb1p\H7]57<<j5iiEeB=WTYnp[N?<iP5q9817f\ffBh0N4mamIQ??aC3>lk
<D`GacpFIh:\h>pDZ`ma]cWb;Xg`In6Rh76E@pRP]hX^=q`j\R\ZEaC_Mc3<>mA2
?=hOGp]_EnRk>aRf6YS[l1\\06WMlG<X2XXU5_YT3qc]nVFeRp_3B<jS>>9TiL;M
?T5Y<RjNjmd__epQN<KHTm^g6m@hkXOH\5MaB1_e:Il5Je\2V7]54@LnY_>C3mqR
`WdilXimNXd2oNd_4KBmDWTY];q19>Mmm5p:<EM]Zgp]R`NSEJ1JCB47EdF]LeVg
Hc]XQopPM2V;2lq^I7ieH\p90;KTYgq5CUBjbR_2=d_Umb:nheH6ejHVM2?RY;GV
N>p<GgfZl:g\XPl96]_pL\`cD`IqALH8MoMkb[ND;K=G`R8IKjaU=I3dNTSq1Si^
b9@pD95d^eVjFn2C]lHoWHWD9Fn6oQp2\`3NiTq\D8m?fW_o5d\2jjDIKIg3cqc5
I`SMjX4<Jbeb:1[bagZEmHCC2pnIaUlOPHI<9i]`WH]J^aoEV39dPeP4pE39>dga
p^?VT=7^6OjAZSmA9C=X:2@imDNeEqJc@\Qd>p6XH?bD9ZE][nkkXS@l9lQPqoTg
W\Q^nNWAinW=BfHF@QJi_fJdXK9SKZe;]EipSDe]>TCFSaM7G4KefR[TBO0ZJ9Pp
gCb1J_oqK:dTVVeIOa4eXB<W4=U]TcI]di=2pTfG@5I_q2OlF@^<3KP\=9Ga224O
?Dhpn3QXaPE@?9[OWhlJ5cDNMlTG^=Qpe04^ZZ8WBSn<5CVLA2NkC_[9D2YdY\f6
aRffj1`g[QZ=3F9NoXTA?N;_2YpZ2B48o1c80NDj<6ciZH@Z^]B2ajpmfE>fL1p<
5_kma1po6PPKK7GYaEG`Z;hC6VKVMdM5jB^o]La0k4ea4qjCUcC[LpZg7Pe`W<4[
T@9=1>=Da^TWTfpGM7G9bAg[JilM;Wc=LO9qf;=]8\S=TaG:ZE[qelL3?jPNdG85
WNOmieK]6:AIKi:\Pa>YEL[q1Kl3eK`qe=>D@62$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_down_IO
// Cell Type : Primitive
// Version   : 1.4
// Revised on: 3/19 '03
///////////////////////////////////////////////
module  pullup2_down_IO (io, i, e, pu1, pu2, pd);

   input i, e, pu1, pu2, pd;
   inout io;
   wire io1_tmp;
   
`protected
k>5dhSQ:5DT^<H7DNe7hWceB[^bP;c@nmOHnf^0epLUXGfAV2KUKUQAY1@;`>b8G
;\W?cM6_b]gm]EW[5iUY]B^;N3]ikq8SoARO32WL@IDNL3b50^W[dRi3[LSMoegO
q?Ci::?pB^WQMfI[UnW>neMZL>i]GoL_C>lpe]fi?UiqFEjZ3DOfFR7PQWVF>4<F
WP<p:Ff6h93XoAIQ>WY9aZTmBcCpBCSZbg?qHnlQd>HUVR1eg<U2@?K[P?0RELM^
h5L4phc0WJ<]iJnWn;\;2eZ2=BR55bV=EoQg\g5;99HQNq\aTP7X]q>:JQX;JJM]
?9=;TplQ9k;hk84ejGjg<Np_o]ST\`SD3[H373:S@DU@`lq>>d?EQ9^AX2L\KSH2
R>Y:Sf@lC6EYE5F2EVnFTOXAY4IPDCoc8gLGOf^pGEVngLV1iaY>lDGom5N3J_Z9
bgL_YdRA4Kd^YGR]F<gQLn=aYW9kHQqCJE<0jT^<El8SJJe?@T0To3<2mQfbkB4K
;Bp]hC[Sf\\nQM[fLmh^YIGb@W<@<5Q?Agp4VShXD?V`d3_6De6><J<mN4_QKJ4Z
b=TB=3fdOmi?d49Y5X1oKHL\<R;5cqE]OW@7Q\eMJAgoc4X>k=l1q?b;R3COjEkK
VWKdk77gq3DK;YMm8D`TWXfehi>@WaQ5`ZjJ=YbqOiLLDKO3cmUJQ1d1AQ7@cJVI
NJ>Il;R4ljAVp`1Z?>N0d0Io94AQ?U:QFMFijlRN;KIWGEU<Zpk]@[MB62;al^h[
ST74Khmb_VTiX[acN\;Mp=lB@`g3URO_N;4Q@9k0TjejS4LjG5BJq_=H;U@CQcOR
VgD7fB2D^WBY\P:fCE1:LM16Y3jG2p`=I@4E=0QRZ=kIhBU^9?aVBIS0l:LY>dXh
>JHSUePJ[M2Ok6O>aS?Xq5>ViUP@F>T2@ibkE0UHFPhkYm8a]]B_?p=JFgdOHoC8
ciNVCKI5Pb^<dXD2cV_@8El:H^Pd?XK8c[_\3pGA?>l@T;SXb6kT6Y5U8^gk`l_Y
YY918A3a0`NWMCjM9>kB6]T@e?bX4qQc@3nVKObbDfC=@PZ3hm0SORQ9fR:l4:\@
hk_0@IW=3`od7GeAVSX[qe8lP?^e:V_hiQkP7`_]O2_2k3F3`VceZn1`abfDhR=`
]GSCq81<T1XLGa`4f`8DR8L[h=8LG=Po<1:Nn5nGK`1anib[L>V3Kqmh40;PTk8V
8jGKn;gnqJQ90AmplRC14b3LdS?JnmLZh\^02fN:Q8oD3HoRRXdU:o6Q;EBa0_qB
:XdhP@GgY2XMhBAoI:Pj;YD6;JR4>5K[7iYg^n3Ic93\?CqI=^gcB<FT;gcVB74=
nJ^7K3eHO^<]?6Pn9K[MbIT@G\;\2W\MM<OCKSF<8_l4UaP51cYI^h>@ORJ9j4pA
kZ?7Aa1XhQI?\IB=dIQZmPkU;KKihI^;AfVT:gF]9Y^2O;epkZ[dbbpRTOX4a6N=
SG4mm6^]mY5c7<nGjabX@O50^DFRIN5@\H]:>XEUL7VhbR`3R<>16@jSVpJ741PR
F8O^R3DA3TgC63]X?LA]R`H9>e6JPo0T3R8b3lXQ5oa_OXFXo?W]0nge?`qlRC1?
87Mdb3bFPXQZOO7JO6L9FLl^MgeGJ07@fmPQheNMH`QOH_:VQgkmEhpb8NgfGqh>
8AKPnBTIgF0;U3ah`S51S4Ql9Mm0B:On3im6OC_bA7TN\cMa:fl@ZqJhch\4pF=F
US9C[dZbIT:h3klIDF<8o7d4lj5?_:fhKn5EVAQCQ:fHqA5lLY:AqT_bhmYXg\\N
aRVCJJAQ9T4RK54=:aS<pX`QVoAS4IfnHeP6m[XFV=0ILi<M@3:0k\C=ITTN9CY0
V8LO0YKS2[F4FDbK`T8qmhGAA\7k1M^lRDWhXTGcHNW[eGHb]jK>q]b;[n\@pndK
h6hlaJ>]c6^Hjjbe_>:2XonbZEL=<Smq:6gYK97hk1k<K8kLjoNp;;0ck7Eq2G3h
P_^gFl]_:]f5N^[T^dD=\BFoq<ceDAnX<o@R:Mf?@@>_SQBZ3G00q6]L2m@>pZ1c
Cici>Ii:a54I\R\l3k4MBUA1Rf7@WGQ_CLJU`JTKJ5eTl^BJk_\o]Dd?SLj<qBOW
WkDNqhiNKAYcSN24F=9BmG]Sl19T?dm=4b[OpYBTUGAk8eOVXCN8kXb1\jIXOgNV
qlGe_4hMqT8_UI40pnVcXUj]L?aoOoWKKF]`MgL9PBNL;e;5R:7?Mo=Ce0B<1oF:
\KYBF1=p^[jiN^OMBEJmDWW3CE?meai[e0EqZeXV;NfqU:2=26hpKG1J0g1g2K;H
eKg7^0AJq^?`Hn6iq`6VGSFodoPHST?>2X^IpT41[0`Rq@7UBd;1^he]0<oiQO`R
hT>?LcahTqY`NeCK1cXD8V`2_A<\1q0N4Nk1]6mLogO6QoGi0fMW;NP5gpmMZhP:
nq;Bl]Wg;pDcakl@jkaoa<lJ8S8;PX>GJVe8CXbVTpJjFRj3UBAnK6bD4EYCV4@@
h8Z9dqG<;<JS[pQi;1k3bp97_U\nLfKbN0OZD[2<V5Pi?mWFAq[clTZ^hqfi>i3O
=Y7c_@7dKlDCXScaA=ZSH[D?K`i8Z\a6DCL9P3:j^fZbgH]>^Ih]DkFJb31DNJ7<
gpj0[aJE5pLndE7j9p7W`SO\:71WHRnf=WHapR19oR4Z943?DNBkjp6U9hSFjXIn
QmEmZ1;gEpn^OXnICp:\hog49EZOij1;j4CRQkNd3=PZgp_@DhWAMp^Zi]70nCS2
C_jCi7Mf;4];V>>6cCqMZ]nGmfFFWpfTjRN\Pp\ZS;Mh6SSnCH88kQ><;D3Q7P[2
CpH7SUVN;pEd<@C[X^:AL`lYU6mo:\H=::^a4G@hK0qa@5dg><pd[]2Yh6p=[A4`
:?q\n1eKl:\6o<JPa87pHdTAOlJpIi2e916eJSIB]CD1n7<8iYXafR<2iSp]cIGV
S=q:J;GSJGlhD>[KC`d>V:JFa84@NgRa78l4WpiNS]eFF5EdKD]Q4hb58`>Y3d85
c8NmP5@K6:c2YoHKjDE7DFBb6po48M:YVVFLEmckMo<QmqKe;IQo2pBdNO03=GT_
mnOWn6QeBTR3\YkRq17;mn\TjVf^10DT^qf31\lEap1@P6Ol5Q]CdMeG3nk;>^qI
MkYGAd36d=C4?\AZN^a0ZeOU_1paFHgN^3p[oJ?:868G8E?dkg7<ohY[IL6FUgDp
k7AT028p`B<dNDg:9c]Z@lP9dB2ApXd_DYOKjMSP0\MNCZT@BdcCM<BKqeI00MAe
[4@PC9`b;[dnaEh^8;IHVJ5On=ESUc^gKo5?<I<OAb6;Q;Tb\k93J;K2p39K7RE`
qZ;Y<eVFKCV[?SSnFHSM]=SS[hXHepQndbP:jpbB7;MbFl=TQh<nZ[mOaRqRA53k
K0;Y4nSed7^5WUm2<`4VmHqC8_UZl07`Wj0<ebHfDUU]JP_io@pGPJ<RRmfbT<7j
6lYNIU8BG0BD63eH>GHGjGSXg7F<830aRCNpPAThid_poNgQQK8pnO6;JjO]3D:0
T0>I8WVq>e3PLc;p9iEP\h@<J8=iSA:kT_2d_:bV`6pm:0?I>gpSJRK:2MDNlnWN
=5XJILDqW\K4:JceRiOS0S78:lEEZicT;V;ph8HHgOTp6\cdS^]@>9GK8]42<gLD
idFlieekU<R85jU9_6g`QhDQ`il<V]5QKefBhiLd@h2A0=9kWcqckI@hRW11KWET
4oJJJ<0ROBTj7`6pca7HXN;qL9[AJnee0n8FVK2D>2GPpR3bHRh:=^eM:W<]Hh_A
ARbQPc]=pm5`M:emfiSA<01[C5KIQW4L4lEd[@XK?hF@JeHjlOPi2GR??JHQ?NXN
N?_onpQI2n2U9qK0^iJ?BE;1lInL52OOD[kKM?dA=Rp]i[2O`mqHUKlZ]X>\E_jC
0lRc[M2p03CH4iP\CKeO9F[>78H^Xi@BFKGpk3>P3W349hFG2JM=_i^YBYAc<KSq
a1G?_gMq?8gnT@mphCMC3o?k`Mkk6PRJ>@qG<mZEZg2?D6SE[fjUiWmmUmQXcC<_
hC58l0i7S[pUSoif_EN88:`E43ZmAaq7j1P3FGq7[Zi?RqSZZ]G7Z@JVAa8m=6kM
qaR4EWL=p`eJ1fh0cTMpSc^jiZfpCdGWlF6W9lX@LMlF==?4SD<KKMGG=dCSm^j7
Jok:4lZLUGOn2R7^L@po2<fN1kiSjj8N>NbXelQ40X?A=fpVi`2;JYq`W_B7`QpH
i`SFJHpKFY9Ul5p1Vb2B53b^5FafigY6OYI6iQ[7IY562mACZVqRXEeD?g?_16Zf
YIlZdpTB7W3h<;TI4m31HjI2Y@>\fDl4PZH4qmbbWmIi2l;>m4@ZB4HELpL>_^G9
>E@B2L;[P2@H<cpgKP>FmbpD^K;<QPLcNf\OeD1fkP^W4>_qd5kP=i1F3KH^Ho65
<?=qcdQ>dACg_aYHo\9a48]alIFb9n_J?cMTl7DqY>mBANlpn@@89RgQ;[F[bLE5
=^0J]k_LlWei<Kdq>oCeVfN]d61bkf0V9?mAL`]Ip0F>5P]6O^o=[];Yjon=q?m^
3;Y^Y:I1fk8LLhb[m]^]2?;>NHD_HkLBqSkJYQUEHRMc^LY[M@?^0eROJfl=CqP`
14<@bp`5XKKC9$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_IO
// Cell Type : Primitive
// Version   : 1.3
// Revised on: 8/20 '02
///////////////////////////////////////////////
module  pullup_IO (io, i, e);

  input i, e;
  inout io;

`protected
a6S6ISQd5DT^<PP]2REX=<?>VlcJFZ?4HZ8Q4`G7bD0K\K8bo;41G6pB1BoO<\aG
8ah:cOn3O\@TDB4o0I=X[=Z[iEBK9K]XbpE\PP^koR;b3NK7L2oIpA3nUmPq]N8Y
6gg8;;>k=R5fiHQjD1;7ECApJ_GG3YkfFW^_<LqD<I\_2:Cd2Nb2S=K=In2a07N1
`Vp@1YF^9gpdgZ;W;ZEj1Qd`Q27okMURWVHpM2TiO^8Dn3JY@hTlG7QBn3UO=ClK
IJ[HQ?[S]@PJeQFic_S74;h;fK7F`]_qLTdX10?elZ=Z^Qma=XbjH:<qVJTJNom2
p]>R>7k2XgT;gVngSgJl1haHC8T>E??p2h6h?m0FqR]C0U?L_Wh\FJ6RpiI^4B?d
ND?H9olcHD]0hnlYlpS9lI0?[=e_JfC3YaP<d167NHF6d]BKDTI;plBL^gL]Jl[b
U3NZ1DNAYdiBPq^U9YbkiCWB7AS\3a01HA\Cq><lQai]m7SOlhko[[bX0>lpXF:1
Y>6J<8eNg5V`80`jbWkb\@dab7:p7=M?ZP1NRPDjh<J4_Ha:k\]TPOnK47`jM]C9
HWf_p\MkA[IcE[2LDMNF<nEF=d;?b_Cc11a9Ppe2@AhS6^Wl_A3j3VA^Ue<nFMU7
?`IRcLCLJ[1Vdh5OOOR1p7kOmW0lPO5Nb4ZF7O@Hh2M^VKZ5cVSFoQN>obl4:Uf4
e<Yiahk428ep0>l^Mg[[64BBLOBVbX_oc=V[QT\Yl7iabBEobno7=\L@4hLqe6En
UPg[h11`Hb=j3h6;Ki[7[8[=AV^Y]ieKh7EpU`_m:PPgI4hWCgbTlL_XqOl3>Ya4
q>m[=0YGSc>=JlSSj7nCX3CHXkO01O2^fpRAQee>Epm;Y5W[2L5QYRRL@l6\1XaP
q4=\<En[qH``HnQVC><O3N?EM7ciO:J2YJ6l^?VTeDNeqaiEY7U0d9nc7d\B:d=3
MHMqH=64TFEq1mmGdVk8VAX?VXJQoUAbYP;NQ0dGqlSTAe0MQcAeIIC;hWTdhW^[
QJIJqU0X]ZDMe7RV6mMjJ@aAC^UQ<V6@XG4A<YDnNl;TCXWY^c?i6kNgfc8fMefB
qTZ4V@\LpAU1N?C<qm<;4FgPb7DIGn@knD303nB23iWKpMf1f>dFoI3ZI58BB`><
Q8GTWX[5`i4j8UmPBA_TVQ@:pPl1O:j5q3OMZGFlp^bZ0Lbmp[433R5KR>C<=gPf
gqD_@nGm<q828SSiYdS@gG[9An?ZUm\Q@m8oYP9TqhW:[?STpJ1J1\4amEG5?5H9
f5[JXah]6HWqBHllbD9q\GJZ<bFdXjfY;?`]cJ3K1AbPk]i<XQ\]GB;HYE_F6`0C
A1Vdh8jiBknIq?F5BYDTbnJdXBIcldbJX69q`XLgBe><?iIdOL35V0G7:l=FoC0q
e_c6fCbqRAaFTF2M`1Q\3gRoC]cNZ\c2C6bCXVB?VZPCTPSDD6bAWYGBR@R@A_h>
5LET?79LJOl0kabAp=Ln7<WEM3Zn=Fk>kN]nifJ1jiK=CpY1mQ:j7qMBa_=CQ35<
U<MjHPVFPUb6qD>Ch0B;V>lUWnBX>8K8OE8b3g90pbjBmK4dp6N:jN@Z9RVOOJVA
;cZ_Z99jOn?KcpaRcYF`bqkSJK^GO1BIU3Rd1Z3DcJG<q2mTQVb:ld\43S_5D_2i
Z7TS`Jf[G2<[B:;XCEUYJ1PpPV=27UANbIUC]K>0:YWGnKjiRZ`qDV>3ebOeMN3R
X?C4cd8B?cB\^TdpOG`fjK9qd?B5962peE6OBkHp^]4E]bTiFeT1L260n]IoB_LB
pIaGdkNNM2k@GK3iX0NKWpY1`0ZL5<:1775f9_1g:2PjUS4lF<dQln7UTk<<A:TO
2CoNnckIWBdC>0>XjZqc79`<k00?Jg049dfk:^?<7d>7\k:Aeib3>Xq89[fnY4q>
BObFkO$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_down_IO
// Cell Type : Primitive
// Version   : 1.4
// Revised on: 3/19 '03
///////////////////////////////////////////////
module  pullup_down_IO (io, i, e, pu, pd);

   input i, e, pu, pd;
   inout io;
   wire io1_tmp;

`protected
4IOc4SQd5DT^<gC1@:94QPP?@^^XQ]T8>Tg3WCWCa^2NV<6TbbJL0d4;7\[WC\AF
HZ9cq:XR?nj6JSF72?:<\2HbmFb91dCX;PcbopS7]f:4VOIFaKO\apme`XEnqjTk
U6?M3F@0PCd[H8alVKBSK9gdp;TO5aNVbF7iAMbjp`d<6mX=1XR_10XLREG^Gfc>
_hPm0L`mcqMDPMWf5@bY4;8INPIg;2Y6a1XZ5ap[NOKXImnAJP21EbG::P:6i\IM
`NFq64n\l[Z7a4;>2=fB6@Bj>BahQ_4@`[UP0?=Lp^2oeX>kKPYiIZGi9Z;bK=6<
ZK\1hin;B=?i`HX6\VciMohd^8dfl1<iqL3QcE6k1C_3Zki33Gd=9YeXMiYRMO1i
68l>gIii_e[p33ZVSWi2Q;gh[O]];[<R\RQ:J=m^M2gh[fXbDWD^;nX[qh6\`CZ\
53BI1M3Q7QXRFNQI9Kj7_Y6l^CBMURj[]GC9UelpgRSK0RBgG\FVPJOh9Di\8lO9
0Z48V[7>AI4FjAOgB:C`g;UdcbUdk4qV^T]ggDjkAHm846>L>YWaSj@aY8MP0:eS
0?3N>F_D<mlU:o<Weq`O:CY;cO<SDleYUeBa\aghlXe@W2JJDkNNbbL6oH;6?po\
e@VJ=[MK46IUE8nJ\]KgjPbkkYQW=le<q22NGi6kp2\3Vn48@Q`jSn2dod3;=f_m
p7a1[Z>9Q9bOK2b`7=P:>IaGq>bX;C4DM2AJCP?C17gTm;[[<_H`MaRTZ_3cVKIW
]KkGnVm?EJEa?`Yk;RoGidZcM5@KLlQp`LO8TaYpfgl:e7]8L\QSI5mU8]Gd1_LE
nN4@S\^nq50[IE>EqL0K<SG_mc_J7ckDp7fD1W3T`HMT_EO]DpC[FCYEV2lNMl_<
ZT6fIRRGXqLLUk5477;n^K17V8g3`BOP`:Sa_KFoScPJfKl58q[`^=19MeTl4QjK
El2RHel1^=S:ODhGOD2M>H:@Jj:[29>C]2>6O8p:IedW30EaRV5ghZ2;`hjV0q:K
EdJL`7I76Hi[OL85XaN`q_LFQSUjN>][J4IP;7PhpODR>j`hhP6gZNg:\Jk:3=_e
\8;2\]4qnB16`YK0McbkNA3mS9k?FcWqYB4KmFlc;c2@Sm=BOJbjJLP7Ll:gam;N
bQq1``E`AT9X05aHX2b7H]02IFlAGX_YFG^`^pd3P0UW0WNAoXl5TMlREjXn<U1C
S7S9@qDY4@h=PSVV>;lc8Hhj?R:5EZlH2oBlJb1dcnTi5Qp=0RfX@?DJ\L@Ki=LV
=LC8>WDIO<3iNimp96?a9jF5E5\SbB6^fM`5o9q230CRZogKN:][S32e;97m`jeL
TW6`XHOC;g6[?=7cKB6a>p=S_DK63>SRW2HU70GB`M11IQl5\_cMMII<EQJ7b;IH
C78c^pZb;CI\G;1GcjB>G^1R7LI@D5<[A0Q19QXVk>enM7X_0Fcn7mp=i0Je_QTh
?f4JYEmd2fGnT8JT<io=gijKO8n\NdlPgfNn0PpGJF3mO2qUAgkD2fA\<niaeKaI
\KF3H<PSCgbO<Tp<0dF?Yo_PDTbMJf`OZl0\AML[icNeEIAp7:a0FVepS3^\56_7
`a0M6?;ZUlNRUEkDn=b2K?QU2=qEVboEVnK[^06\M^@jgHd4Y>7FIZD0_=6`BZ8\
[01YlUPB623YjeR4RPpRCc;`lb[O@j6QX:A3<<qggPd^UfqZ3^<7YBn><96CXUfE
>?@;hLY`X=epQF1Pn2o]73=hX:MmEGi6:bVcHP7q>CCkG^4p`dKGNWVqSQln[`]B
`\aXB<Z<62H^[FJQn]iKaf^]`cQ=b\UB?lEYS^EKmlD^=4:p_e5gRNgVib3GdQGj
01MkAgO3UISPnfKp^G1`^fC9^?EVK?9LlgP^1PVidLgq13L9MB@pde\H=\eH[`;M
FPZ:EQ97j`EQD1L`VHGn^[DEll1JT18PWN8^MV<;]j>pD_Noj^Kq@o?[m\ceg9dc
0@mACJC\TNaBEKlq;[^8`6Zq>B57h]0pN=E6VU`qOh<kEKJLh4B0UQXRUAjpVG3\
Nc;lIBPgl>cb8B9Ci4g8l^gD@BoKgUAcYe<?Y\ZARZ0S0X0pZh[nA`ZqaJ]M<nLa
MaTKd8kZ7LLePehlij7gpH0TV:=<:45_6O3AWJQBQCT:]>[hp@`7U2Jbp]]lBalG
pN=X]h1:fgXF6;dOREMnRdW<B\dQ7RbXpHe`JE^]d<g5OCZ88]hV7P_mgnCMq?=d
R0gJp_W:Id7Xp>hT@f?V[dM2n<EpRPCI05ABU9T8mn8g@=^m:od0WVmpV;lSYPnq
n=PZ1iSq4VRnQ4npLiSaVS_hAU\md;BE>Kqa3]gVZW_Kn:oag1OjjSp;Ee`Jb1q<
W\3kkUGU5;0968<l3DE`4G60\Vp@XW];9cqQWBW9Za[4=IjLg_gJSgW<7kBmf5Kc
i?Kb1oNIKn7`o=JMbJk4=H636<3iDlaI[AJpNajV36YWaWpe4BKg`=q^Z;OXhR>X
?j>oRZV??HEHGCl2\EqK5RTAd3p<g0WZiUaFc[Ph06F@@YUaXm3faW@W`_\D:ZJH
`1fI6h<<UQm;9\[g0q;3]oZF?p9MUiiF<pT<O7ibUp8Z[mH2gnFdOgNnfBqOUZ=J
f\qK8NZgbd@bh82mcY<=_F?C^6F7LRlg`q<=Q1J:lpU3hHQ0:IOGCZNbJ>M14720
AjLk?BoGDKTgp9PH?oePKiMFikGXdk3[]6=DO0CeLK4ENk^^1?kAMQAM9`5_EkF>
k5O4DJD3j^NZh?HKU^GIq6UE5bF_2WTVLibbbZVHpX;hn]BSpm2=ldl:B8792WCU
f:TL8W15V:BpX3cWRc>qXOjU;X<8>VJ2RTTamhd<qi?W9UBiWW:Z9@Bj?0o7l<aD
E0Ye1n7WMq>QhA<0VnW5=Wd=La`ck@W9@@gG8qP[o7e\QqPGL`DQH0XiNC64KQ?<
=jE7<6<ZL2qSNQg5DCp4_j6WCnfO\VCN[h9Dm\TqBj4@9_nWj6>53UVKAnG1i5;4
a9<qnOKlKKlqNU:8GfD2NW07FNKU;oB>C=7JX:Yopi=@YW[fA7ZN:[jd]R7897]1
cdRD;=9HZg]3?acj8eTo8Hm:85@PEV_W6Pe`hcE;5B4CnQOGpE]3A]dkq4f0kZiY
FcgOL[k<XgR9hqLMcO4d62kRd?PSXhgH2WDQO1QajqTSjWBEGHo]PfZC138AR>mA
GN7?TDZ1URH^_MJ=CcGkPELU83WiF_DHWC9<c32M7Up\I?7QAImn>g7[9K?Ri35F
`ViTBeq9S`>f\Gp909RQm1qj?H1HKacKH]^XR]3g:9qOeAaheUq_fMn59=?c`l5Q
_nWCM0T[::0D1EMA09TV6MgADiog23qf[[QB=I1iNiC?Ac\^gR7WAh^aMql<fc41
>p3gRCD=h914KRXOhE^33:qOWIck>6Um@JaH;X]gd]o=c=IiSapF^g?K\R<h_:7Z
4hI;\UZ1IjEcOWiH8fqh>`2W:7pZdGfmolhFaaKFZ;kbdDEiCX76nimqD?o1b^hq
8X15;>6BeU650U4^RV2nf[R\[AWqA9\;1KQ?7bTO`famkJlOpm1akSWH>mI[D;l@
QUmjGCKkJag4qE\E;3Fbqf3AhcCHOc5J;YOAI=9RRLHBFPX[^ql?182g7pQF;;T:
oc?K<[N>@1e5>dq[3FNZ>=N?W19b^o;DGe26>YURhmq]Km=d5^JlG5m\<:SIKBiI
?6Zo?7pILLM7VGpF5KV[<>e1F`Q?^S8p@148MZ1p\ika7@;TJ8GR3mlN28pj7ZAl
<QIUXC;IO8oNW]q8MMHDi=q0VgkEhqiH;Q]4CpFFdaoAL<D?ML;a<Bc1N:]Zf2NU
985U?XE9\]D_0[XBH1p`P85f_K>@gqGYOV_9Jq2LZb9N^PPmjHmNF5`EMhbhafD@
CplS]^W6XqKIb3W]>qZ8n]`Uaqjfj_lbj??D;7g4M;?2nkaOSDLXJZSbfdT\Mbjc
qVSTZ>_dqN@2[bN`CC>FWTbach_6^VgMQ36dMV0W>MidqX>l9ZE651^MlJ]K]EJ9
e1MebDMKY45qGjN2R\\c3c@TdnEoCM??q@bP<OVF=MFD[?1GRK_1;0Gj:F32D[VT
dPU9RGJFfUN4\PLYl[bdMLNX9m1933MGp?mKd[47jU<mgNG>YZbX@pNiD11_Npc7
m1nCDF=SQTGl7_=jih4fbKpZEfZ^F\2WQkZ;\CiAR\Hn_K9iIqVVh^3^N280<^1B
EHS6nqiHdfY4<2`IDB6?@=]^Nbom7T8ZJFL7GO`6@qCI_\Bm5pf4eHe\9UV;lZ?N
VOWISeeHEjq9iP@\j^;50?:HH?lo:<pRMPH1?eY@_IeIfNPRA>;OXe3GVEIkdkG4
I`q`]co?`fp1WBY4X\=1L]BA?nbUJ3768]OiYESLMmRcY4@QibkPDmR]9JhG\[l`
XJTn^pPd1eo4m$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_down_IO_IEO
// Cell Type : Primitive
// Version   : 1.2
// Revised on: 11/18 '03
///////////////////////////////////////////////
module  pullup_down_IO_IEO (io, o, i, e, ie, pu, pd);

   input i, e, ie, pu, pd;
   inout io; 
   output o;
   wire io1_tmp;

`protected
M[]1>SQ:5DT^<h=`7mfV^np;OQGZM?2HbJQUH3;\CaZ2lKdIo3WUZ3Q25nWRo^E6
[C0^;oNiY2a<E`N40P\TnkdR_;=;gq6fdMH\4gWS9W>I@MolP^:9Hi63n]hH_YSX
QI3f4pQ22oaDq1eI4kAVgN_\_3jY_;HoEXR=MIhVqdKc0fEZqFWU6:LJEQ1>Le1m
6Oh0k267p77:W]ZifU?Ln[Q462MM6i37pX:X<j?SpeJ2Z2P]>MYAG:Ughfbl6eJo
BTF28cR_^B9O@=A^60bY1kf^jLK`q:_kiTa<iN[mb9mhU2HH;SF@2eK4;DXNDpFB
_MmOnp=;AA728bBOSSK<bpBk6bK[W99N6<@0;_M;A:fW^TJ9Fq1IDHn?2@9;N_G7
>BFdWm4J7EN9TgEAUq1S:gR3Em0Nk5V_U?EmLgbiKMmWbe:Vid^V[kHWZN0>_JQ1
G4idIS47p7Jl_6UPnZX2DP?=jJ1NPpGC`<VVUNi?Yhhja8B[obD9qTY>fbOYc7Yc
U?]hilmhdR`p4;DBUMU@@]92GjF0^=5iB]0RZRk9UfULPk?_FH<S>9dU@B[>l53f
Q4:oq>`0g_4a<;^:Td_2RmH^q]GHT4@fUBigT8]6TaG59QSj3mRNDa>p^NDaKKVW
52caoJ;71=X0qW[IYO47XV53;BbT]XTEdpjFDgR57DCkmP^K0jmZAcf31eR63`B^
bplaAO6aB7[WhSB=9B<A^JTNJ^TT]kLBq\EH>l57o5]F3gf`F8O0FK13D]a8]>;L
]V^p>jAJC\eLS<YU9m8E^bmgfadJbQk80XR796q<JlVMEl10@@BQVg<ToST_Ddb3
HNNiPjqX^3BXTQQEce81dM\\DLHM:8Pl44@UOJ5]cpRiF@NVF2UZ]f?o[nAGOYJQ
W6HJ[UjS0Sn`SPX1EWac;m=5LqYclUO:92@Sf2=lVI^4b]qSX01ElBS4@O[BPko]
`NBLUg6W\ca2_^5=\chV>>hq]Y3hF;<CiKD6ndHaf1EBIEQ=C0R4Dd9_p:UiblOb
e6oS[ZTn9HAo<P0669fj\EFYZY\bp]b6en^QF`0WFK7SGPN]O5oD>koZ`30=>M1k
Sg>35=MSA>>qh`4<YZh3W4WR4_1;\\Aqd8:HPHl275:@]\a`EO]366^b8M1UmUE[
1=R63fo`YfMOSa9pJLPif8bl5>:h?DEPQX]X?:;8a:H3eX9J1kAiL1VmB^a9LKQ9
pC7j<A;pN?TD9RbfUX8hlU>Po:U5gVJB`HF5IW]edIiSG^73qm2K]CSnhH`TPOjS
dk=72>```:\7g`^:8:JbAJ:6Sp[b_5PP@X\V=1R=Cl4X_9HC2WSf97@RNYl<E2WX
nH<3;qj^gcPjJGWGKL9d7ESLS^>T0Kh@oF66=2VWkSfC\3;lMgB]01qNaILmm?7Y
5BfAlBafHl3^=Jh87a;a:UfSX[Q[iLm:4]fGNiVn?=@78WBPlEhmT39nQ8pg=LZ2
n^p58C27S3;JWP`V:I`JF>0CjDff]@>=O8:p1R2bnF2R_mjaUkj=I<0ESL^>Vk]>
S3FW0Rq@bW]nZOpf`2==JGD5=j]^0GKnAQVpIn6`G4k:X]^InFO1Y0K7WkahM=p>
RbAjdoak5=PhF0@poTe0@YNq0VOf?QCAFU]FTgTn=V1cm<mDcm9C^jR]F6q2=De7
DBqF_b\VP;MhW^IB?Jo:P2_PZaL;0Ale3O3PoSkonPA@Xk0]Sp5mJMZUBTQUjKBO
NS4aL4\\IoEWTqLU3`i4`aZHU1JTaRMR`k=U3kVk7Gq7MdnJHjq4K_3OB6IQ;3]Q
FKJkN47ZDhIC^[iN5da2eXaSP=INbB:2bebi1J`m_U_H:LBTiCZN@KP`@qZSi9QP
Sq=Xk_P@7S>YMDU^c1bo_BKFWHmA53BCGjqOVNoKaZqRYd7Zc9jC_Jg[;oU754<C
:bkOVf?qh0FeOfQgMDPW_4OT;=?lg@RHFkSSPBA2hXM5K>2mc7HhVcRmpH4A6Bn0
qT9GIXZaqo??_@:Ip1`m_W8[M^Y7NkldPHXGEB8GPWnjIqF@Z\Ec1qe\c7Q_RqT0
ARefb[GHi[o?OQd2M9@o<eg_WGkW`aIJ^W38M=fW>n^mH4jCSLEg7SPRhH7Y8amn
ZPI?Wp]]1m8DCp_BIJ\FEZ?4hS1Ui9X=^:K9Z4]X6MeZn5^Q`cpMH^\YBM0GGbC9
OMZIkckaQDC^DoMp1an:S^@q];1[S\dFJ=XhLVkb4]If>iH>B3MJqHn7]Um4qDIk
8MC^X<ZAeP?fJZYm<GNdlGW5aimN1kU=\a8BaZYH<UkhjpfODVeQdEHI9[2PW[qH
ImVNiSpMSTGDbVMHoY=6Jj0XnK_h;bhA[g:qk3FkS84pSN\fO5dK7XQ=YJBVU3L^
_OfZ`6O6<8qISb]fFDF2AqOSYLD25pjUWOKW3n2MVNRQ09mj3EVD?NF3c8qdLU^l
?hq9JPo\N]qd\nBcOhY`_XY^XeBX]B1QV`h2e:Z?Hoog]WdjDDK_VCK[0j0cDTdG
Uo=j:n]qlVQNhhJqa;8knQWqA@OiS;PV9L[nP2LHdZWd=\E;`\\j]]:?I]AR9GC`
Y6GlUOHjo8eg2JmXL7iPq^IMW:2LpHKjORUnR]IC=^kDSUB7:QJ\8QjXP;\_ponW
D>O\bQ9;fWQ\H?9`j7KiRIBONK39\qD5Jo`e4p@DNm8go1;ZR3KdHLi1:gN@=Df5
R2;o>\X]AqF4aah``1?5gmLS`p0Qn\OR4l\QPj\XYg[SQp]@TBgaZpoiIlOH6>ZA
bH\[lD7AZ8clk;9K90pT]feJl]3J8`@8cULg4[C__g5L_Wp=37e<gPpeJd2BcLq[
gKA2iD<_din7gk6ha8?<;^jp1^4Y=52:KG@lo2e_l7]YOG[27cCQnN`pV1SVIKmQ
600;IEFa^7fCb?HWoTBqFT:T:5=pKmRD1;kq7W3QQXXR=?MY<5Cn9Xm[k_65TgUj
9B][elXopHV[GilF9m\N7iBkQ?Dbo9;4;5mnq2YH`gJTpPlL>h`:qDZSNEH?B@K;
`Ml7X]IfeHWNA7XWCgCKqSce2ed[qbF[15m]?S128?^AbQknqONaBHbBq@:HENGd
OPaB4Jaf^kFD@37f?4]akYhORkhqXD?TbemqiUIehMME1;R[03>OoWYMR3UgWl_`
pB:d9OR2O3450WC2=D[K<K<IRF>aqD;<Z19XpdBloMScWSW@3ZQK1QNSN^A4K_kR
f@amAH;[`l<o?2J\G7ZJ\q2Id;3KUq2Q:okF0415Pf`MFoLOC6OP3`Gg<>@imqK`
mdHJXLP;C\BNGh]InDiH\Y]Y[p@DJ;W[Ipc6o>6n?3n;D7LKieT;0[`S5Cd[^qd;
E_b\^pRh?]LU>?LLnm_@ee[Y?]PdJAl@@pCK^ICl3pJCn`]0Wq8F?__i^qjme1_W
Pk\X0e[lELE[]Og_Y?VRg^\dIg@X>c^`[:]OdnKi34H09cW0@B>6PO4Rf4bL4_pk
[66Z8b94Z^OMo4HhDbK322=Y]GQ13VIX7J?pC@F?L``>I=gV]]g:g1XmFnIjXUhp
=SE8oU7p^9UKmhe4`ZQ`O<;@li2jj6E8Ef0p?^UZJ_;q;WiQ=SIoREkPOShqQN:k
U3W9;?m?A>jB81pbmT;TCPT@3W5:7JgbmlpP5Te]lXpbF`BOlf6@bCWEL^GMZo[E
Y>?lF3pOZbO8D]p^L<:?g;I?7pXZ4DT]`cXi0_AQ@O2Jan:RS[O0]36TPNAZVMRj
5F;DSop^AA;iG4pN]PQgo>o9dIL<G@PjgggYEmfiQGqHmB3<2Gq7;6X9aDeDRj0N
DAT=\GB9160Y<FZ2dgaI:Pa=a2NjSLYT^8pkJ3XYmUq5Y58[d<pKmG\?K1qOgJ28
>IR7fh63P]ekmmm3gPYkkCd`4P3BI2oCXkNjHeD:ggg`M<=f\pk?@Am9iSKBG]P8
mgqFQW=bBYq>YIgBiee?BM0k[HnZ[HUKoQS7V=d6Nq>\689FSQ7E5EnTXbNR\[XU
1nA3ODHW7k^LGe?\I6fh^GPM\eXO2h0g`:3THE2ER\EeqdR8CgVKp\>mAj>Rd0Uc
?Zj>mo^GWA>TYU];E5kFOLM<p<[oeVj]RB;ZSEUg>\c6qJ76bio1p7d5R`fn0oB1
]]kk3nMn<]_9F9Rq0hFCna4qK9oUnG3LAT]H9@QES\VMqIje]K0HC[fVKlh]Y_Zc
Lk@PZIGFGkTIBJ7C`P_Ad]d\ON;=VGRRN67S8SHa2Mm3AO_PY[Iq6>BD_hd0MBSD
Oj^9X[:==Rf9JZ7q9eQXK^6qPAnC@N6V\DDTSGN:[M\WmD;Q9@\dq^M<0@dfqbVn
7^iK:^:maW0I@:c;Kqc`N]P`Pg@1^@HG61g0oViSMBVkjq4o50FXgq78AX<m\Sm1
SJR0o<_3FR[AH_U<CZqL^ZGHnKqYnP;XDHb]Un\P?1H6Ri1Qa4fT:kfkE9CnfLVN
1m;TEXUXdEPnVeW:o5m;:kQqLCS\mVOCbcT^QBihj7^jqU?f^ZfGP9jWT6GGC\P1
H7neD=D3pf39g;3GcF5]eHZc[g6J>V\@[[K2qDN<8[dNq@bG84X2pifbE@Q34a3c
8cR5h`Q3pC_[ngHO1dlfE9:;GDDN0n=J0nD\cS^RI\0A;5e\V@Z``8lp:f8LUNTq
ThcH^<GX<FAlnR^1V>bX2kLF:Z6D9NAT@XpAgdH0k>qPOAL2h;kEk0ZT]nA`kIkH
g8hNQkS88^eMJnVYBVE[eN>KXAH^M?N4R3HO`j4F@3D7Enq9KM:4Mkj>2X;JLNG5
AniF@M:<1pG89VgbDpWMc6Y2XZeT7iW501eD0Tq__WS]QID>IcmlQ@M:66]?]l3?
c:plVL]eL>pEYB;YGdgGB7\^aIdIjD9ePJe`eMCp9SgK;HHDdU[^lWJT^^OJNO8n
0SKFPm@2?dU0lMAoFX<i68kUk7oKk;=qa]S=hj3q[Qn2:N[eTCXCkCC8MDNgpW70
<BN>>0Jm6\Qn[N?OG[1\B0;cpiT6^ILZqXLfSCamd`6YL`TFJHCSBc8iH5d3np7m
mTc`mpVm42ES2H1lo9GFP9>9d<pocNaF;44EY@Z\a<VmAnnW6FRGAEp61Q9QTRbd
gc^I<SMDQ@gRTJ29DeUoA:<9c3:I>g8m\A1]Iqk5nP6n:A=IZfOm^@LPdmVGm>`k
2qZ3L3Re8q6[c@eXjqWT39\g07^N^SJT`2HJ[UjS0Sn`SPRUInaNoEq\8mY7=KnC
Ro25868d;F=hYXE@T@q=>KcghFpB[ca:JCL;\WES1=0FlWcajk:FGPp1_KAlZTqR
WSPm^did]d7U80Ia?pl1UBWS9SiEjNlQNh>@:ND:52Lb7c]19CE8bDAGcbQ16:p>
FmWSL5KEJaX52fBS;=p=La9E4Cp5JQdQmp>BMUcm=pRYb;cP?eE6q29W02\Tqi@S
ea<P0IN>Z_RcELH>`RjCX9cWp1=I[KhCq^E`^7LL7Pmd<:@CVi_`pN9XOLD]qf=N
TZHZqb]@`m>gqBI^BN3>RP_4_1:KLRCL0:N^UKb=70GR9TXUq]b0ggbQi]ZQ<O\J
WV>O_<ioWAJVFPIp3B0?i<JHS]^n8=?K26Cip=0cmXVce=J2XCn6@6dWlpEPSbVj
oq[F8Q0WamDJP@iVH5X\J0N\`lSMd[b<q;cRBCgLkFc>\L?AN=WEn5ji2BkORh^n
ET2a]qDW6ESY]j8\6ogN::E@3SfIJ_?X`k\[BpI?OVRElTUlO[^T8d@A\;KCpFSV
BQNDU<HOS>b^7XBcF3Kp\NKOiCCqkfZkZb48k59U:9_kNgU0XQCiqCY\PCHFHVTJ
[P[HgH62qm24Mk2CYX=CcOaSX[4o_iL\onnoI6@\J^o]pegWH_N30ojPKh`>>q>X
6SIEapf8I2P`=Uj^GNmeUE_9CN1Fc\=ApWmV^eCb<^4B79fcAlbVUpgimcmZ3oIX
@AfMC6<NoMcKcAJa1i]BSJC6F9qGUj<G3SpTof3VGi834lGg9__F[j8qoHJ1[iJc
MQXY@cjAkeUff_=aqKUl0;AFSmHcE^g9kQLGqI3oYclYkY=BGdmZ3bn3\M>VZ16d
fbV_N;3Ap9SUkolgp0D<^_ZW`<n6joNHZYlZlPI@66Mp106K1_^Rhh2emOdVe4>o
p^GU=FME960o]Z?g`?jZQYI?LKZP6:d`4l51^q0WKSkAQHbb?nE4i8hLiLg?qnNH
lGcipFSjEWOj$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_down_IO_PSCN
// Cell Type : Primitive
// Version   : 1.4
// Revised on: 3/19 '03
///////////////////////////////////////////////
module  pullup_down_IO_PSCN (o, io, i, e, pu, pd, pscn, ieb);

   input i, e, pu, pd, pscn, ieb;
   inout io;
   output o;
   wire io1_tmp;

`protected
NZ>B]SQ:5DT^<N=]]m`2<@=Z5[ghAh0^F14pQI3DnXRiUC1OaibWYiIAAnRn7M2I
pSBZU8;6C?a8o2hQ_]kp9_MA`Kqa_2:EHS^]D:\eHS]BTQNh\K=?SEpPQfQLlObS
BFS09Pp^ROGO40RSb`aoP2j9\>6h=Cg89@\=:qb]8LmEQhMIU_eLDkBoiAi9=@XM
U@gQ:SMC^PE?qV]J=Kgei_CR6g0iJaaeUU>i;g^;So:PD^T9:_L_qIiL29cZOaVD
f6KlBF9fS_:Q9`^jd6bV?8VjjBe24hcf?HVi?U6<pJebM0gQajK?1Ld45XNn2g[K
Y6V5=\70Ye<iaWE`qhN\k7N=NRW?1fLl>l_Gj[cg[M@dAdNWATUo:eljq=WNBP<`
b_SiKLLB7;EPF`K`b1@SU9k3Mpl=FmHiGJCO6T>@^hg`D7FTAfL5bQWidm0g5jo\
dgX9^p^M<<W]m121HSLEiE^lf8H9S:\D8ZWnh^S>SIa8^bZom`jT<pL;NcRNXjgM
GPC=bYLeCSNDLAfijH3Cn`8Bqe8H7NJife6iC<^h4fXl5>`kR?hZ:J`cBE2po58L
ENfj\<Ra=CJYEiG7Q7_5B;KO]NTA0_5Bp]O8<cV:>AE6>_0RZ?WY5[W>^Qh<>NaQ
4Egb7A>LImlq`]1AhkQ<YKHTOF6M\8nG<MD^K7I1ZZW6GV=`fMESXTTmq^gEcSho
VOJNge^8L6\UKCf<TaWU0h8=<53Y>E>f56WdOaRpNOgR\a>?TBFO\A`NpF_o:IX]
AEc_`dgdV?MgJ`c`@m5_NY;AcoeRo9e^DPb^INYBWhK48Bcqmb0fAW4iJ54_KZ:C
Cm<>SRV@;9hcF<C\[ECeD=Wb1:ip7O4P\PH25K`Bgf[7FE3Q\DL72>kEj2m@ebpD
AEW=[0nbXUFb\NPdJ:W>\G6]WZ5f]klMHn:?2`h=7mQ5>bc\37ImXKU?7_aq?_QD
64c1HG8lE@GFKO9?1=55VIf[e@FKQgQg>QPp0>41IkL?Z[8UW_DO13lGLCCZBE8l
FSZ>ee`4K;`@0J_4qlTmk`Wq?OKAK]VpKc43@FI1a[bG[^n17e0`Jb>qgn:i1Qln
:OaRQ[4[cOmg8O<pRH?c\ZRb4C@\iUP]5VkM7KjagRIbngM7:JEaq1QJVX8:p=SJ
?@@^4co_RbMH[gELTG>LDja2KXVE4p6HAe4^Hp3gbKLS>`0>;Y]e1pk>cSXi7g;l
oVZ=[`qWF>mb\iIGI5_qY1J[`gD4V7hB=YW`Uh45JQQ?_QfRLPEWjnHGHB`pWhaC
Vi;\n5VDB\No;4cKPb8qlUG@_i>Ni8R?Y=]NKbdBm1SUhQZK[_i`2]Fmo59p34j`
3fjS`N6dA]delI6l[`qXgRl;VlGYoeL1=IFK8oMGYp98IPaX@oli7HKV0i;6aqFS
oWI50CN9kRbOj9NBV[[^;=\N@?NEphKRD26GAf3nW@Z70OnaMblV0>Qc\>bU>HAp
Yc[;SXVTI8KlG85X<KmjjNmf]ZXV6jD_EkG0V?<kb0a2LFEdcf`UADnCAcDMS[e5
aT2fK4nGpgbS1nXCKVieVgi<D[MY5@hAeQ=m9e=0d]MpJYfJ5=;<4GBH8E1ZH@MN
FlV3WSS[2;8pCfbGo82onSWWL=gg_`knibbiiagQg0RXj4:c>^3ph`G^Wm0nX8N?
CB5hMS?o_aKMaTLYf^JB8m0g_HF8;[NF?=1@KU\ip\PQ5ZleCe0EPNS76:5ZW:Y6
<_mGCnMJ_Hl@]@HKa@dpce]j3kg4KQehhl]jk5F3mgg0E;ZMF`hPEYqZI0M6Lnnn
9J9:D=lGEb0J0Ke=U0>eQMV:U03OB]2SE7=>`pE10bE5?GNjPAf9EL9\Y@I>VP>0
SkkfD957GQTPP^9]S]Kl[qLJ346oA[R?VD]P\GeaTIo>:6`?f0MCPPPGFBY>:BOf
117I0q`jU<8R;nbHFIB4X9nl3TTQJm\WP9EiKdg4_H4E0iZOXPJPDGpC_Od?eW>j
30TPf@[QK>IaVKDTcLPCfWXhGU^K_g:GNi8nYHjR:l1mHTQD0;S9V5n6h3RnLnK^
aaE]YYQqCZY5U\?q[K83X0m]l3cHS9Mo8BM@@McGQUm`J@5_Jid4p5S;f^09j\g9
n^>dQMgKTU=7qfe=faVhpZPefZWn_LHbaoO_Z@?cSlHRJ5dlg4EB?T10GAH;MT`?
hD[o\=P<YOWdf=[MWc][`o@epVEXNB54A?a;SOQT:V[<BAIclTNlp;ROIQhjpR3I
JUNEKndZaJ@=C^_[Znkf:H^P9lT9\L[H9nlW0k[8CO7Rm_M8:H:9CQofkDGIqV0S
5cQc0j^6>OL8]lZCH28[@4cZXaf<\mPgqm0?XT=XqeekmU6C=`@gedc@N0INaMQX
C][Em`=BqOHdRX4aBh0EX1Q\diBKKoOTgU2<_]1M9W7>cqS9HE2Chp5I:`d;6jhD
R4GU30@c]B0aO7>RgdpoIG1\gCIQTRSBhR4BKC2kO@Ag=4q:S@AeJ:p[UnkLojJf
jYJZ3a364MeiL0=>ei@eWeF7iAIIk_^;YZAkjPgO4WQFWG`eOq>g7<TAgp_c0CJN
VF;SekMKYeaLT16Zl`V0XLHPbpNPBYDi?nkFLI1]27CLZm1GA:90AqCid5al4pOW
mj=NbpI18jU5eQ:MNn[Nl==_dK6nNU:D<p2k2cIh8pf=7oi:gpjQ2]@29^OEABSQ
bhnadb9dEpF\akcG[p93B8?UOqT0e\d^Pp^o=63n8<djnk]TJnL>_HBUhD2^0QRC
Z94g`GNJoODQ7qYLYGlG3gVE4<:jPkGdBTcbdAhR=iWK<0q=bX81L>qUl]R1cLGi
4e_<6<P\W2S`21g]okR9OIUDIlh;RaT5<_]ln>pXJZ48o3[2>Kb81eCa6P`q>[G^
S@7Bm\L6[L0>QOd@m20h?VabjYpVL349mJpYk1A6EMR12A9Pf@?aQ@lEafY_fC]p
BBlP3eS6f1VfPaj14@HS4eGi\XJqh<>V8YJq9FdE?V6p2ZMoEmmPanLl4d]Y6cdg
=lM6]9UkF7lp_kJ74b;9:B8[XfG:NEnaF7;cX?PpCIbT_BXq>J>UfD`p:N>8^iaB
\Y:K6OU7^mAK:777@>3A=>kABUhk6`o9Qg2?A]1[\X<Rg0eA0nImdSCRdMUp^Ykj
?iHT6TE5JM6gLUDh>8j0?4HqCfL>DAGqQR]`XL3qd@hoI62q27kaZJ@RFG<cCc5]
?cn2bY7T6:GMIYec8e]I3U`q8?9Lc95if6jjU<28F^bXpe`6?GjDp0cSohme\DQY
`18jl1CgmeWNnVL:Xq5?D[:5Sa_VYF21AfHfaeKL3ETmeq9gESYJ;pW2lbP`Qq:C
PD5U1Kdk\54R];LM`YdeA6e3e1b5Gq\II3;\h2F6P<EYW5=W_TcmF__nnW>5OK]<
J4<S@EEfI>kQ39XPk>ccIKK;M^9ElCPlVpJ]LnE;VJZM[o8XMHG\[F]@^3MObq3S
=3oi<p2[ha]SIqj`WgL_XVoDObC4kj0S3^05T;h@_pLKDlQ:2qe6a?HG?ZRYUf8>
4T@`Z_R=p@L=n0f>p6dV=ZGHpc]jOIgRlj6bPCm=fH_0pa@34?=SWU4bQK_33JLb
<q9A\5l3:SC4beke:NB7Eio6O>JR6gPl;W[5p<Y15;THpKHnB64j[DEkB:K3YNM4
9;bBO\LBq122lfM[q\E;aNA07mmq4=02R71qMk33dBW^2k=]14Sf4[kn4>=o>>H:
H52?8fV9gch?S1o7FapmLU0NcIPfPRL_Eb[Y9Ri<^:3IY6plVej@ZmpJ@o6oU7p`
Tl7lgQqMe^VSBGq0cCPSI_pYYBJ7<KXi]=[0Qjgq8_AVFH^qG_g7`LY[00]fnT;g
feO5d[q]28?@TG8D[2c4OQ`WK?;3IUAf55Mcn65eDB>q?Tmm]6^qn>m3[C2=6cnF
O9O^g_^7B\P:B]MPqLoXFSS\qdQ^g[Y=^YoTgdQ`>:2WRp6=3PkGlDDVD8]K2^GK
PjE@mB5]Ip^M3@jElUD?YP@L=F2kkAYkgOqY@6H0a7q:RA\QjVhXmoTKb^^m`I[=
WG>KeeVQEjp^HTFiFGqhVWD^C_od_OV5fCO^X4ipXHeA7L4A]3T7SkZJ1^G;IIYm
fG8j[:2nWFM_Z79qS>MSadFXYL8VBClleNWd\jlk[UYqTG>\UL`q5_j1@OSVgUMN
G<S:n9Pa>k@5\I99pM8[49_hpQ?X6AL^6<n0]K1Z=[KAa8]`;:395Z<^;]C7UT`g
7:kS<qiFNmXnlP9lSYXP2SH7TWqD?i2M:jZgOWg1i2<ffU?4l?QLaWpiA<4<^Rgl
DKQneOEICNNYnXCbFZqW>4X6mUq@9<1?:iq:O0LZ7ipN8CUlc_fg=P;mZl@po_:^
9i3p9d4K^k;42An8onN=Kh<oDid^Q[jnOepET>oAgipYY0oMeMmiL0bNQFfGN:MG
9dZW[Z<]118hVYYJUm]LBD9j31qi_]n11i8H=]kc_Z228jHphGW]k>]pVF:?kKl`
1:baFen9O<9G8eY]PdqgCiIdZmp;<V\boCALon=:iid<\V3S4ff>JJ^:CM@6Hgi8
]B<^]oAcE]oB?I?fgM3Oe5XFRhcEXW9m[qo<>:@Q2QWF>E;5VULb`=pS81f;3ThV
5PhIVET5g[^i@DRm=\p_d653a<p5l3;m^iF:nYaDUQ0N@ihd59?0BgKq>Ah7k6]q
R;1]4:oRGkSb0dCC`Dj=poRXTM:QE;GKV2:7PhH06=4_QImGkUaPWO=:ae5H1RKE
aOdI?2DEDm<n8:?5qUaXK7ZbT=^G]6;L21X<LCneRliGp6De<9FPq@[;0HE4\jG8
ic[:_AZBL]7:2cV[`qXK41<KGqlmXSQY:@bH<8P_oZ=cCKq;gWQK1j0eM:l1L78J
Fg9HTMd[djqWCn=REa>[h=o8RTbU0Gba_DXQ]gp_CgY?Sd`^:kFIZ6LVF`1j\iNK
6qYU4fNAXqhZ`c9d>q@;ITcfm6[eT;KX;Yg0D4pDUnCl9lq5Z=^<ing^4Qm2=1J5
aBL[QXQoHq2G@>\1I91L688YU\71B>oYSgcMOR8WF_n7:jjD4EYGT0ZCWC_FZhH1
pQZ=R<6bqH:M1O;TI?aC?iMPMC\QZpWHKK73IaOjj94S:R@J@b6c8d9Q<p8>IUKK
cpSh5[XKmGURj];i5PF<H0j^^WOi:Api;;b9E`p];c9@DGSo=@@UkINKXb6pKc[S
f?]2B:gDb1j2;M0Tb4lCga=plke50:Jq3AJ<R?Y=gZPNXH6@ki4`diRNaY2qAKgk
e?mOMJH\giR5^k4^?JB5ce0Vp`V4AZZ:pPQB>ARa>ocLRFY[@O>WopQ3^HROfjnl
k?lJWSnZa7^JYVFNZqKUPOe2Q9_V=cYb]=0FDH\Pd=h[8q7D`b86[qA5COD5NpL6
fW>9;>VRUPJIEEjm[qm<PJL6XB^fB3_d2PH@XFMaV]ehE98?YO=KU0QoG><WJ\kC
l\A?R5^ZH>qfE?mPL65g8mge94NDU\@pIn`n59Jp0gOI9]p@6b2P^gq7>S5hm`P4
f^RJKZS\=;N@[ZY2>0cWN8f6ZfJ:7Ei9gJEWP7Q6[BA28B;lVKbW0_2qcSLI45o9
`mq\3h]de^p2<:eai>S3TUmbM9j_XYT0aWfa25q3nh9G`7pDO;1igjqk[]oIgG<N
2LPA;K:<b04MYpl;1g2X1pAQ6OU1aq8OHFOETqf8j2cYmR:4PVIcK6hXNhU4S6Kg
J41HTe;28qX27V<\linm:VY1lTZINjdD<nU@@U^npNF_oJW7F\DhHkJ@j;83FqRE
^0kY<i@S0Fh74oEndNO=f]WKQOMRTNRIV_J?\WA@98^c?l1PIQ:F:DZYpD;B1A_o
0hOF`]8YMG<QQpE3^42nhqlF1a?d6C0CZh`]cVXlKidCZ;pm[Bj@k0k;TRVo@mQC
Q@qdXbFKZam6R4cA0KoPX9ZW=A1coUoKYJ;[9MpiC9`EW[i>5njbl19dA0I4]HdB
g_B_]<b[1FEJ6mBJ;d[F6pb_c[iRMpoNL_=7Gi>FQncn]@okSG1Ed6q`dIQ2X?eZ
WEoM`mDGcWp4O:C6?L@Xg_Y]TK4<Uj[hW?XWa@BL12C:a0p_Dc3bNEMZB@S2BN40
F\0h6^Li<0F6WqUJBf<fmq>>>f@G[$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_down_ene_IO
// Cell Type : Primitive
// Version   : 1.2
// Revised on: 3/19 '03
///////////////////////////////////////////////
module  pullup_down_ene_IO (io, i, e, ne, pu, pd);

   input i, e, ne, pu, pd;
   inout io;

`protected
XZAoRSQV5DT^<?QiQ>N382C?VK]53ZfBhDF1K0<PX\i??YRIq3lD_K\4OPBMLYJ6
IK7OJ0lb>;UcY[cqb<cf1\<C69AUS39_JcqPkFmAPpGZiU\VXJZQQik3?9jgMeNf
kl]mHqKn]RNLApR1@h;oj]a2Blb>FUaR8iY`EJpPjVka;I@26YRfDe:6fU:Ua7q2
c`ln6VXp3APgkDF;Z\ndUP;PNEb2OiH;\kS]ndBlq]IG9bNj?<:<SB?I[9[5MNEn
gW7B6;VYG2DG?Gmqk4dXG0d`p0MdiKYqAl8DUaW7Zg_YJGJpgkdjJ:c<QiT8`]?k
qi<1NmioS4UiG6QAdq2F\MEA7PW2YLk8POi32kFn@@OU5`SJ]H>_=:X1oaNDiT@1
j8l7q7?6CFNKR1XeTGMhKi[b9T:qj[VC;=qNVPld3l@0oj4Yi2cACh\WIq56IkTT
IgIAWg>^=p?T2XkAI\b3dcL:oX@:SqK2ciN]om\;n[I1]Wl>LeB^la40M@G`p_O]
Wj2qRSK50J:BH7YcJ?7G`cZQWn<WSE607gl]bnqT?;^fockDH\@g5VhPg8n2iZ6c
`cXC7LB`>qAPYkD9;XM>MMD<Pe<GYV4@VFAc3303f2nCCb=i6WO[aPZI4]HSJ`^R
91b456GAeWE:p`^o>hZB7_Pi`U52;S`[59]N17YG6nHnpJPL65CeiAfJ<?UWTcW1
iLo>m]IM49<WYYbqe134QCqVJf>K[<nBagF^[nE<];:9jF30@d2]G3NZ^\@1U1Ep
=W3j01YiRAZYOFe\g@E8B[`NJIAB=k`N[\b^MUS8\D`ec37];O^pLbL1;Z6E0OkY
Man1^Q>5p?=34:AaCZ0GDCVd36AhQ4oH4XOXajc=W@MZ=4XTE^G<a[W3pVX^3jYH
PZ1?5I^0Zo>k9`]c\HZMl[3GeKHKOd?EA3@9]JXOLpmO@G::qS0?3kj:_]@VFoCk
P>0[B5a>dkUnkEf[BM_ch;6moU3mah1jpZ`17=DHbWHi^Xc\coWq?DJ:^gHpCA:_
9h`U10l6a5A]TAJ_f1<LS1L\\j=p]4W>a6W;;kadLMoX9Gamf:;6DkdhYn9mqf1h
oHB[Le]N;WPO[=IF?87epoP;<MHLpXba2n4QZ27LB7@8gAbc<oTcOkjkdFM[3>Bq
cZPf8odff=N`0MB<YJTpMOXmPB=qWlm_]M;@1fb2Ke8We]b^MVJiI0l`pnY157DF
ZD?6^]1m2E5`8MW4UP]dplNQ>54gq48CaATiqBNNNW=NG5ck7IXVWdd6[4gSKX9J
SZe9A@4YnekB>>DH>EkC_]fhGDlj7pe2=6Ph@l]VdUPCA8H5ge\?_1HUi1m[^qDF
cg76gce`>TBQ4h=fcI4iloVQJp[]1mA:nq6FUDi=9p=CFbN[;bC]kEWBEF?B1K?Y
nYZ_hpWi6b;LWplYfb8jX4\d:NVC=?Fm9e?Y?8h2Dcm;ZFMeDqUf_RZD2qKnm[_N
gpXXmA^44\IT;X?6HjmPGpEOJDGETq6ZI243>[_bo]>^2amZalM`DBc8]]pi=:]Z
D]@^^1;[3`CGQ6]2bH^3ZHD[FUKlQgCk;n:0O3BpPQf`<aMnI_5f?o[Lo7=a:VdC
DPfph>]<KYmq[6WT;_lp8aUgOjKkaRR;SZRn9@3]KdIHPR8QfWaq@GPBU>F^VbDI
QOBN9lEpf7[U>=IAiNiC=J]7=0kDPaWKkUZq1\FbBL>qRKO3nbFqVGM^7HLDB;^H
XYA0WVHO=:c_Akk:LF3Q44<J?SkKVSOp[IPR\ZnoZYPHQcOI>7T=IUkRHCfp?m\]
Rn[pGj>jfO>qIH\c2Ncq2SEK4;JhZ[UK1YcVU?M9>[NLA1fl4@Y6B<AdSnq6V[_o
h<JF`i8niI[kCq[4MKh4]=<\>DD^G5XZ=p?<S8bn<q9D2[IDVK]inB0FSMJX;^MN
:X7HVo7[`caDMRJ6pfD:;TgSlO0:oRbP87Bo]0CJh@70qbW>2\@Eph\_TJb8hlJq
2R31Rm<qH\9XjDE>7D[5LX22:cZ1kBJI9fXq:FF[88\8^bcOG@C\YQ\]4Z@ZQ\kk
YilYCEgPq;Ckj7mXp05^3eYGqgeg=k_GpENoO4k>pDM3H<EEBVELQj[8Epe4\BB0
hWZ^IcJWYFZ<<MLk:]8<^Gi7mp[<g0li=pPE7lk4=W[XiUFR_bC>b7o?Uo:oeBin
q`^5Zk8apBiZfJFEWjIj;m3em9haiD7R[?O=T\:49cNqEC=:3o^XN^ZRaRMBTU>p
a2L_6fA0B2i3_RgN<Ggn7JDOqAOBBXYaqG346737GCEoYQa:ZXimZWS0Ej1qUl`0
E7>p]O?R]WPGXe::I[::hm`Fq5`ABGIe;IS3MW>1>?c;:844^1`Vp]dTRA0Eqj@V
JG_ae]`Q6ceE4CSM^P7JOAhDjpZfoJYh3qVP2;b6Zb@T1k@_Bk1;CCqaC:c8^4CV
:[4=?MHoR?cG<pmB3^OE_Td=QD_@XMm_D@K11EJkLqfRhaM2NpF;OCjN8PAO^]8c
N^c_cgAn58cedgq7o;@E5?=TL27J2kQ0n]c3__gQRZ\KUhARB>VSQY4=?lEq`bXJ
1\2qjBRIoC7TS1glZ@gPk^m_pIG19iaS4@PoVfW?mP2OcN2HS39TpF>PhX?Q9BSj
c\ghfJ3_6X4Tj39QqZhNT1K`qBBRKW7R5mRoJED2KGJLIG2]<C1>mG8C^hC2i1mp
I<3jQR[qSCl2Nl?>\ONR8N0]hZTp7m9H<?fq=bIA=6E]aZmThgdLFLVVm2oEB1p3
Nd\k4Cpii6D11:DCQ1PkN^S^hEl6iZ\OgJ5<giUVU]DC?HK2i]en`QSFl\O8iMEm
;p@1K4l4T5h6FAm:gTmDV^qZ>g:<?1A6ikBkK^^ILmlE:JTYEJq^ceW@]CqochFG
7B2XnMGeMPUl;3gCBk4J0ZGpb2FD1kfpIfR7oW2`HTaX[TUi5IHeDLF>ko;GiS5M
MdZTb2ZNHQdaNQX>bA<GQnUaF`2mqfokN5ZB55OiUoiBQ>Y<1q\oKHaSc8U;[RSH
oc44`bJ_C3WO>pm^g<0mTqI76B7@YNjaJm:@gR>A\]ik;6GN[ApW\9;=:aqiBfQV
WXJc:9V9=7lD9KGpcD?HfFc5c;n:B6lSCGfYIj]N86GpO<S>bhP2;fKMSCAMUK9M
CAXVF5\JC=Xlf:dM[o[]<Bq49iCD:`[^hPmiYn3BX;b0fe;\@Pq:>0LD3?pM\77D
0cpCXdKkX2LQX?>8>fc<6p7m[oHemNXj0nkX2PQ9apgd`9hHipd18^b7qCddh6X\
@4nTW_Vk0dknFR_J^P2n:W6qg65:LF6qG3d7jTGoW2pFBf9?OMpM6_;><J8=?G=E
Ik90ibW>jXU:A6;Le9N9i9a5WclFIq6\IbF0Y_m<7^TQSWUULF4g:L]e\qn?2Zkd
3qoHMS5K4pLnXBc\8q4c9?6mFq\l6AmdMSJal18[0b]<UXa>Idc@g@O]CoA9TpG1
P6P`@VgVc0JL5e3b4]q]h5lO6=;D5[gCAZ6<LXn0NY5MMN1DSq2=VhBSP:l@Q<17
JnA5YLqOPVZfQGno8dP40hZdFCRpVPT_??hp91Ke^Ve:hobl2M:DJCmIPQc>pPa@
bOGgN41WcS]LaC9=qT69]L=^^1=iN9P]i]e`I@A\8?niS=4\U_J4p5\aF^bdACX2
Y4;<GUKb_mRZ51cCq@HFcJImpT53@\FDB8TU3J33c5OfRTZe5pS19:0\SigVN_:o
acW_MpZnN<mGTO<dicl3dPgE[I?DM8i\@dmjQ:C1Nd0N\7q2B:U;j_]V@VIoNB4i
ON<c_5bcEEV`36S<g9qV\e2C;[pTAdkGJ_$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_down_keep_IO
// Cell Type : Primitive
// Version   : 1.5
// Revised on: 5/12 '03
///////////////////////////////////////////////

module  pullup_down_keep_IO (io, i, e, pu, pd);

   input i, e, pu, pd;
   inout io;
   wire io1_tmp;

`protected
A>_7MSQH5DT^<>WXam34^0[Z@d2k<W6kiMEbNl3kLZWgO9eYbm7QZjo4GB\YKopY
D0kQOT@Po`NB5XJem1k7AaGBkN\Q<<`5I4pS8C3b_2dcEYE\IAMZQS4kkCp=>Im0
cp:gOcG9mlZ^CN^`?bgN3AVB?@6S5p>k`1aijJefAa_43p=N1>YU2he?3<VJSjDn
UOg?hd_?molLVSpTA\=G\FHKNXA_L0M1\?]B\aW4fg]q6V[S[4^^RKdF5e>2\Ve@
Z4N1::`Zqk;Lb6[Jf>3NGk0dM:on^obMkdjTQn]>IV9MYp5`lPKJJZOmW5:Z9oL>
AefI`bkA3i70UgWV^Eg@oSAepTO7akIfJE_mloGQqbZOY:01K1LG5i`7\cTD>H>_
k`cQZ_kRTPi:LG<feSJ<=qLj0<ZSb8\3VBWS=XWnVZE?UI?8]n8?2[48KELo7YS0
2:58p2Dfc5m5H:TWSi1J7NYe7P63I\cdZfoZbkW[oh5gS^S`NcLJ[i^XAXeqX;fj
@j1jjk@06=?cTUV`75[M>VdHdTB24[]Mc>E4G_X^elBOcPe3:f:nHTpD2AA;Of0l
ED`nLKi2efW^Oj3BSg>V77QoBfa0c;RLOlqMhH<S=qLTJBCC19G6aYhA]VW<_ImG
3Q=58>q9]0PB3?aIfnS;en0j@Y;_ZiKnWp1MbjeSV;1oM?BQcb6d@iNa<2[1@jJX
M;VbQ?XPkq;G2V864L0]Ie4=@28S5^B7Yq:V<742?Dnc<Gf@MTo78[JMER]nIQIc
f2ZFLqhOXb6@=ph<WiZMaK=2EJE:OnTFRc6eSqFm6ZUjAC>Z<DFWK=Onl0h=XqZm
\ij^8pH[]UP37MMEYhUgMI4R6?l@1RIHP7NXaiq8G]BZ;7<QofSel2F1O]=9nS\G
c=[d9O6<W6W^2qfI?5ieHqcG>d5K0O[\PA]IipnL7Y[>4oo7:Ra=K2piK0@ZoRmN
`R;S34H;hL3V60qVhbf5XBi6FOBZK[QbgnB<8b9gMfh_H`a^GEbj33pAELN;<TNX
_ND`QnTW`Eg_BpTEEElckA4nfWN5[d\CHBTXp^M7jkNI2]aTnkKdEf29q`P7Bi6m
hCCb<iDn9oMQ;ZCqA@GGg?UemW6bmUWO7\`_FWcmF4qGi1=^YH40_Se0[TbI^Qi@
W\MJO;W6Cpk_XO0CfY]oj?b@nmfER_fN_BfCPQ>J^9f=pclkLm?1n@YD;KX4=YgJ
=9:0h@KdC72;h`7q1aNkGnHj2eIa0kCOaZCLmTbRT7UA4\jq75FS2eW]M4IhFF=\
na470H;B@ZKRRXJ]70Wd1o:@pXf7E5n7WUebEehlN[K]J_9VAYXV^d2>i7H7J4l6
q4l^IVQMZh9O8hbVPS6E?73hHN1VOf`3Fp9g[d@n6bN7BjFX_f?fRk_mhCM[3Z0J
WN3SW6[3RgDGM;ihpfRcmV0eI:a6lI65o]f9WG?ZQ8YHY2kJ@dL2\:VN6DOf1U3V
qJebM@g?9>jnIiRE`XNn2g3WaBUl5F70;eg>B?<k[^<Q6YP6Wq7_<fLLXKGKJn@l
W=4TTQQnZPSDT0R9[q2U1l6Hm<fHNNSSUe6IEl15abg=YI>iS5S]K@gaJ2H[?Id<
DqK@MZj]5qcQKOCNgW=gE2j7XR=U41=J75PVCHd>fp6?g=;41T20g`ao6G8D_h59
L5jm_;Zn7HqTHiDDVIGg]QS`U;6;dX3dj4=]R9U@Y_aR6Mn3XWg]DBh3fiaSFem1
9eqaMCWk`WqTKn<c59AbjbKPlgUa0B<39N`9:SKHT2^UXpW4I?QG:Le\meA6S35b
eqXBVKOHCql9jNH=I<C>[MlPQ\nm_bGl6d<TPhq[=>SIU;63djBhn`Ho\??NVhR6
i>p>\?5NX_qmk=oNdYp:Dk5m@SY;7Qg94fFF67AMl\AL[\dEa7kc>DJ0in6oOKD2
S8D\BUX9AE0dl^<ddVbIBCm0bDJq5GflmHc:K;j53`g=hOYi<^:G;28E^U1p3bZZ
R;QI>o\D;>]?L\9nTWNfiZjpH77[gmZq<RJibA2pm87XDe1FHfl=@`X_fEOZ`GSm
c[mqGQ>GX6<qMQOgL5<qJMj>O;WpUoc\T4P@f?i?42H>VN:pgnd:QJh`oX[`JMMg
lS5XIlZU6<k_0QcV:aO7jIoR5;CDU]?^n??MpO_3SH_MpLk0VcVYN;17N>\Z>>Fj
5n83[Tie4qPl1@aA?ncZ6VicgCKjLm=mJDG5mq7YEJTF2p;=dB<>Dq5a72BohA?d
E;]55Z0e5md3hNP=71^PSqc\Rf19WR`C_dk;6\6ejfF^OKQd6AcPDU??Sae_55mO
8pO7DgHR\SX2l[DjL_EoCY?3mJ>81pmZo1GjZpd^6:d86qiJnPYa7gF^_]^POm:Z
610o_:Y_1qRMBV4GLqm<9YHU2pFDo9Rg1pFMSTLi;Fe4HSU7hCXNTp1MWW?6SpJ`
joe_1fi^WBgDJUQccpHoHD?WP\cSE[`g6m1ibWHAYMJ=Xq1HX45`DplPkQmYO3n8
XDnY2\ScJp6BGK_KmpCJU<^XmEDHT2:8`hbo9cg:R`ZU;d`>qe43<Y6kp4`hOebD
cEmp5nW2Ka^pcEWZ848oLo>a_61o9jn[o^bDX>ipUak4J8CjfHZQh9NMd[GD`F?`
@\[V0Nc9p[49X]FKpUo9<ZKHqncnfIIGqE1`4Pc@pTnMY?nfO7jASMPYQpZJU_0@
Q:N1BYPMEbHI9[oEhdm`ZDci=AFK6I@5kZ[o8VeUSUPSe2YJc1_W4FK]39oDfgom
jqd@_5=;XqLGkhK[0Co[XCG:5k?6P=[kXdZWe3=9p^nEJYD2pg<]kDPE6jnKOgb6
7R:Sq@4kJfP<inGVgmO<E\PL5ZZ;2T:_4jUi@6KqJT5XEoU>cF?Nkm;R0ZcpKWo9
[nAp0UeYF7o:UZ6o\\LAAWLK9KN7MJqK6RT:mXq27A9fL=kSVl\nCejl[XMqej>R
c::]gcIil^M[gOn0hVkXoc:qA`ADC`1q8flV>WM;[9DWaS2eB3[Dl;T@fHSI4Z2O
fa^q3I9EY32]b0=6F=nZfGZ1N0E?OC91pAl11h_Mq21O>42hNo[Pc1eiBZBJQq9h
>2J`l]gAR;ChLMlNb:LL=8eemq57QY`kCKB>0<oclDQ6S[VRP\PQ89jdQkb5c^p\
_[5b7>qF`SLNBKaHYJ1SH2e]_O?XM@6oAKAp<]HX1MCqdHjGj5RMbkh3YbD@V\Wo
qJRS1ZKZ9;l:PDedR?M27a`^EoePp?J96Q4Uc?UB^Y5YH8H7J@T<9<`[p4FfdZd<
YK;QNbC8m:iW3OlM_K3\JOba?12h7A6>5dG]?J\YCpdnEcOL>pKk8aI?Dp=7A<N2
5k3]5^HAi:94LpG7XQ4`DpF\2E4OjYWF=;F[2P@m@VpBRP13dZfR7RkCg8:4nGFm
W4P^0pCAB:F7Vp;6=^PlHeZcb_nD\nE=lWphbQm>\naEXKV^EIcbCVm18m`[hdp^
f5N;Hnp6`LZ8QIEX0ITDT;gl0^Kn@C1_cAZq^QJPHeg9n=9P1C>aEMJ6bXc2W6WK
G_^HPSZ2jTQXOhnpC8eoSNcq>Qjo3[3?R;\FL5g8QH3jp]F:a63Zo`3G7NZ\73[O
Oh\Nh]ZbqmL`8<hM_4^0gYN<cM=GW0NJMkPG:pAH@M1EnqHgD5A?<<DL9\3QjHS3
`aNji?XV9RpBA:AfnBp?FL?gV7_]6@B8MoJ406=qmF8NZT36dA93OIJMCCeW^lB<
S>3qZ9aCC=Pf@WH@Old>H[T=AXcZ8[0pEFG9NLhDgd2WA>?Ak5h;_C9n]mSNa=Y2
]@eDAX\:2ORF]L2o@?qfmHTQYGqA`PXLVGq:VWXTh4Y:MGm<C0E0l_pfjVi=h:q<
=9lV]iL8STJH7Tm9_F^6fe^Qe:q^6YJCl`pgloY8311SBMcDj]:Fb7qf67BXNW1^
Yc[[XpCm_CXXCq8>_kP5Ra4l?JaH]b[9O3]RWI2GoP3iq68CT[iCq\m1llnREA6p
BYdhe_Mq6@S;eQfEa<VkhJ=2T4hTJZea`B4pdVIcUncqm^L=OXT5dddgob_Vp1OS
l[YBqKRW5LkCpcaTgl6]qUk4SN^8KKYa6_A5DEh;fbDJ_KKKaOZfM`;lpWVl6iO7
2>KALZm:WPS<@CN0oN355Cbq`9=fmaT30VGOPQI>^ZHU^;JAieN^?N4qOS>A1L\5
m_>]W0K[P8[Apno4c8FM75?hkY>=7o_UopPSWUEGUiZNji?\5T:mX1>?6qoW^iF@
8qWGj_IVDbR4gVZe[qEbbI3UVALQN4gPDVnlL]MZLVpfhGWH7g6FGakC@;8>LVp;
6aE2VE0IPJ7mo_KKgRfUAIY7`;W70dPX0Spk6ei7SJqD_P;M9fh\N[a]1;KdFN`f
:Znp`mJmMPH^8F^Z5jPAQd<pM3E8L^@c55D:6ndOk=@glXC?meh1@I6`W_<pb?7L
nmI>RnIk^NBXlCZ;[hf[T;1ekK3iY`DmCbMoYjG^bo9XJ1Z4H3E[L\ClgUV7_b@q
UiGOE6npMl\o>a4PF6o6D6bHMgJ1Uh5=KbipSS>RN^<S58bcom5S\n[IHlq>I>7H
L1e0aN1O>]5iC0_7epehX[``T4CHOlaI;<=R>HgW5<d6DKeWPTSV=JMTIibRMLm6
LXMmqOK3oKNlpl@fh`6Z$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_down_keep_IO
// Cell Type : Primitive
// Version   : 1.5
// Revised on: 5/12 '03
///////////////////////////////////////////////

module  pullup_down_keep_IO_03us (io, i, e, pu, pd);

   input i, e, pu, pd;
   inout io;
   wire io1_tmp;

`protected
:1Y8VSQH5DT^<<IM]:dG?;MC\_;DGhg4fij6LE^L7B^PkbNBM@I5UAD9WRU`P?lP
?3h3iD0E_4DLpnlcC[`LUOhI61o;qL`5<=6Vk@N6jJK0dl@]f4bS9Wi4h;0DMe>K
_UMaAhjHN1IVcEYTXhCELGNC8SPMbj^q=ab\Zmp^aOSTW^ZWgL6KLJn8ChG^fQUY
^?qB:JHCUfo3c_kXZTp:eAdMLc@h15bM;D0BN9NUeR`mg5``SNSq47lRT]0Q>7HM
n6AMeK6E71SM>OK8qohFiTFi8R>Clf?WU=;PZ2f;kU9^jqOEOh4c;XG_NMH_`0T`
kQB<[i9QhFTeiAV9p6jP_EVGlSjR<Gbib2eXDgBFg`cjWgCDC9Qg\p[Mi>bGYFPJ
8@<Fn\iW\J11D>f<6fcXFB>`OOb7HTVmp1^JD>7n34`MA6k28g\RA4<SiWg__CU]
jIN?kn\:9VemfqLb77=;0\G<>jaP^flh1<Bd1aa2JCinZ\59o:g?Z3H9=\:XgKdn
6TDO>]0_@dKNpnYIULi`\@f9@@gNMR1leomPWWjOQYj?AfTk=oW9iR@80Amq3Go>
WjFWIDWU7nM0RRC0GHk=aFM^P6SncZg3Q`^HN\2R@XicjGIV4cpfMb2>Ng^@l>DO
3e<OH^`\GX`1oQ:oV@LJcJN4hda9WXqGh9?dhqJ6GFYQ32[2c]HUb[9]?2ULOTbL
7mqaI]6i663H[eN@TbBSn0jPKHclopEBDXF\PHXeA>PmaYh3[_OGo;@8_IZ3iSq1
[;X1hMY0I=4m7C8Dj9\GliM[3nM7_JbTiK>UI1qT:ChQR965=oMLK\@N8_ZToJDi
CdN3VNd4E^qjZ_RY]Lqb@HH;<79B2N>Y\]9IGWLJhgp1\5l5hWmWJ_?E4Scj3N=K
TVpZOTlDn1_T415MX<T_gm:O^S6X`[pfR<Ed6G4l@3K<Q:_HBoMY@TQ4[C6lXp59
m9QL`q5cPU<jVE[N1fg64;K=[XQY\G\@eUOL]iqSc1RCd84QhYO3ZSl[a8dko[W>
VA\`M6_[07qacJ`UDmc8SDL?ZR?7C7U7`?1PENdicQQ>24f<klf;D:laalXkdcJQ
JM00[2p40D5Q4Cpmg3MS<e07\?T8abq^5cO8Sn03NBAYYocpoZaXC9kKW8foEVnY
4IJd3l8p;agMM_WJj6G>DkU^kX6G5_O7]SB[cWO>YQ8mmRaqfTd:]?9>_?J<oX]i
1@eHA_p>naGL:QO9l[Z[OJBMoEeCkp82BXE?\dmbCjg6hb^U7q75_FSn58hV>PhN
d[bocMX64>1kp@4=9@HoCUSK1Kf2Ha`JBXdqZ<8hKT8M@WnNaMO^QL\E3Oh3Fi6O
OPpglB;eeP29j[I@la85I?_C?YW9G7TJnG<Heq@:8;moFdbIUeN8C_eRfk92VU7a
XS:bNLF=pXJ:6e7Z`?TNbDkdPWj`9bHDTX2XaYI]p=mH9nkZH7Ba120@=PURjMZ3
NH6k[Q[a`[Ni;@93CpMoG_i61mENg<dEb05YSSdN>UpV?P;`DOQM1fXll[boP<6k
7bH2=mX_S^YqC9<5@8D^h<ioiH[<72W^P:5UafLMW5=NN?[Ek\3_]ic:H8pL:FJZ
3RQO2DfjA?ImhZ9PS6Vl=E_b6LGS>BYJbY73:N;0LjpNIDZGJ:WKKR^cl\Y?=<J2
ao<WC1\hiO41Gjf8?HA]gO>h`j\q65ImTMHh8E<G7RYF<VcEeSKje=U15jlg4`Pm
ln\4KZMmA:>p]C4XnCXqfS2BS<m@eI:W^Ab@OWDJ2`XR1T]hdTBp=GW1`H4FlAjh
E4=:N5`15`2Om6@AbfcMqfifbW^@qVe=mJY?Ce@A5[V<GnEXh1:oNkbL4b7b>aS4
gHYb:PBbSp[:ZP9D5e>N3GcaU2159<ThmJ8?SAR8QIbgq2FaXP5f_@07O6a?BCcn
qLIJZU\_qXKTYW0kBPjgmXfJ^ga5JnNJ5^L`cp`im56lF_KUeDS`SGR4<BY^RoWG
m=9ki_0WiF\5E]Za6U\OWQ7NDWRg9S7@1qc6h[U;iNH3gUoR>nGRH700b<m=Kqf_
fR;V=qF`?]icXpa_NE8LQ8DoPHE>5IUCWKL_@NG<GH]P>pa:UGYgheGRljKlGm?m
V2MYJFEZlp`l`;0n:qP`dR35Nqb`ATWWg2j1lf0??l<f:Dd21b0X`p_MBEH97848
WB<`o5`j6Ba0J:1^L4k2EDMOdXD4@CM[ZlSE5<qI;>[dUEq=kM09gHqcX7>]B9q]
0cbQBDE\dY;\XTQ_U7pd=XR42Wq^Y8LAE8^cW@An<CD;eHNJRBWCX\dqQfBm>[6B
]J?>K8G\:`[ljGhOF0bQp3CP_KHJJ7jZQ5I4W4<oi<hA2kJjpBDgYg66q4IhLKk3
p7keeAi6^Kc>IQ<MJ?h;9k;Ae\3ROGH;qb8XH2FcHj558C2Gg45^2E\fm08AqnTl
k?ZW`bAh3iS<Ua9M8FG`Bn`Ni<SL?3@V<mW3jpk38^`^<pF4aViWMqFfeoLY\CfQ
2a:1P7]4cg[0GF7ZQqT?K_Ym1qMNOOngmqbC<:EcLpGQNI1NV]Eml90BCo`c2pAe
]<?7QSiogR_BjFU[WnF:[M5J?Qc1HEbRa:moq;9:AYE<qA@?4hjd_K2e:iI7_ZaH
_dQmkigBqXV2c\F\paNlgcGO<[lkSVL?^84<pf`[^@EZqMSRCSTD[Ah\Gfek6I9g
9n<A_bJHo^<p`iEXZ>63]H5Ygn?mYA9MCYMOINR35d:n@hoWh?mEG6qYmm54j=pN
nFG5ah<f^qZBJifdYq\@Ra2G<UXRTMle6V@;584b]78X:qS?a27RT8iOLG>cKl8\
LQJZ8?kT[q=I]Kch8qTl8h_bgqNBfG8i@pWMcD3neqMGFOn3\:\^Dj?^i1Z`\\PT
\Of07<Snapc?2D^FVe0S>^G>4HqJNG49<1pia4aFDV5mI20<869BhcaN=]LP2Q\4
2q_VS:m[Up5=][FO;gQkk7@:XUiG^>dOCfXI9F_RO1\Cq_89fNLDf;]QZb2`a0D:
qYcBJJ\Qp9o=o?2YYoc9c9[D5B5hbFN8X?6pDXkDXB1pEVm_W66lQm8H]4SNSiTF
;?HX4?C:1I75aB<]iT_:]P`?:E[`WJV4hRTB8VmiQ^5q19TfjhbXD_HQB<``Z8Y;
pag<<kWk<\dNm4@GFCAFFB;ME=_4p1PNFn[=p1`R<6:M\4Mf]f@>kQ;OWYn@1djQ
JplKZc_KQpUlI5RE_LFc7=`K46TNGlpXCaSQQ5807e9<3H4TKN32\hIEc6qJo;0m
nI=eZ1>b3H9:87OfFD_;RA37f<hTbH@<j1qhc?MnCUqW1Wg<SCLF2;^1EH@MRMU`
OK6Ze`Jp_iFHG8fp34:=bObT;:OKWoo3`fI3q`iX:^n=IhcKX4CYfY;O^80Amd4f
qj\PkK<BLhClSTVG0i=B1Uj\6=dMpllla9IdSIY3Hoc:@N2lNBmoE^hiA<W3XC9o
Hp2X:Kj?3pmIj7RXap:Q<AOYYQh5e?iMDZ1hZqLo=HU:0qPUHH9aTM`fIIW0cRU:
45>P``GQqZ?anjZTq4S9lOUCJNQJn:`GD8_jfCAIgTO8AI<gomEoT[_>`oB9jqM5
:58D>AWik0kIEE`Y4;qZFAjkU]]FZ=4dO7Y0=B9QJTZdd;p0AW7Q5hpCGe?HO;R0
RDjCkDI3lH_3ISM<5?ApPR5JoPhqTfPG7KmhM:>IUQ9NSC7:2c]<d=U=4`fGAX]Z
bnF`5OD56bg4cllq:RLmf`b?Aak10l6]0kKBqE4Ln7W5J<BMMgO?G3eQgSRKXeiH
pAJdI;L7pH6lh^DC`\EcOT3T`Hgn6bg46_EnNpgUWnW_IpSD=4;?WkZdXAOH5Ueh
dUp@PMK=ELK\<I[Fb33:T?Ji_W63F8ql:n7?4N?A9LNNjE:@7W_[5\:2kRqWY:fN
U3qM5g]87nSJ80DOkI1ZCJXQjcM5VadO59HTh:K<a48gWOS3i5fnh?@W\^OYa2W_
c@hpS430YB0qLUR\B;XXgdPAge]4bU0p1E5]<:nq6=A@K2TTaSYN5Wg^jgGbclQ?
9Ldq>5JO4m8pln0iD2b]ZamjR[YU=2YpMl@k>_dqPQ4^m]W=_:UZK>BlH3i2FV13
4DP0if?L^9pF:Fk9RPgWU9ZkCefIdE8DchUjg6\`Wpb7<h=YYpSL\1_V3S:bq:J@
D>JPpZFXOd`EHGN><SGdYVHL=V>VXnZ7pbgn^:9lpEl8EV^3pki_57g>piI0d]B4
q5AmliLWi9I5bFKnQ]Hb:e?gmLLB?kOGgCkq:8bh0ID7LS]@C]8>ShN9<17<=c=7
\mY0m_jq4g<`0=[15oYA_7ALNeBEo8>1HYl2Q6qD=`=Tb4MRd^?fil^;P48p^oeH
hgA>D^HQ3D:fl]<=qCm^gKB4VMNI@bNVhN_08:acq:=>a6Uiq0AA`oLPFTP9KSeC
\^;5X@1=LVDS]p9fkoShjKnh65lRMJ>0K@cg1ApnaTRH\6oc;E=FMbKi4<qGViW`
c>oom2m=<KSaNGAiX7CY?[]`<=n5\DqmBlQ1ARqXQd8Xo]emQ7A]@>Aa[2Z:d_cq
ZRa[nUjhHHS=DN9=\2epJ?WU2`dOQLg7_l<:[2gEa_lBDThAl1bP@WGgD6@p]o7l
l]<qal?m0ID=6\SeFUma?Q5H9DDdaZIq@gnGP14WYJSF]GM\NGT;JIMFnl[4QhWX
8IU4iP:NfFj[\AW0L0dm4n?Kb[OLiHnJS_hVDgnQqLeYVobnZ1bOa@e:VNQCR^Cp
kRne:H`Ofk0lNW>@H9Dk?6qMIg6HBSq8Bn4@Dl$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_down_keep_IO_IE
// Cell Type : Primitive
// Version   : 1.2
// Revised on: 5/12 '03
///////////////////////////////////////////////

module  pullup_down_keep_IO_IE (io, i, e, ie, pu, pd);

   input i, e, ie, pu, pd;
   inout io;

`protected
jOMCkSQd5DT^<=XMe`1?17dIB5j1[=p0E9P_X9@D_TKXE5;J6IK=H1`3TM1@<ET5
ISiPZgh1AXLfkYSoh7C_6=[q\BC_RB3^0L_hDG]TKMZY[Sj`Cg];OAo@9Mq>ELbB
1qd6b8c4nX4HL@599EeKXNCJoSC0:qF3dMm?6p9?EB2KVC@_hXG^BPI?oD81=Iql
1gUZc:gH83E_EUIMWJ<kOoqdHY;SmYPp=S\MfILmdnGk3ffbFQ519>iR^JWnBlU\
pL7:D7fenp`oHIY><B6IYA=Wiq9o5n<j@NIQG[?ZAb5F:KCoYA2gaG?H9B<\8bNA
;qLX@Rf^1?d3m8Y_SDqb8_NF40gfe\XATbW699Z40=pb_hijH[ChDA52]B;2CR<1
IZF;In=oM^Z`ScGG\IpWY46R\dicGc?algg^BZC30aGJPT:WJ3S6JQGVLoB5i:Ma
;PLED^JTjX7pn?7B\ZKa5]>=MLg_WhbmQ8p0I`8jA[Wa<NF428JDMAWYCpVeP?k2
b1X6TRa7Un3Dbpe>FW?>A7h^?aHWUhC_FM_6p6E<Bc<a@`@4Qi_fAg:K^HDKYd\l
\>nqV_[:;=jJ^k9^bkiC@Y_kfbR4[Y_;DdGh8Gp`iUo<6ScI:OFR^`9i8YU5oW0h
Y7Z:FKGIjqD17@>L9H_C<iENZ=0]V8^AjnSSD2m?3\dO_Jg:`VX14537e=O9MOU4
^_4jLNNMDgpl_^65ahkG?2RkEn4fQibW@@ZiRM:BThqYCINZbFIo?3:iAkVjTEQ3
hcEYe]U`DO>PDp@Ff?mBoLG<_5BHf]YE_n>hmfOh1hNJIo^eVfC04]q7beP3lbZ=
blbTWDPESN:N\?^I0naQo47q[GD[Kh_J7>ITkNLh=<L080Ya;INURZhFn07P3Q^2
RbPch1q`aJi1Z45=O6l0<_[Sn=cOg:AM1Z?eg@X_eKAb0No6hUgYI;qMl7Rj_]6L
\bNXJ;\d2_jSDKI@RXKRNc7mX<Y21Pj?Q20MN:mpk13DLm7\iBU5;aO\FD[W4aJ\
\Yh=mWbf^K@c]A`ckd0[o85dV7n;hN6=[VoOp\U8mXPfk\B`7XoOcnWg6[LEpb?f
8hX]pi`oFjL^EihM2l`Am<ScAH2\GdaLM9@QpAJZ^RG90EU;ek;;QC8;X`a`IGkX
4SBb8pO<14aZlq`BlL2]Em@S<GIAXIM`\S4<3Qn]X:?60eM<omPEiUJRkOqcSHN<
kWHjMhkDE`>H`DNp?`dh^c?3E9I8=m9bJk=;qYBGoX]oaj^37RTi88hPTqWfJ`BD
2fRM=eRQJ\;O[G0KJ^5Z=Hp:QW;O_`h549NO5>^UVDfq>@T72ZmphJ`jm7E_OklT
jeB^G2AC<:7:<KOJp^fK7QcoVbWBb4WRSZ<>?\_gnI1kp;@6O1m8pI?`oYgSq9P3
<dT>G;4NF<D]GhnXCl`Mej\T?3PSq8OF?Y4HU<1NWBe1J_h0nmdZ49\iAI4>c>Xd
NNYn:_H=g>j7h0iIP0HZ\E06^CI@f?mjq3SF8QEJGim1N1J6hGD_M:EI3QWcp>[m
[Z25qJ@YnYcfpO\:XgdAEcB_aeol:]^iMOcjOM0Dqki2HHk5q6jY9f\GqN2RO;<>
\O6YeAEc^T[[c1Im:Nckm6nQYI8Xq^5dH@FDqmhnJ5o7]E8HIAX5CheGVpj2JNfI
IOg[6F;HM>K=@1qR>^Ell?TV2o^HAjB\4_cqmJ60iMXaNAZU97n8OUOYq1i=F<Ia
BY2AfO`K6jf`4qC:AJV4\0@ULkSG3=hVC=dG1p=o[kd]fp7\2>>43Z[Y<ObRKL2M
0n>Nbd>KoOqh[Z85JjN=84;>k[BVjBESa0T\;TqSDkbIYMpgaI?c6:pO1I[_`SX@
UmHE2l]CU;g5j6?I>G\HA]hdMFFcm`[bI82ZJZ`@Cg<3Som_HQZDjRGh:p<LSn=9
flbjliUg3LB2`4YNMlfLn_PikpjeBcFBY5:3VUGO3Nmjl85Fo\:MEpIZk>FgPp0K
o298>p1`Bfg50[NUBfV2EG]TlF5c@_YoDqM@50KY2qkfe7oWaTIId<XOjopKU5KK
[]q<;eD7A2q:HWTTh4Yoeb5Q@`?e>aBp[;^>G`H1<danm7?1fd5kpd>Z:m^gi^Oh
Jcj;aJf1<p]fQX>bbc==U375OH_:MWpPKPBo:T5R3S<In;A^]TRHbf=>cVjWnVlZ
[iCKV5`[eLj5IcOS=2UPXmo<X@MiFd;cipJ>Sb5c9pRBaeGQQFTmTeP[7e3T7Mj_
?0lDdph1Wbo:6q3L?jS8Sd\eJmB_SJJP1kplglXZD4qC><S`;a;_PEED:G_0<k14
UMe\;A[biqlB3Un4kqC4=0dNf7RB_@XP1=Dnp0Tj\Fd=PI9qIHTZJ\0p402Rnc@]
c^oXjG7[dZKngmLLecYphi`NQh\pAb\UUndqJmci@_kKBGC_[CC7WbqWXgPcj3q[
RQVf96qLg\9;KhWFa63<4IVpjeD7UZOpT:A51VK@8RT3HARn8=jUSOHHDK`0eaqa
WV^h1K2m9E@KI3AiWFdBmcmKQngoX;66>NZ\FeeZbMPcOdU5E<^F9>Oq]oAfinep
<Q\\f=4?RLXXH^<S^dna<kDnSfU8W4nRdiXgJ:e9O`RCpOE>mS`nW:T[>DWUOZRS
Lq=Oc78cHBO2GbR:U@WL:4pj?glgK;;a\a3ibV0j=6Lp^RCN67`L`N7bjR``LWOX
p;aWJLU7pf]f2SkR<ViM?c4=j7S;iRJCnF`aT9Zoca0naa@Lm1R:8k7E;e:@:2>h
cgM2?JnQqXc?Nf6lFQjoo27cX6GPC7=efYJp6bm3Zj9q46A^@aASbKR1JdoKSNPH
pR3D2<VMMGR6OlY^M:NT`]>C]HI2pA@]0OL;qCOi_=]nn;3DiK[o1<DGYEXNbago
9pB0o9]Lcq5bBjofAQ=j>HO;LflBjIj[V0aea4b5qJD0F5j=1WZ0QcFleUHTcpNo
eSnB;FgW>F7iD=_f5=gl=aW^aqS110oPfp;d0KC<PDWmMFoCUROcFjX1KUnMDgpT
^77Qh`p>NPEY:^Q\WfTSoT\JQC6qFFfY0OZbYU]I1MO:bfEGGm3NWBaqb0Zf;oU:
O^48GW1bNj>Kh2V@>G@C2AP?Uh14HPo`C<lOTNID^0SOnfbY>]X23E14pFgg[`1Y
4Udb9>XZ^BLVbZTIFOPcp]U5VfiBqaR7RQ\MpK7eE[:MHD]YOcVXGW:00p:EL:1N
[k]6hc4D4M=6OMq8FEJjBQ6>LZ@eLF]^f;NfA>8foU`G_W><Kf[N0Qql\L:\eZjT
^UYCSMbdG0cqn:El3S87iP4faB6ggGbUqY;1\_=mE4FQ:o;ehX3@`p^]fGY6hp@I
8f543c5@NheP@Z`]KAP8c3LGAE2W;Sn[NlH<[YID7XpZ6aB\[L1GdhSVI5CnW??E
IQB;5pf]EKmZXqX:U@gh=n=eZg2WW@<c::p64?^jQ?_LIZ=3cJAFeaObIgR6=5pn
W1ZoEfpWPf`SljcEmaYg3f5kbM5C4b3C`>lpA2\cl`0qEom5X`Qfef^]?MP>@5VX
jZa^O`o[qTbbF?=\^TR?F`YK=GZd_qhi?;m5IVPT?Mda<N>G5CL`Zhi8ApE?KXWN
kqk1S475QMoMlXmc?O77>13FYg01@OpN7R[GnAqNen2O36nnkEW\:@hK?EDp>dcO
Rjof>;BPKD_QnBR:a4YnMc0pbNj;4G]Jk`OjRe5ZShaLc=6J61DVMc7qi0oXR<jb
SoPT\\a4e2=Kl1W^bejpD9kTY:_qjSkZe2CpEbmHB3=TB9UGBW@??cjn2oUkfa34
Ukp^L2JT7TSe84;YXii?[P=qdj^3Q7FG6n?Y^cPXj12@qJ=2e67VNG8Ge6l]@L3k
MpcJ@A5bl6iJAGLV8iCi=\p]HTRXWlqMiMUf^jU>UoTok6\6c6?M;8V1j6pQ8mDM
MVqlR2AL2g7hd7kG[MHNSLaG`lFh[mfB1:A3R_G;KflN?7^JbD1W07?Q0IHaWpUJ
V0B?5OU8R89aan6kTTqJLmJK=9q4Ycfml<@H2TQHD?>>gOPJ\o?Ibc[NWpoF6[9]
aqEijlQTd1A;HoWN;AbjfOR38peS;Q`7<DJ1pOL@CZ;=qmC\^XP>8Jgl1hiE9aQK
D_2:o_D0pTYH^6Uhqi39nJXEpcM59>Lapm>;D<ahpAXoMFE`41@dZUOA=m`PPLec
;f8lkm_KiV71;0Voj7ISP5MpoD3k[35k5NNefb1kmUZeEfB916h_B\SRh63p?>F=
kSjIVdOn6<7MQo=kG`8[Nn7c>Pp_3UM_hL6A@E6RP[>?JMopoS@;804AHG5dVb3N
HINbqI\9^B>>j6gE4hKl_0OlG<LKpnEmW?[?q:OJ<2n6cma5c9=E<><l3BfWLY@W
jo:gdL3Vd5kF[4nUV9<:8FDW^TFklJ8;7CHSp;KR3WdbOhk@GbPXLhT@EJRZaq>2
PXVPflJ3LA<9PZI4Aq_ZD[UW;bj[BencWfi:I:M^genQQ28BijIe<pcH0oVl4p0G
9P=1<aE9]@ASm;I5FO@]Cip4UR4KG<SEV<k7C\706Tq>Y8aCLI=_VYOEhTS5_ER5
;LVLiJ]U1^XD6KpK@SBf20q=ERQYP_jkbdkO>Pm`jPNB:URi7?8Ni:cnk`B[c7EF
DRf=?NAf:M2Oc6gJ\iqb1;A>@NeRG9<I@64G_Bd04\7L?]pFELnCWKA[Y[?AO0<G
c6Ojnqen9U<o@P1J2TWfgX2VhFV`pi<e`XLEl3eeldcU0ZTf75@B<nBbjMlgq4d5
m9EBpOe==gam$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_down_keep_IO_IE
// Cell Type : Primitive
// Version   : 1.2
// Revised on: 5/12 '03
///////////////////////////////////////////////

module  pullup_down_keep_IO_IG (io, i, e, ig, pu, pd);

   input i, e, ig, pu, pd;
   inout io;

`protected
@2`EHSQ:5DT^<:Vh]L`ddgdUR@0^T;;l^QJlIdP5O[JqG1\5JG[8EVf:a;C6SDT@
JI=bEGU4pHZSi_CaCJP?j_Eg_@cE_XeR?q?R8VZ=qai1o6MH0Mk?K`fDG76LX=@R
J=@1p\U^MFi;ph^<8^_^40j`cBU^U^gEJLRHXqK3kka:VN\5Ii@BSYf[BoCE8q<a
@;W`Aci5AYK`iE<C47U[lpJn<gh;22pBBK:LkYn@JYH@`noMgQD;cPO4OES92hnp
63gWOKkFp9IoT1QYA@`@F`LVp1Di?S[2AMUZnHPS_qn1RibN`kHBgeg@nDDKmXcb
3pH7N:8i=kg^AmZUbApO@lbUPn?WT8]2]\jJ3TY6F:PCRaHa7=?AiO1h>ZqVl^>[
^6jgfCoXGaHR7olL_peBRWaCN5<K]QF5]GXMC:FPqLKkPj6`5;LCTM4WWJZ7qbA[
KiRh2E2aL>PCQS`oh\Cq^jL[Ff>7N9leR4:\]1;=<l8:m5<l=hp]15N:?mc[Q5:8
BXM[RUE@9TBAPnKcVpaDREf>bbLHDjYF\KU^?6dHfm[PUJ_nZZ;]p^lXN<]:]QWj
U59e:U^=Pn[gR:MT`fJ>ElnpJjee1G^Wmk22]?RdfhllfQRFCM2O?9Jqh?UcRC^[
UFVQ3JG0KJSg6fFkI__N7j4_EVpCmmGQ9DFkMfYh\3:FnG1UN82d2CZR3_Zj?LdK
JeKqBK4A[Bl[XYGRm;m3ZB47Rf2hT[8KEFc:qL9Dg<Ffc=R;Mo_fU;kd<hM>2f=P
WCJ2R@7hWJMdNY0A4]]pe2@AOIi;cXhNSU:mZHE9b7gT40Le<ZAP5;;3e6gYY911
EMHqCm:?R<70<POZQ\9YiS17ck0iE3OPeEVqV3NYK9PJ;bTY]4>d5APlfU342Uhe
gJFACFmIKdOY<5UBYReSq?aE\IeGXO>NH;GDS?e=ecAK=`5W0jnUUB[iag;ZYQI1
Z=9f@Eg<Dn<_N20X3qkmXJP_`pUkf_6b2d]`bd7Q_5E?`:\GJ;B5JZJKkqWGi6Vb
G`ALm`j]XZ5:BQ8C:4\:X7i`P1q5^gOV2>ZA7JI<Ck;pJhUHMZGpBVm@1m_C_Tbd
=ZZS6;hl:0WMNLfN0h=oReRM<OT?5M^<q6ndAUf?_T22ni?Tj1NKJp8[nmRNZCaX
B;dWaiC@H<p:a@k:K0jRUHNc?HF]P@l3G4;F8]YE]m<Akl@<2@lV;YhOK[;hTDU^
^0Qgk:p<Dk>G5JA?=b4B:hCEWCYqf2BIT=SFeE=CJ;W9LYQkqPiel6THqQ;9Ai6;
B9g:V=o3?WH_pN6BfMi?6kFLI1d27gKMZ[l[j=8VcpAVddhW4ZfZOL=9Z9hEkPPZ
W@[UlpSgimADCp:PdoFH`pdd54QVMWng55hPf@G_1n:hWA802Z_6?pLJ?9ek3>oJ
0]IDRg^LC<U6RV7=]pm:?3La8e^[59=<kNUhKq5^Pi@U9pgack:k;qKe^6UiPUH6
M<jRQHNI;J^QlXgcXqVc;`0h^pn?KD`\MqJVkBanZqP8d3H`d:1MGSL_[1@JmOq=
4Dk2_\_ef1ULhlIq7o?8Fl1_i=Do1jGeLObcqj43;jE@RB0VY[if4n^:BpnammC`
Tf;6>232OmW@`dpUmm[aBR3PlcT<N\V;nggq5lG\D?UqVb?TaCadoeXb]6C\BcXW
M=<Ca]MQpn5LRAb^@bHFKa:oac8j\UagG3=JpDb4\XQ8qo6PL4CeqTWk>jn;_0DG
@Q_S8]5KmIQSXS\GALnKc7oE6R\LDZQ_K>hjqdaHMZ9SHFnf8@<:HVRXdTXDQR`U
CG=jq5[QEgFM0[Tg:3KWclk1_YkjVFd7pbLIE@^TqC>G^H^[i=6R7QJJXFQlEeWW
6XPN]=2d`;S;XVSTqnOe[T=7qL1?i3ECmX`M]lff[il]bFLmNS_Tq[B_EmLOpcSn
EWeCq8ZnG`j4p7]`[]HSYVgdSSDRMcV[OQ0aDh0IEjU8OR2j>797Z]R`NphRgmPb
8[[VCeVdLK8ib]qkfRlW^b9MA@X1;h>kY<ipBb@0Y@1`ZD4H]eB8^Kdoq?T`Q70T
>SZj76LWMce3JpL2Z>4^KpF1dnb8F1:Qg\iI8g93@RM9KcVkGqM9bEe22p:ZE=;9
jGG1U\3cO07WNdX>6TGHX_QVZ]IR7iQXKPlXB_I>8G59DoC1V=<X5^>nCp[aRV?N
C@kaTY?oE0V_V3qDmdA1?9q?oM6Ae3^]21[B?W]]`S=FO]RgkZ4Y[qhN5Hjbbq>h
0f9HiRTop<Uc8UC9pZO\kGeVCWal0XOo4V\GBPGniFL;pC?Z7`a2p=nfiYdII4JD
VQafaaG^4:;l>STFQn[eeA0IP1QiA^:lf\R@X=5UFG63hN\X6h?]<iT9bRecqE=K
W]ekpe6LjWjmpgkWa[i>qeU5H\keo`_fThMcZq`]YUg5YqQ0Y^Ie:\iT^1`[0]hD
g8?2>;R<F]6Yq[FAEF40qoDnS:]>\>EcDZY[SS?[3FPUj]dd[ZgRiddaR@eZ8e?a
np57k9jInFh86cGDEolIJ>qU:dnJmZCQ^fBHPk6FQ@K]gZgmj3m05c<JCepLDB;X
d;@eblFi56WdEW0qdhOahoWMUld3PUeC3G5oqW4[YbjQWkCAaTkj_m379p?J]f96
=p0S`Wo]F<a:]ITfJJ1:<=6GO6K?p`F:=b?WpS==7KFf=Y;dc@19nHH:XP?_e4\7
0@8H;QImZgR5niBVlQ0ilg`09cmCb1`onij23MQ^:L1q[4NZWESEZ3`O3DEEV10`
pSi5NMa9B>L4J_2A26@X^cd0`niTpUUJ<m^7q5b^0dA;BPiECEIAkL_Ll?\TA3RG
RqlCWe8J0q_A3SF`0_;JFde_`PI?OQp;9LP;]LgEa3MTFni2^WWIPohS0<qRQg`C
lj4DZ_X;\E[R\Jfm[0FUCZ:nE`P`8EJqKgPkof<qR4;JOZj`6LWj>HTfVK:1?O16
cO94q[;GNIV5pi;ZSeJXP3C0Rdd=ebX`8pbZIV_GP8cg1fD]No:Me^6?6;3i^qC`
[=iglKTJj;YhnS8oEWLZ@U`DM]a6??]KeF_CA70XNe12A>kY0q;TYo_Y7n@FTeNY
a@C[5S]oZI8b`qcRl^Ua<qWPNn<>bpZLVm7S?b4PTUTaBnI4OaqnbkCNW73;JE@:
ZZC3LGLpiWR1>878<oP_`7CclE:Rqe56IRdKXia9@>[42_S3mqhDo@@@0L4ML6Nm
Rh8?CgpVPoU>8fGfJXCcUNN4Q]=>DmI:RRN@5D@cX[dOG942NYn`PJe>LHm6K8`W
WfHO>G=_^ReqYhAUkdBpiKMMYCD:Ef1f=C\;Q=MjJ@f`cYp1BlA0b_p=mSZSVPLf
PEFNEX42N1OqbBnBHQ>@B3da2RilAD>6jmF@;6hq;hXd6F6qkc22][O5WlUOgbPQ
6;R1i^Z?gBD]p6?UAo:8qd^D3VZZ?^B3D9bYlG=Wi<kmB2ATmLD\BkjFic^J1k[H
fja=Y`b0MPD>>WKKONe@]dgpJ?\D9CA502OPeTEWg]>ipggWjE7OalC1B<_?9fh;
7coCbX@fqh4Uo5DeqmH6>9a9a`[MMS]B:`X_;R8?jFF3Yp3c?BK;@q:8KREH^kbf
CWYg4]QJ^]pNSj]Y4@[ThfJSYReeoSoI4G@E^Xq^>i<4oc<FSnQ0QjLngS01V81=
94q4YCb6j_p@^[EZLLAX_JUbT7Yb?36Um2JAMg8nmJT]<M0>K^E5bTYb?gkhf]:e
\iPOoaflb0AP6b>D7qiK7F@ggphna[SDaEe=^`67k^PEDnqbbkKNi1f^YdUji[9k
[6hpakVYdJT<:NBOhVl3B^OVpVCjl4MJE<mh>GAN]L41jqFB\`Jhl?j>[A_SMVcg
GFgQ^R<oH\>Kl;kFMb7e1aIbbh>@S3o_aIC3Yg9Ya0>7SlZKCP54Nq?L>RR92p@C
kVkn>27fkVahE^Ji26XgKIJaYqA4IAQhXqOk7_3i>C8E6a\4m`DIC:qNjGWgC:pa
NUg]OJ@kJ@BS=>RKGV\\^Aa<[XgfNqUb@o>Q6h^bC?`Sa5c64DL=<6dcM68hq2V1
Hmm4qEM0k0Yek^mq8@GLO`Tqh>a?[4cZ@[RC;=5hl1@>:c0cjGSpKhMPgJ3p^SJ4
OAmpUf_RZD2pkgg48H`1SfO@k><I9\Q3TS3[7S:Jk3MP=0q4U[bRb@q48YdmRF[>
IEP6eD@dP>?YD[;6CZAOhlbE0hp@cSIJM2S=T5=75kGTVB`=7De\2O4K>p6<m@mb
ERR=5ES=@eiBbip\faAZ^ZO[=ZkE`QDn>X8pd[^>U?HZP\j>LliBh7fcHF2qm`PE
0K`pjg[9[E3mGS1Z^M:ndd[5@HN@pe8G4?Rla]kU?1H8OB4nq@RlTUB6>nnCaBAg
FYVB4?YbZ`H;Cj:\Z6h^ERN5_`54oC1:^8m4c0jFSJDbijC3p]]KZ2aVjG[EJ9b=
ed7NG]eUdHi0dm_a:TIfq6;_Y3`OphZWB[odE0LjdKMI0Q7Q1:@eeqP66UCGf1bb
ZR\Udk65Ep]84?8cJiUW<>02UC1fgS27`G7_O[b<LcZ2PqfV2bgb0qjh@_O<T\Vl
:MAJBMDbh==MKmbA0qkI4=T_RfSjd]82IC`]Y\CkqcRLn\Z[?Cfo3gY4\9V:aA:q
ckAeWLIgkmHW@01:@nV`cIp=feJ4LUq=UfH[6Q$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : pullup_inv_IO
// Cell Type : Primitive
// Version   : 1.3
// Revised on: 8/20 '02
///////////////////////////////////////////////
module  pullup_inv_IO (io, i, e);

  input i, e;
  inout io;

`protected
H9lg4SQV5DT^<U`:7g9e:im[3><jjKmoF`L=>go_798e=6XFWe<f4LiIq2TD9;4E
[Bo?PSYcdk^h7UHo\FhaLQYcW_h1XB5Q=oe[NG9@Y8<ET9J9L[SmKpnCZY;2N@5>
@oX;RTaEb_mf3;7ne@h2Bg`cUF2jo<\WT>D@Wh<4PZ7eh4P89S>X=pUOK4DHqlIV
i8C<d@]M?79_4gZMDgWR3^f2p5S3b:ki?Y7kYNSqdEne=cjU=4HFW6=Z]DnD0dqc
=7k4Sd;;kPjB0lc@5;^0lil3fnpFCOBDV;p\b2AB=Bme5WJne:_dFn88H<[qG8NX
;nATFT?1[j5\8OXN]BZqRN]7SJO\pJ8HPO[:]VkN81=kEN?k6>]9\ofKG>_pUoCQ
aP?SqO5gCXOhJ`FVj0@=pkbo4jfFeI0nWXZCi0lWinKOEpYMR91eoFN2C2MQ_0>9
oI46C_XFZ:LTYMUZcO[93MgAa]D``Q866f[Xeq;gB1X0mk;AQLQ;H_5]8_5gl5?L
1N:mF<:cpFkZ^\<AG<Ecl547UK@W56bp0lQEBZCQNe?M;Q9FV51IC1q[nd`8@Yg3
F@0kELoXH`0P]L@g?fEAC8q;@M[ZR;P[IE8ZA3g>k4Oo7POIY?<5Hm76Fm;G38>q
Rng]1h]5bjgZOPSe6gMfc[22NY5=:[j2qCV?iMB8GF8hP^L^`SCaL>ZO3k5k8>OJ
0BMBMWWn4T^O9R@pg3PGP<i64Yk^N?_UMVM7]0c]nYgMD>l0mQCaj7=9hIj8VFNp
0WGH`Je]D]h^o`RGVMO0Rf[INK7_4ig6i6m<g>QXMigmTPZ[h^I^Veapd6mB7VUc
]HlC^^9HHB63?DK<QQPB^=HaBXDQ4jGq4kYR@:UC`P:f]l>B00^cq=nn`TN^q0[2
VWdPTe2U4d`_El>J00\VNYdX8G\=bq2KSdAaFpR8HbYnI78:T:<LJf7^bmP^pPSZ
>`:3pdaf\05RS0QZA8C0KL;gNb<C3eogk?iAkZK[pl`]mJ6PpFQCF0B4;RH6LE_O
NY`iaI_@NK6Sb3g>ADh4Oqb[?7D_d4CEE>;EATc7SgXklDg_L_pgkac@QnmEbGkE
@o2?8KF>W[G]6:qBh?k=?;qJ3]lVU]pLmC[c1D_M92<ZD`6>=T;0ZWLH7=pfGe_O
iSpkY7`1Y:OLJXIH]GSZ6]Cd>LMS6Mo;fHf^79F2BA5@BIUiKa0[`6JH\9NQLapB
a>1:nTqJ;Gf=ZlqoMU_BhJXe\[g@FoFqZXd\_APBND9`AJ6QcYVNi1G>HMclWKQ@
_``MIfMkFYPB=NFdlC6jJj\SKZBB2UW<MF@>qhkYWC9mp2K5oTMHR9fl9<A;PdYd
5N7@U`Sk@Y[qmDm0=:bqlHmi16Wad;3aXMdi[^ON89^DeXpYMlLT:aqYE0>HJ@E^
=G?Wkl^NU>:A\p84H7ddD11:U7oQ?H[Khlj<oWbc6jXX>j@QPEmXT^4FLP?;fO;I
^X_TMZVVMA_`pJ][H^NJGAP=7BbN6TZjbhJiEkeLq2;H03l5qkK]Z@YDIF<J4n;=
J7f<c\]3GV`ghpofd_8[MVnLYjlgnIk7B7UQFBK`fiC>C2V^pAl11h_gqGL@kA_@
@PLF13j1K>^IR=AqmaOTd4D_@AH]YY5B?CRaEge0XP=qTYd09HmpPQhC0cZIDbDl
XBEDIk_g1kFAD[?Tq4PM[RiLf9Ljfa=<_ZVT83cHG9=hI7U?1iDU`=h4`[N;qHc;
24AhpGE0dHS@X6`GXo:hPc;Il`Lp1l[ZoZRk8oQT9W4;Ci51JS\j4iTpjg><LeMn
<GfOoASMcSVY:o?kTScqZFn<PZTp]UG6Y9bh=ROJ^?giWO^R25>PcXA`FkfG0[Kp
K`ZU_:lqOANT]=HpEQCcc;KAooObCH_dW[PD7OFaqh?Q6VGF>^QaG\MBe8bJcUM>
UMOjjABQb`\Zip@@JNc?4PL;LdS]9dL56gp?51DU[ahW6;3C;5Tm1_g:0n5f5n0c
HOeiEAqRRJZGg`q56Y9n?4$
`endprotected
endmodule
///////////////////////////////////////////////
// Cell Name : tffrb_udp
// Cell Type : Primitive
// Version   : 1.3
// Date      : 11/02 2001
// Reason    :
//      1.3  : Modify protection method 
//      1.2  : Deal with unknown ck.
//      1.1  : Initial
///////////////////////////////////////////////

primitive   tffrb_udp (q, ck, rb, flag);
//
// TOGGLE FLIP FLOP WITH CLEAR/STANDARD DRIVE
   output q;
   reg q;
   input ck, rb, flag;// Clock.


`protected
Xn\23SQH5DT^<dmHa0>Nc[J2lYQo@RG6?MU@TiP@IY@LjJRIhjbmc85mRIfa[f6[
WfNEJ3Tp=mPPbSbN_SIM\0i48M9c8Y[EXC]Z7QC74VmGSB8Af?j]3WUg_6C<OBcV
70^m7bM:IXq=Nd4U2lJH1VH7\2D\9Y7`6l:KU3SdGkWn<V7hecU32Ga24Mk`Bq@Z
YYGXpB^f0DU9qWV2Rl2o@Kfg9ghoHf]Kf5^fgpmO__j?B:f=8CX`ARnk>WcGlHpB
9;4OT;mh2NFI=]I6WjEF<4:q3PLH3\TDO:DPG;Apc0_D0e8]c5L`9aoBY;Pg`P3^
C?78piU7k66qNZRJN5gh_JgLbEglQ@1Te35>MX6NpaLmA73oEflKY=P<W:hS7Eml
jpoA5ZV=Xk7an;B2NkRi8<i7eYq43JW?mT_c_VRYa^imBCmiG`:C`E`RZG<9d=A_
iP]>9JV2TYQWdqd8S4F\T$
`endprotected
endprimitive

///////////////////////////////////////////////
// Cell Name : tffrsb_udp
// Cell Type : Primitive
// Version   : 1.3
// Date      : 11/02 2001
// Reason    :
//      1.3  : Modify protection method
//      1.2  : Deal with unknown ck.
//      1.1  : Initial
///////////////////////////////////////////////

primitive   tffrsb_udp(q, ck, rb, sb, flag);

// TOGGLE FLIP FLOP WITH SB & RB
   output q;
   reg q;
   input ck, sb, rb, flag;

`protected
ho;nYSQ:5DT^<<mRL^OdYTe9q\^603SF;I5]a?Wi^na9hTG?UneNV_kp8FS>Aa<B
OJQ<^3EL;[_a554lW?<aB7PipRobfeDqN]O@I`jp?KNdZEFdLSW4SJ9W[J52LMKL
I0Zp<ZkG@L7nK\K3Q1LcVTd66foNG`39JaGDh04;>g@[7>9VL6][9HJn5KS8;[=p
_W<i0b2^i^H5bFb;6fP`hejfj=<p64RcAU;6?agid6eZ4SOmFZU]39VpLl`:1b`@
^aYgAHP<ik:?P_G7]`WpUb27n@cQX`f2iFR]Yce\^nJUZNCA>ThpT<mI_^KKl;ce
omN\J@E15nD7MLap0gl;]5<<_[LR3JhBV31:S\1Ek7:pDZcYS`aS7Q_chROMLk[G
8?L;bP7p0Y\`GXae@OggO9<Bh?moUfE^D6cN\LYUe4Rp:T;6`JNW?djFG44_U[Ck
MBk>JOoqEh@P>Cq]XD93YDePe_HTWjke5W?cM8?2f_A`P@pIYVUjAi>[29Qc;j_=
NRZ2G1i:V>KYhFS43U8\QA=pD8hXG8TTiD18JkH?iO7;;Ge0G`\h_0DqFYOjNj9k
0ogUn=S]DP10ni3DQanpVOQ?H]B$
`endprotected
endprimitive
///////////////////////////////////////////////
// Cell Name : tffsb_udp
// Cell Type : Primitive
// Version   : 1.3
// Date      : 11/02 2001
// Reason    :
//      1.3  : Modify protection method
//      1.2  : Deal with unknown ck.
//      1.1  : Initial
///////////////////////////////////////////////

primitive   tffsb_udp(q, ck, sb, flag);
//
// TOGGLE FLIP FLOP WITH SB
   output q;
   reg q;
   input ck, sb, flag;// Clock.

`protected
DlM@RSQ:5DT^<m21DBg0aAT6a@X>@Vj[3FSAKPpU\kkEnGEbC1o[mbc[\H:CHj62
`IGBXaCR?Zp0Uk[ZTXOJ6j?R><XUSS5U2@AT;ikp^1ea\0qEmYJ2AXqnCc>>@?;1
Jd4_1Ij@YZ\0:_JplTX`\K?dFYEZ2M1?do;@PXGnqLo^86\LGjTebTRe\S7eRKS1
Mq88Ebl\CBc;DGXX\fI<L6MKhl3J0lbQUbgFU0MXS]_[E663fFWVhq_7NMC\6C@;
35he;@m5=l_PIIf?_]q:\DRD?p?cmMT3ZR39<bL0J?MXb]GYH]dMFNpe]f_7]mWj
77M49bMhI_?_Xg8qkoQiC23fD_?1_>dbddB[9MB5pMUKPESI$
`endprotected
endprimitive
