NAMESCASESENSITIVE ON ;
MACRO CORNERC
  CLASS PAD ;
  FOREIGN CORNERC 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 235.6 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  OBS
    LAYER metal1 ;
      RECT 0 0 235.6 234.76 ;
    LAYER metal2 ;
      RECT 0 0 235.6 234.76 ;
    LAYER metal3 ;
      RECT 0 0 235.6 234.76 ;
    LAYER metal4 ;
      RECT 0 0 235.6 234.76 ;
    LAYER metal5 ;
      RECT 0 0 80.01 80.01 ;
    LAYER metal6 ;
      RECT 0 0 80.01 80.01 ;
  END

END CORNERC

MACRO CORNERCD
  CLASS PAD ;
  FOREIGN CORNERCD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 235.6 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  OBS
    LAYER metal1 ;
      RECT 0 0 235.6 139.28 ;
    LAYER metal2 ;
      RECT 0 0 235.6 139.28 ;
    LAYER metal3 ;
      RECT 0 0 235.6 139.28 ;
    LAYER metal4 ;
      RECT 0 0 235.6 139.28 ;
    LAYER metal5 ;
      RECT 0 0 80.01 47.86 ;
    LAYER metal6 ;
      RECT 0 0 80.01 47.86 ;
  END

END CORNERCD

MACRO CORNERD
  CLASS PAD ;
  FOREIGN CORNERD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 140.12 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  OBS
    LAYER metal1 ;
      RECT 0 0 140.12 139.28 ;
    LAYER metal2 ;
      RECT 0 0 140.12 139.28 ;
    LAYER metal3 ;
      RECT 0 0 140.12 139.28 ;
    LAYER metal4 ;
      RECT 0 0 140.12 139.28 ;
    LAYER metal5 ;
      RECT 0 0 47.86 47.86 ;
    LAYER metal6 ;
      RECT 0 0 47.86 47.86 ;
  END

END CORNERD

MACRO EMPTY16C
  CLASS PAD SPACER ;
  FOREIGN EMPTY16C 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 9.92 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  OBS
    LAYER metal1 ;
      RECT 0 0 9.92 234.76 ;
    LAYER metal2 ;
      RECT 0 0 9.92 234.76 ;
    LAYER metal3 ;
      RECT 0 0 9.92 234.76 ;
    LAYER metal4 ;
      RECT 0 0 9.92 234.76 ;
    LAYER metal5 ;
      RECT 0 155.59 9.92 234.76 ;
    LAYER metal6 ;
      RECT 0 155.59 9.92 234.76 ;
  END

END EMPTY16C

MACRO EMPTY16D
  CLASS PAD SPACER ;
  FOREIGN EMPTY16D 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 9.92 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  OBS
    LAYER metal1 ;
      RECT 0 0 9.92 139.28 ;
    LAYER metal2 ;
      RECT 0 0 9.92 139.28 ;
    LAYER metal3 ;
      RECT 0 0 9.92 139.28 ;
    LAYER metal4 ;
      RECT 0 0 9.92 139.28 ;
    LAYER metal5 ;
      RECT 0 92.26 9.92 139.28 ;
    LAYER metal6 ;
      RECT 0 92.26 9.92 139.28 ;
  END

END EMPTY16D

MACRO EMPTY1C
  CLASS PAD SPACER ;
  FOREIGN EMPTY1C 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 0.62 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  OBS
    LAYER metal1 ;
      RECT 0 0 0.62 234.76 ;
    LAYER metal2 ;
      RECT 0 0 0.62 234.76 ;
    LAYER metal3 ;
      RECT 0 0 0.62 234.76 ;
    LAYER metal4 ;
      RECT 0 0 0.62 234.76 ;
    LAYER metal5 ;
      RECT 0 155.59 0.62 234.76 ;
    LAYER metal6 ;
      RECT 0 155.59 0.62 234.76 ;
  END

END EMPTY1C

MACRO EMPTY1D
  CLASS PAD SPACER ;
  FOREIGN EMPTY1D 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 0.62 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  OBS
    LAYER metal1 ;
      RECT 0 0 0.62 139.28 ;
    LAYER metal2 ;
      RECT 0 0 0.62 139.28 ;
    LAYER metal3 ;
      RECT 0 0 0.62 139.28 ;
    LAYER metal4 ;
      RECT 0 0 0.62 139.28 ;
    LAYER metal5 ;
      RECT 0 92.26 0.62 139.28 ;
    LAYER metal6 ;
      RECT 0 92.26 0.62 139.28 ;
  END

END EMPTY1D

MACRO EMPTY2C
  CLASS PAD SPACER ;
  FOREIGN EMPTY2C 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 1.24 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  OBS
    LAYER metal1 ;
      RECT 0 0 1.24 234.76 ;
    LAYER metal2 ;
      RECT 0 0 1.24 234.76 ;
    LAYER metal3 ;
      RECT 0 0 1.24 234.76 ;
    LAYER metal4 ;
      RECT 0 0 1.24 234.76 ;
    LAYER metal5 ;
      RECT 0 155.59 1.24 234.76 ;
    LAYER metal6 ;
      RECT 0 155.59 1.24 234.76 ;
  END

END EMPTY2C

MACRO EMPTY2D
  CLASS PAD SPACER ;
  FOREIGN EMPTY2D 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 1.24 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  OBS
    LAYER metal1 ;
      RECT 0 0 1.24 139.28 ;
    LAYER metal2 ;
      RECT 0 0 1.24 139.28 ;
    LAYER metal3 ;
      RECT 0 0 1.24 139.28 ;
    LAYER metal4 ;
      RECT 0 0 1.24 139.28 ;
    LAYER metal5 ;
      RECT 0 92.26 1.24 139.28 ;
    LAYER metal6 ;
      RECT 0 92.26 1.24 139.28 ;
  END

END EMPTY2D

MACRO EMPTY4C
  CLASS PAD SPACER ;
  FOREIGN EMPTY4C 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 2.48 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  OBS
    LAYER metal1 ;
      RECT 0 0 2.48 234.76 ;
    LAYER metal2 ;
      RECT 0 0 2.48 234.76 ;
    LAYER metal3 ;
      RECT 0 0 2.48 234.76 ;
    LAYER metal4 ;
      RECT 0 0 2.48 234.76 ;
    LAYER metal5 ;
      RECT 0 155.59 2.48 234.76 ;
    LAYER metal6 ;
      RECT 0 155.59 2.48 234.76 ;
  END

END EMPTY4C

MACRO EMPTY4D
  CLASS PAD SPACER ;
  FOREIGN EMPTY4D 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 2.48 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  OBS
    LAYER metal1 ;
      RECT 0 0 2.48 139.28 ;
    LAYER metal2 ;
      RECT 0 0 2.48 139.28 ;
    LAYER metal3 ;
      RECT 0 0 2.48 139.28 ;
    LAYER metal4 ;
      RECT 0 0 2.48 139.28 ;
    LAYER metal5 ;
      RECT 0 92.26 2.48 139.28 ;
    LAYER metal6 ;
      RECT 0 92.26 2.48 139.28 ;
  END

END EMPTY4D

MACRO EMPTY8C
  CLASS PAD SPACER ;
  FOREIGN EMPTY8C 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 4.96 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  OBS
    LAYER metal1 ;
      RECT 0 0 4.96 234.76 ;
    LAYER metal2 ;
      RECT 0 0 4.96 234.76 ;
    LAYER metal3 ;
      RECT 0 0 4.96 234.76 ;
    LAYER metal4 ;
      RECT 0 0 4.96 234.76 ;
    LAYER metal5 ;
      RECT 0 155.59 4.96 234.76 ;
    LAYER metal6 ;
      RECT 0 155.59 4.96 234.76 ;
  END

END EMPTY8C

MACRO EMPTY8D
  CLASS PAD SPACER ;
  FOREIGN EMPTY8D 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 4.96 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  OBS
    LAYER metal1 ;
      RECT 0 0 4.96 139.28 ;
    LAYER metal2 ;
      RECT 0 0 4.96 139.28 ;
    LAYER metal3 ;
      RECT 0 0 4.96 139.28 ;
    LAYER metal4 ;
      RECT 0 0 4.96 139.28 ;
    LAYER metal5 ;
      RECT 0 92.26 4.96 139.28 ;
    LAYER metal6 ;
      RECT 0 92.26 4.96 139.28 ;
  END

END EMPTY8D

MACRO EMPTYGRC
  CLASS PAD SPACER ;
  FOREIGN EMPTYGRC 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 3.72 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  OBS
    LAYER metal1 ;
      RECT 0 0 3.72 234.76 ;
    LAYER metal2 ;
      RECT 0 0 3.72 234.76 ;
    LAYER metal3 ;
      RECT 0 0 3.72 234.76 ;
    LAYER metal4 ;
      RECT 0 0 3.72 234.76 ;
    LAYER metal5 ;
      RECT 0 155.59 3.72 234.76 ;
    LAYER metal6 ;
      RECT 0 155.59 3.72 234.76 ;
  END

END EMPTYGRC

MACRO EMPTYGRD
  CLASS PAD SPACER ;
  FOREIGN EMPTYGRD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 3.72 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  OBS
    LAYER metal1 ;
      RECT 0 0 3.72 139.28 ;
    LAYER metal2 ;
      RECT 0 0 3.72 139.28 ;
    LAYER metal3 ;
      RECT 0 0 3.72 139.28 ;
    LAYER metal4 ;
      RECT 0 0 3.72 139.28 ;
    LAYER metal5 ;
      RECT 0 92.26 3.72 139.28 ;
    LAYER metal6 ;
      RECT 0 92.26 3.72 139.28 ;
  END

END EMPTYGRD

MACRO GNDIOC
  CLASS PAD ;
  FOREIGN GNDIOC 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 34.1 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  PIN GNDO
    DIRECTION INOUT ;
    USE ground ;
    PORT
    LAYER metal1 SPACING 0.28 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    END
  END GNDO

  OBS
    LAYER metal1 ;
      POLYGON  0 235.6
               34.1 235.6         34.1 0         32.47 0         32.47 4.58
               1.63 4.58         1.63 0         0 0         0 235.6 ;
    LAYER via ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 ;
      POLYGON  0 235.6
               34.1 235.6         34.1 0         32.51 0         32.51 4.62
               1.59 4.62         1.59 0         0 0         0 235.6 ;
    LAYER via2 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 ;
      POLYGON  0 235.6
               34.1 235.6         34.1 0         32.51 0         32.51 4.62
               1.59 4.62         1.59 0         0 0         0 235.6 ;
    LAYER via3 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 ;
      POLYGON  0 235.6
               34.1 235.6         34.1 0         32.51 0         32.51 4.62
               1.59 4.62         1.59 0         0 0         0 235.6 ;
    LAYER metal5 ;
      RECT 0 155.59 34.1 235.6 ;
    LAYER metal6 ;
      RECT 0 155.59 34.1 235.6 ;
  END

END GNDIOC

MACRO GNDIOD
  CLASS PAD ;
  FOREIGN GNDIOD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 62.62 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  PIN GNDO
    DIRECTION INOUT ;
    USE ground ;
    PORT
    LAYER metal1 SPACING 0.28 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    END
  END GNDO

  OBS
    LAYER metal1 ;
      POLYGON  0 140.12
               62.62 140.12         62.62 0         60.05 0         60.05 3.28
               2.57 3.28         2.57 0         0 0         0 140.12 ;
    LAYER via ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 ;
      POLYGON  0 140.12
               62.62 140.12         62.62 0         60.09 0         60.09 3.32
               2.53 3.32         2.53 0         0 0         0 140.12 ;
    LAYER via2 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 ;
      POLYGON  0 140.12
               62.62 140.12         62.62 0         60.09 0         60.09 3.32
               2.53 3.32         2.53 0         0 0         0 140.12 ;
    LAYER via3 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 ;
      POLYGON  0 140.12
               62.62 140.12         62.62 0         60.09 0         60.09 3.32
               2.53 3.32         2.53 0         0 0         0 140.12 ;
    LAYER metal5 ;
      RECT 0 92.26 62.62 140.12 ;
    LAYER metal6 ;
      RECT 0 92.26 62.62 140.12 ;
  END

END GNDIOD

MACRO GNDKC
  CLASS PAD ;
  FOREIGN GNDKC 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 34.1 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  PIN GND
    DIRECTION INOUT ;
    USE ground ;
    PORT
    CLASS CORE ;
    LAYER metal1 SPACING 0.28 ;
      RECT 18.05 231.09 32.09 234.98 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 18.05 231.09 32.09 234.98 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 18.05 231.09 32.09 234.98 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 18.05 231.09 32.09 234.98 ;
    LAYER metal5 SPACING 0.32 ;
      RECT 18.05 231.09 32.09 234.98 ;
    LAYER metal6 SPACING 0.6 ;
      RECT 18.05 231.09 32.09 234.98 ;
    LAYER metal1 SPACING 0.28 ;
      RECT 2.01 231.09 16.05 234.98 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 2.01 231.09 16.05 234.98 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 2.01 231.09 16.05 234.98 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 2.01 231.09 16.05 234.98 ;
    LAYER metal5 SPACING 0.32 ;
      RECT 2.01 231.09 16.05 234.98 ;
    LAYER metal6 SPACING 0.6 ;
      RECT 2.01 231.09 16.05 234.98 ;
    LAYER metal1 SPACING 0.28 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    END
  END GND

  OBS
    LAYER metal1 ;
      POLYGON  0 0
               0 234.98         1.73 234.98         1.73 230.81         16.33 230.81
               16.33 234.98         17.77 234.98         17.77 230.81         32.37 230.81
               32.37 234.98         34.1 234.98         34.1 0         32.47 0
               32.47 4.58         1.63 4.58         1.63 0         0 0 ;
    LAYER via ;
      RECT 18.05 231.09 32.09 234.98 ;
      RECT 2.01 231.09 16.05 234.98 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 ;
      POLYGON  0 0
               0 234.98         1.69 234.98         1.69 230.77         16.37 230.77
               16.37 234.98         17.73 234.98         17.73 230.77         32.41 230.77
               32.41 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via2 ;
      RECT 18.05 231.09 32.09 234.98 ;
      RECT 2.01 231.09 16.05 234.98 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 ;
      POLYGON  0 0
               0 234.98         1.69 234.98         1.69 230.77         16.37 230.77
               16.37 234.98         17.73 234.98         17.73 230.77         32.41 230.77
               32.41 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via3 ;
      RECT 18.05 231.09 32.09 234.98 ;
      RECT 2.01 231.09 16.05 234.98 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 ;
      POLYGON  0 0
               0 234.98         1.69 234.98         1.69 230.77         16.37 230.77
               16.37 234.98         17.73 234.98         17.73 230.77         32.41 230.77
               32.41 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via4 ;
      RECT 18.05 231.09 32.09 234.98 ;
      RECT 2.01 231.09 16.05 234.98 ;
    LAYER metal5 ;
      POLYGON  0 155.59
               0 234.98         1.69 234.98         1.69 230.77         16.37 230.77
               16.37 234.98         17.73 234.98         17.73 230.77         32.41 230.77
               32.41 234.98         34.1 234.98         34.1 155.59         0 155.59 ;
    LAYER via5 ;
      RECT 18.05 231.09 32.09 234.98 ;
      RECT 2.01 231.09 16.05 234.98 ;
    LAYER metal6 ;
      POLYGON  0 155.59
               0 234.98         1.41 234.98         1.41 230.49         16.65 230.49
               16.65 234.98         17.45 234.98         17.45 230.49         32.69 230.49
               32.69 234.98         34.1 234.98         34.1 155.59         0 155.59 ;
  END

END GNDKC

MACRO GNDKD
  CLASS PAD ;
  FOREIGN GNDKD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 62.62 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  PIN GND
    DIRECTION INOUT ;
    USE ground ;
    PORT
    CLASS CORE ;
    LAYER metal1 SPACING 0.28 ;
      RECT 2.41 135.36 20.31 139.5 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 2.41 135.36 20.31 139.5 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 2.41 135.36 20.31 139.5 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 2.41 135.36 20.31 139.5 ;
    LAYER metal5 SPACING 0.32 ;
      RECT 2.41 135.36 20.31 139.5 ;
    LAYER metal6 SPACING 0.6 ;
      RECT 2.41 135.36 20.31 139.5 ;
    LAYER metal1 SPACING 0.28 ;
      RECT 22.31 135.36 40.31 139.5 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 22.31 135.36 40.31 139.5 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 22.31 135.36 40.31 139.5 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 22.31 135.36 40.31 139.5 ;
    LAYER metal5 SPACING 0.32 ;
      RECT 22.31 135.36 40.31 139.5 ;
    LAYER metal6 SPACING 0.6 ;
      RECT 22.31 135.36 40.31 139.5 ;
    LAYER metal1 SPACING 0.28 ;
      RECT 42.31 135.36 60.21 139.5 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 42.31 135.36 60.21 139.5 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 42.31 135.36 60.21 139.5 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 42.31 135.36 60.21 139.5 ;
    LAYER metal5 SPACING 0.32 ;
      RECT 42.31 135.36 60.21 139.5 ;
    LAYER metal6 SPACING 0.6 ;
      RECT 42.31 135.36 60.21 139.5 ;
    LAYER metal1 SPACING 0.28 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    END
  END GND

  OBS
    LAYER metal1 ;
      POLYGON  0 0
               0 139.5         2.13 139.5         2.13 135.08         20.59 135.08
               20.59 139.5         22.03 139.5         22.03 135.08         40.59 135.08
               40.59 139.5         42.03 139.5         42.03 135.08         60.49 135.08
               60.49 139.5         62.62 139.5         62.62 0         60.05 0
               60.05 3.28         2.57 3.28         2.57 0         0 0 ;
    LAYER via ;
      RECT 2.41 135.36 20.31 139.5 ;
      RECT 22.31 135.36 40.31 139.5 ;
      RECT 42.31 135.36 60.21 139.5 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 ;
      POLYGON  0 0
               0 139.5         2.09 139.5         2.09 135.04         20.63 135.04
               20.63 139.5         21.99 139.5         21.99 135.04         40.63 135.04
               40.63 139.5         41.99 139.5         41.99 135.04         60.53 135.04
               60.53 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via2 ;
      RECT 2.41 135.36 20.31 139.5 ;
      RECT 22.31 135.36 40.31 139.5 ;
      RECT 42.31 135.36 60.21 139.5 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 ;
      POLYGON  0 0
               0 139.5         2.09 139.5         2.09 135.04         20.63 135.04
               20.63 139.5         21.99 139.5         21.99 135.04         40.63 135.04
               40.63 139.5         41.99 139.5         41.99 135.04         60.53 135.04
               60.53 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via3 ;
      RECT 2.41 135.36 20.31 139.5 ;
      RECT 22.31 135.36 40.31 139.5 ;
      RECT 42.31 135.36 60.21 139.5 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 ;
      POLYGON  0 0
               0 139.5         2.09 139.5         2.09 135.04         20.63 135.04
               20.63 139.5         21.99 139.5         21.99 135.04         40.63 135.04
               40.63 139.5         41.99 139.5         41.99 135.04         60.53 135.04
               60.53 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via4 ;
      RECT 2.41 135.36 20.31 139.5 ;
      RECT 22.31 135.36 40.31 139.5 ;
      RECT 42.31 135.36 60.21 139.5 ;
    LAYER metal5 ;
      POLYGON  0 92.26
               0 139.5         2.09 139.5         2.09 135.04         20.63 135.04
               20.63 139.5         21.99 139.5         21.99 135.04         40.63 135.04
               40.63 139.5         41.99 139.5         41.99 135.04         60.53 135.04
               60.53 139.5         62.62 139.5         62.62 92.26         0 92.26 ;
    LAYER via5 ;
      RECT 2.41 135.36 20.31 139.5 ;
      RECT 22.31 135.36 40.31 139.5 ;
      RECT 42.31 135.36 60.21 139.5 ;
    LAYER metal6 ;
      POLYGON  0 92.26
               0 139.5         1.81 139.5         1.81 134.76         20.91 134.76
               20.91 139.5         21.71 139.5         21.71 134.76         40.91 134.76
               40.91 139.5         41.71 139.5         41.71 134.76         60.81 134.76
               60.81 139.5         62.62 139.5         62.62 92.26         0 92.26 ;
  END

END GNDKD

MACRO PADPOC6MC
  CLASS BLOCK ;
  FOREIGN PADPOC6MC 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 72 BY 56 ;
  SYMMETRY X Y R90 ;
  SITE core ;

  OBS
    LAYER metal1 ;
      RECT 0 0 72 56 ;
    LAYER metal2 ;
      RECT 0 0 72 56 ;
    LAYER metal3 ;
      RECT 0 0 72 56 ;
    LAYER metal4 ;
      RECT 0 0 72 56 ;
    LAYER metal5 ;
      RECT 0 0 72 56 ;
    LAYER metal6 ;
      RECT 0 0 72 56 ;
  END

END PADPOC6MC

MACRO PADPOC6MD
  CLASS BLOCK ;
  FOREIGN PADPOC6MD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 72 BY 47 ;
  SYMMETRY X Y R90 ;
  SITE core ;

  OBS
    LAYER metal1 ;
      RECT 0 0 72 47 ;
    LAYER metal2 ;
      RECT 0 0 72 47 ;
    LAYER metal3 ;
      RECT 0 0 72 47 ;
    LAYER metal4 ;
      RECT 0 0 72 47 ;
    LAYER metal5 ;
      RECT 0 0 72 47 ;
    LAYER metal6 ;
      RECT 0 0 72 47 ;
  END

END PADPOC6MD

MACRO VCC3IOC
  CLASS PAD ;
  FOREIGN VCC3IOC 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 34.1 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  PIN VCC3O
    DIRECTION INOUT ;
    USE power ;
    PORT
    LAYER metal1 SPACING 0.28 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    END
  END VCC3O

  OBS
    LAYER metal1 ;
      POLYGON  0 235.6
               34.1 235.6         34.1 0         32.47 0         32.47 4.58
               1.63 4.58         1.63 0         0 0         0 235.6 ;
    LAYER via ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 ;
      POLYGON  0 235.6
               34.1 235.6         34.1 0         32.51 0         32.51 4.62
               1.59 4.62         1.59 0         0 0         0 235.6 ;
    LAYER via2 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 ;
      POLYGON  0 235.6
               34.1 235.6         34.1 0         32.51 0         32.51 4.62
               1.59 4.62         1.59 0         0 0         0 235.6 ;
    LAYER via3 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 ;
      POLYGON  0 235.6
               34.1 235.6         34.1 0         32.51 0         32.51 4.62
               1.59 4.62         1.59 0         0 0         0 235.6 ;
    LAYER metal5 ;
      RECT 0 155.59 34.1 235.6 ;
    LAYER metal6 ;
      RECT 0 155.59 34.1 235.6 ;
  END

END VCC3IOC

MACRO VCC3IOD
  CLASS PAD ;
  FOREIGN VCC3IOD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 62.62 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  PIN VCC3O
    DIRECTION INOUT ;
    USE power ;
    PORT
    LAYER metal1 SPACING 0.28 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    END
  END VCC3O

  OBS
    LAYER metal1 ;
      POLYGON  0 140.12
               62.62 140.12         62.62 0         60.05 0         60.05 3.28
               2.57 3.28         2.57 0         0 0         0 140.12 ;
    LAYER via ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 ;
      POLYGON  0 140.12
               62.62 140.12         62.62 0         60.09 0         60.09 3.32
               2.53 3.32         2.53 0         0 0         0 140.12 ;
    LAYER via2 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 ;
      POLYGON  0 140.12
               62.62 140.12         62.62 0         60.09 0         60.09 3.32
               2.53 3.32         2.53 0         0 0         0 140.12 ;
    LAYER via3 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 ;
      POLYGON  0 140.12
               62.62 140.12         62.62 0         60.09 0         60.09 3.32
               2.53 3.32         2.53 0         0 0         0 140.12 ;
    LAYER metal5 ;
      RECT 0 92.26 62.62 140.12 ;
    LAYER metal6 ;
      RECT 0 92.26 62.62 140.12 ;
  END

END VCC3IOD

MACRO VCCKC
  CLASS PAD ;
  FOREIGN VCCKC 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 34.1 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  PIN VCC
    DIRECTION INOUT ;
    USE power ;
    PORT
    CLASS CORE ;
    LAYER metal1 SPACING 0.28 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal1 SPACING 0.28 ;
      RECT 1.91 231.09 16.05 234.98 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 1.91 231.09 16.05 234.98 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 1.91 231.09 16.05 234.98 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 1.91 231.09 16.05 234.98 ;
    LAYER metal5 SPACING 0.32 ;
      RECT 1.91 231.09 16.05 234.98 ;
    LAYER metal6 SPACING 0.6 ;
      RECT 1.91 231.09 16.05 234.98 ;
    LAYER metal1 SPACING 0.28 ;
      RECT 18.05 231.09 32.19 234.98 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 18.05 231.09 32.19 234.98 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 18.05 231.09 32.19 234.98 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 18.05 231.09 32.19 234.98 ;
    LAYER metal5 SPACING 0.32 ;
      RECT 18.05 231.09 32.19 234.98 ;
    LAYER metal6 SPACING 0.6 ;
      RECT 18.05 231.09 32.19 234.98 ;
    END
  END VCC

  OBS
    LAYER metal1 ;
      POLYGON  0 0
               0 234.98         1.63 234.98         1.63 230.81         16.33 230.81
               16.33 234.98         17.77 234.98         17.77 230.81         32.47 230.81
               32.47 234.98         34.1 234.98         34.1 0         32.47 0
               32.47 4.58         1.63 4.58         1.63 0         0 0 ;
    LAYER via ;
      RECT 1.91 0 32.19 4.3 ;
      RECT 1.91 231.09 16.05 234.98 ;
      RECT 18.05 231.09 32.19 234.98 ;
    LAYER metal2 ;
      POLYGON  0 0
               0 234.98         1.59 234.98         1.59 230.77         16.37 230.77
               16.37 234.98         17.73 234.98         17.73 230.77         32.51 230.77
               32.51 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via2 ;
      RECT 1.91 0 32.19 4.3 ;
      RECT 1.91 231.09 16.05 234.98 ;
      RECT 18.05 231.09 32.19 234.98 ;
    LAYER metal3 ;
      POLYGON  0 0
               0 234.98         1.59 234.98         1.59 230.77         16.37 230.77
               16.37 234.98         17.73 234.98         17.73 230.77         32.51 230.77
               32.51 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via3 ;
      RECT 1.91 0 32.19 4.3 ;
      RECT 1.91 231.09 16.05 234.98 ;
      RECT 18.05 231.09 32.19 234.98 ;
    LAYER metal4 ;
      POLYGON  0 0
               0 234.98         1.59 234.98         1.59 230.77         16.37 230.77
               16.37 234.98         17.73 234.98         17.73 230.77         32.51 230.77
               32.51 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via4 ;
      RECT 1.91 231.09 16.05 234.98 ;
      RECT 18.05 231.09 32.19 234.98 ;
    LAYER metal5 ;
      POLYGON  0 155.59
               0 234.98         1.59 234.98         1.59 230.77         16.37 230.77
               16.37 234.98         17.73 234.98         17.73 230.77         32.51 230.77
               32.51 234.98         34.1 234.98         34.1 155.59         0 155.59 ;
    LAYER via5 ;
      RECT 1.91 231.09 16.05 234.98 ;
      RECT 18.05 231.09 32.19 234.98 ;
    LAYER metal6 ;
      POLYGON  0 155.59
               0 234.98         1.31 234.98         1.31 230.49         16.65 230.49
               16.65 234.98         17.45 234.98         17.45 230.49         32.79 230.49
               32.79 234.98         34.1 234.98         34.1 155.59         0 155.59 ;
  END

END VCCKC

MACRO VCCKD
  CLASS PAD ;
  FOREIGN VCCKD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 62.62 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  PIN VCC
    DIRECTION INOUT ;
    USE power ;
    PORT
    CLASS CORE ;
    LAYER metal1 SPACING 0.28 ;
      RECT 42.13 135.36 59.77 139.5 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 42.13 135.36 59.77 139.5 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 42.13 135.36 59.77 139.5 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 42.13 135.36 59.77 139.5 ;
    LAYER metal5 SPACING 0.32 ;
      RECT 42.13 135.36 59.77 139.5 ;
    LAYER metal6 SPACING 0.6 ;
      RECT 42.13 135.36 59.77 139.5 ;
    LAYER metal1 SPACING 0.28 ;
      RECT 2.85 135.36 20.49 139.5 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 2.85 135.36 20.49 139.5 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 2.85 135.36 20.49 139.5 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 2.85 135.36 20.49 139.5 ;
    LAYER metal5 SPACING 0.32 ;
      RECT 2.85 135.36 20.49 139.5 ;
    LAYER metal6 SPACING 0.6 ;
      RECT 2.85 135.36 20.49 139.5 ;
    LAYER metal1 SPACING 0.28 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal1 SPACING 0.28 ;
      RECT 22.49 135.36 40.13 139.5 ;
    LAYER metal2 SPACING 0.32 ;
      RECT 22.49 135.36 40.13 139.5 ;
    LAYER metal3 SPACING 0.32 ;
      RECT 22.49 135.36 40.13 139.5 ;
    LAYER metal4 SPACING 0.32 ;
      RECT 22.49 135.36 40.13 139.5 ;
    LAYER metal5 SPACING 0.32 ;
      RECT 22.49 135.36 40.13 139.5 ;
    LAYER metal6 SPACING 0.6 ;
      RECT 22.49 135.36 40.13 139.5 ;
    END
  END VCC

  OBS
    LAYER metal1 ;
      POLYGON  0 0
               0 139.5         2.57 139.5         2.57 135.08         20.77 135.08
               20.77 139.5         22.21 139.5         22.21 135.08         40.41 135.08
               40.41 139.5         41.85 139.5         41.85 135.08         60.05 135.08
               60.05 139.5         62.62 139.5         62.62 0         60.05 0
               60.05 3.28         2.57 3.28         2.57 0         0 0 ;
    LAYER via ;
      RECT 42.13 135.36 59.77 139.5 ;
      RECT 2.85 135.36 20.49 139.5 ;
      RECT 2.85 0 59.77 3 ;
      RECT 22.49 135.36 40.13 139.5 ;
    LAYER metal2 ;
      POLYGON  0 0
               0 139.5         2.53 139.5         2.53 135.04         20.81 135.04
               20.81 139.5         22.17 139.5         22.17 135.04         40.45 135.04
               40.45 139.5         41.81 139.5         41.81 135.04         60.09 135.04
               60.09 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via2 ;
      RECT 42.13 135.36 59.77 139.5 ;
      RECT 2.85 135.36 20.49 139.5 ;
      RECT 2.85 0 59.77 3 ;
      RECT 22.49 135.36 40.13 139.5 ;
    LAYER metal3 ;
      POLYGON  0 0
               0 139.5         2.53 139.5         2.53 135.04         20.81 135.04
               20.81 139.5         22.17 139.5         22.17 135.04         40.45 135.04
               40.45 139.5         41.81 139.5         41.81 135.04         60.09 135.04
               60.09 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via3 ;
      RECT 42.13 135.36 59.77 139.5 ;
      RECT 2.85 135.36 20.49 139.5 ;
      RECT 2.85 0 59.77 3 ;
      RECT 22.49 135.36 40.13 139.5 ;
    LAYER metal4 ;
      POLYGON  0 0
               0 139.5         2.53 139.5         2.53 135.04         20.81 135.04
               20.81 139.5         22.17 139.5         22.17 135.04         40.45 135.04
               40.45 139.5         41.81 139.5         41.81 135.04         60.09 135.04
               60.09 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via4 ;
      RECT 42.13 135.36 59.77 139.5 ;
      RECT 2.85 135.36 20.49 139.5 ;
      RECT 22.49 135.36 40.13 139.5 ;
    LAYER metal5 ;
      POLYGON  0 92.26
               0 139.5         2.53 139.5         2.53 135.04         20.81 135.04
               20.81 139.5         22.17 139.5         22.17 135.04         40.45 135.04
               40.45 139.5         41.81 139.5         41.81 135.04         60.09 135.04
               60.09 139.5         62.62 139.5         62.62 92.26         0 92.26 ;
    LAYER via5 ;
      RECT 42.13 135.36 59.77 139.5 ;
      RECT 2.85 135.36 20.49 139.5 ;
      RECT 22.49 135.36 40.13 139.5 ;
    LAYER metal6 ;
      POLYGON  0 92.26
               0 139.5         2.25 139.5         2.25 134.76         21.09 134.76
               21.09 139.5         21.89 139.5         21.89 134.76         40.73 134.76
               40.73 139.5         41.53 139.5         41.53 134.76         60.37 134.76
               60.37 139.5         62.62 139.5         62.62 92.26         0 92.26 ;
  END

END VCCKD

MACRO XMC
  CLASS PAD ;
  FOREIGN XMC 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 34.1 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  PIN PD
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 9.29 234.08 11.17 234.98 ;
    LAYER metal2 ;
      RECT 9.29 234.08 11.17 234.98 ;
    LAYER metal3 ;
      RECT 9.29 234.08 11.17 234.98 ;
    END
  END PD

  PIN PU
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 5.57 234.08 7.45 234.98 ;
    LAYER metal2 ;
      RECT 5.57 234.08 7.45 234.98 ;
    LAYER metal3 ;
      RECT 5.57 234.08 7.45 234.98 ;
    END
  END PU

  PIN I
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 ;
      RECT 1.91 0 32.19 4.3 ;
    END
  END I

  PIN SMT
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 1.85 234.08 3.73 234.98 ;
    LAYER metal2 ;
      RECT 1.85 234.08 3.73 234.98 ;
    LAYER metal3 ;
      RECT 1.85 234.08 3.73 234.98 ;
    END
  END SMT

  PIN O
    DIRECTION OUTPUT ;
    PORT
    LAYER metal1 ;
      RECT 15.49 234.08 17.37 234.98 ;
    LAYER metal2 ;
      RECT 15.49 234.08 17.37 234.98 ;
    LAYER metal3 ;
      RECT 15.49 234.08 17.37 234.98 ;
    END
  END O

  OBS
    LAYER metal1 ;
      POLYGON  0 0
               0 234.98         1.61 234.98         1.61 233.84         3.97 233.84
               3.97 234.98         5.33 234.98         5.33 233.84         7.69 233.84
               7.69 234.98         9.05 234.98         9.05 233.84         11.41 233.84
               11.41 234.98         15.25 234.98         15.25 233.84         17.61 233.84
               17.61 234.98         34.1 234.98         34.1 0         32.47 0
               32.47 4.58         1.63 4.58         1.63 0         0 0 ;
    LAYER via ;
      RECT 5.57 234.08 7.45 234.98 ;
      RECT 1.85 234.08 3.73 234.98 ;
      RECT 9.29 234.08 11.17 234.98 ;
      RECT 15.49 234.08 17.37 234.98 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 ;
      POLYGON  0 0
               0 234.98         1.57 234.98         1.57 233.8         4.01 233.8
               4.01 234.98         5.29 234.98         5.29 233.8         7.73 233.8
               7.73 234.98         9.01 234.98         9.01 233.8         11.45 233.8
               11.45 234.98         15.21 234.98         15.21 233.8         17.65 233.8
               17.65 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via2 ;
      RECT 5.57 234.08 7.45 234.98 ;
      RECT 1.85 234.08 3.73 234.98 ;
      RECT 9.29 234.08 11.17 234.98 ;
      RECT 15.49 234.08 17.37 234.98 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 ;
      POLYGON  0 0
               0 234.98         1.57 234.98         1.57 233.8         4.01 233.8
               4.01 234.98         5.29 234.98         5.29 233.8         7.73 233.8
               7.73 234.98         9.01 234.98         9.01 233.8         11.45 233.8
               11.45 234.98         15.21 234.98         15.21 233.8         17.65 233.8
               17.65 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via3 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 ;
      POLYGON  0 234.98
               34.1 234.98         34.1 0         32.51 0         32.51 4.62
               1.59 4.62         1.59 0         0 0         0 234.98 ;
    LAYER metal5 ;
      RECT 0 155.59 34.1 234.98 ;
    LAYER metal6 ;
      RECT 0 155.59 34.1 234.98 ;
  END

END XMC

MACRO XMD
  CLASS PAD ;
  FOREIGN XMD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 62.62 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  PIN PD
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 33.47 138.6 35.35 139.5 ;
    LAYER metal2 ;
      RECT 33.47 138.6 35.35 139.5 ;
    LAYER metal3 ;
      RECT 33.47 138.6 35.35 139.5 ;
    END
  END PD

  PIN PU
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 27.89 138.6 29.77 139.5 ;
    LAYER metal2 ;
      RECT 27.89 138.6 29.77 139.5 ;
    LAYER metal3 ;
      RECT 27.89 138.6 29.77 139.5 ;
    END
  END PU

  PIN I
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 ;
      RECT 2.85 0 59.77 3 ;
    END
  END I

  PIN SMT
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 23.55 138.6 25.43 139.5 ;
    LAYER metal2 ;
      RECT 23.55 138.6 25.43 139.5 ;
    LAYER metal3 ;
      RECT 23.55 138.6 25.43 139.5 ;
    END
  END SMT

  PIN O
    DIRECTION OUTPUT ;
    PORT
    LAYER metal1 ;
      RECT 39.67 138.6 41.55 139.5 ;
    LAYER metal2 ;
      RECT 39.67 138.6 41.55 139.5 ;
    LAYER metal3 ;
      RECT 39.67 138.6 41.55 139.5 ;
    END
  END O

  OBS
    LAYER metal1 ;
      POLYGON  0 0
               0 139.5         23.31 139.5         23.31 138.36         25.67 138.36
               25.67 139.5         27.65 139.5         27.65 138.36         30.01 138.36
               30.01 139.5         33.23 139.5         33.23 138.36         35.59 138.36
               35.59 139.5         39.43 139.5         39.43 138.36         41.79 138.36
               41.79 139.5         62.62 139.5         62.62 0         60.05 0
               60.05 3.28         2.57 3.28         2.57 0         0 0 ;
    LAYER via ;
      RECT 27.89 138.6 29.77 139.5 ;
      RECT 23.55 138.6 25.43 139.5 ;
      RECT 33.47 138.6 35.35 139.5 ;
      RECT 39.67 138.6 41.55 139.5 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 ;
      POLYGON  0 0
               0 139.5         23.27 139.5         23.27 138.32         25.71 138.32
               25.71 139.5         27.61 139.5         27.61 138.32         30.05 138.32
               30.05 139.5         33.19 139.5         33.19 138.32         35.63 138.32
               35.63 139.5         39.39 139.5         39.39 138.32         41.83 138.32
               41.83 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via2 ;
      RECT 27.89 138.6 29.77 139.5 ;
      RECT 23.55 138.6 25.43 139.5 ;
      RECT 33.47 138.6 35.35 139.5 ;
      RECT 39.67 138.6 41.55 139.5 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 ;
      POLYGON  0 0
               0 139.5         23.27 139.5         23.27 138.32         25.71 138.32
               25.71 139.5         27.61 139.5         27.61 138.32         30.05 138.32
               30.05 139.5         33.19 139.5         33.19 138.32         35.63 138.32
               35.63 139.5         39.39 139.5         39.39 138.32         41.83 138.32
               41.83 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via3 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 ;
      POLYGON  0 139.5
               62.62 139.5         62.62 0         60.09 0         60.09 3.32
               2.53 3.32         2.53 0         0 0         0 139.5 ;
    LAYER metal5 ;
      RECT 0 92.26 62.62 139.5 ;
    LAYER metal6 ;
      RECT 0 92.26 62.62 139.5 ;
  END

END XMD

MACRO YA2GSC
  CLASS PAD ;
  FOREIGN YA2GSC 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 34.1 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  PIN SR
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 30.99 234.08 32.87 234.98 ;
    LAYER metal2 ;
      RECT 30.99 234.08 32.87 234.98 ;
    LAYER metal3 ;
      RECT 30.99 234.08 32.87 234.98 ;
    END
  END SR

  PIN E
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 15.49 234.08 17.37 234.98 ;
    LAYER metal2 ;
      RECT 15.49 234.08 17.37 234.98 ;
    LAYER metal3 ;
      RECT 15.49 234.08 17.37 234.98 ;
    END
  END E

  PIN I
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 27.89 234.08 29.77 234.98 ;
    LAYER metal2 ;
      RECT 27.89 234.08 29.77 234.98 ;
    LAYER metal3 ;
      RECT 27.89 234.08 29.77 234.98 ;
    END
  END I

  PIN O
    DIRECTION OUTPUT ;
    PORT
    LAYER metal1 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 ;
      RECT 1.91 0 32.19 4.3 ;
    END
  END O

  PIN E2
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 18.59 234.08 20.47 234.98 ;
    LAYER metal2 ;
      RECT 18.59 234.08 20.47 234.98 ;
    LAYER metal3 ;
      RECT 18.59 234.08 20.47 234.98 ;
    END
  END E2

  PIN E4
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 24.79 234.08 26.67 234.98 ;
    LAYER metal2 ;
      RECT 24.79 234.08 26.67 234.98 ;
    LAYER metal3 ;
      RECT 24.79 234.08 26.67 234.98 ;
    END
  END E4

  PIN E8
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 21.69 234.08 23.57 234.98 ;
    LAYER metal2 ;
      RECT 21.69 234.08 23.57 234.98 ;
    LAYER metal3 ;
      RECT 21.69 234.08 23.57 234.98 ;
    END
  END E8

  OBS
    LAYER metal1 ;
      POLYGON  0 0
               0 234.98         15.25 234.98         15.25 233.84         17.61 233.84
               17.61 234.98         18.35 234.98         18.35 233.84         20.71 233.84
               20.71 234.98         21.45 234.98         21.45 233.84         23.81 233.84
               23.81 234.98         24.55 234.98         24.55 233.84         26.91 233.84
               26.91 234.98         27.65 234.98         27.65 233.84         30.01 233.84
               30.01 234.98         30.75 234.98         30.75 233.84         33.11 233.84
               33.11 234.98         34.1 234.98         34.1 0         32.47 0
               32.47 4.58         1.63 4.58         1.63 0         0 0 ;
    LAYER via ;
      RECT 18.59 234.08 20.47 234.98 ;
      RECT 21.69 234.08 23.57 234.98 ;
      RECT 24.79 234.08 26.67 234.98 ;
      RECT 30.99 234.08 32.87 234.98 ;
      RECT 27.89 234.08 29.77 234.98 ;
      RECT 15.49 234.08 17.37 234.98 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 ;
      POLYGON  0 0
               0 234.98         15.21 234.98         15.21 233.8         17.65 233.8
               17.65 234.98         18.31 234.98         18.31 233.8         20.75 233.8
               20.75 234.98         21.41 234.98         21.41 233.8         23.85 233.8
               23.85 234.98         24.51 234.98         24.51 233.8         26.95 233.8
               26.95 234.98         27.61 234.98         27.61 233.8         30.05 233.8
               30.05 234.98         30.71 234.98         30.71 233.8         33.15 233.8
               33.15 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via2 ;
      RECT 18.59 234.08 20.47 234.98 ;
      RECT 21.69 234.08 23.57 234.98 ;
      RECT 24.79 234.08 26.67 234.98 ;
      RECT 30.99 234.08 32.87 234.98 ;
      RECT 27.89 234.08 29.77 234.98 ;
      RECT 15.49 234.08 17.37 234.98 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 ;
      POLYGON  0 0
               0 234.98         15.21 234.98         15.21 233.8         17.65 233.8
               17.65 234.98         18.31 234.98         18.31 233.8         20.75 233.8
               20.75 234.98         21.41 234.98         21.41 233.8         23.85 233.8
               23.85 234.98         24.51 234.98         24.51 233.8         26.95 233.8
               26.95 234.98         27.61 234.98         27.61 233.8         30.05 233.8
               30.05 234.98         30.71 234.98         30.71 233.8         33.15 233.8
               33.15 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via3 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 ;
      POLYGON  0 234.98
               34.1 234.98         34.1 0         32.51 0         32.51 4.62
               1.59 4.62         1.59 0         0 0         0 234.98 ;
    LAYER metal5 ;
      RECT 0 155.59 34.1 234.98 ;
    LAYER metal6 ;
      RECT 0 155.59 34.1 234.98 ;
  END

END YA2GSC

MACRO YA2GSD
  CLASS PAD ;
  FOREIGN YA2GSD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 62.62 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  PIN SR
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 27.89 138.6 29.77 139.5 ;
    LAYER metal2 ;
      RECT 27.89 138.6 29.77 139.5 ;
    LAYER metal3 ;
      RECT 27.89 138.6 29.77 139.5 ;
    END
  END SR

  PIN E
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 33.47 138.6 35.35 139.5 ;
    LAYER metal2 ;
      RECT 33.47 138.6 35.35 139.5 ;
    LAYER metal3 ;
      RECT 33.47 138.6 35.35 139.5 ;
    END
  END E

  PIN I
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 24.17 138.6 26.05 139.5 ;
    LAYER metal2 ;
      RECT 24.17 138.6 26.05 139.5 ;
    LAYER metal3 ;
      RECT 24.17 138.6 26.05 139.5 ;
    END
  END I

  PIN O
    DIRECTION OUTPUT ;
    PORT
    LAYER metal1 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 ;
      RECT 2.85 0 59.77 3 ;
    END
  END O

  PIN E2
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 14.25 138.6 16.13 139.5 ;
    LAYER metal2 ;
      RECT 14.25 138.6 16.13 139.5 ;
    LAYER metal3 ;
      RECT 14.25 138.6 16.13 139.5 ;
    END
  END E2

  PIN E4
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 20.45 138.6 22.33 139.5 ;
    LAYER metal2 ;
      RECT 20.45 138.6 22.33 139.5 ;
    LAYER metal3 ;
      RECT 20.45 138.6 22.33 139.5 ;
    END
  END E4

  PIN E8
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 17.35 138.6 19.23 139.5 ;
    LAYER metal2 ;
      RECT 17.35 138.6 19.23 139.5 ;
    LAYER metal3 ;
      RECT 17.35 138.6 19.23 139.5 ;
    END
  END E8

  OBS
    LAYER metal1 ;
      POLYGON  0 0
               0 139.5         14.01 139.5         14.01 138.36         16.37 138.36
               16.37 139.5         17.11 139.5         17.11 138.36         19.47 138.36
               19.47 139.5         20.21 139.5         20.21 138.36         22.57 138.36
               22.57 139.5         23.93 139.5         23.93 138.36         26.29 138.36
               26.29 139.5         27.65 139.5         27.65 138.36         30.01 138.36
               30.01 139.5         33.23 139.5         33.23 138.36         35.59 138.36
               35.59 139.5         62.62 139.5         62.62 0         60.05 0
               60.05 3.28         2.57 3.28         2.57 0         0 0 ;
    LAYER via ;
      RECT 24.17 138.6 26.05 139.5 ;
      RECT 20.45 138.6 22.33 139.5 ;
      RECT 33.47 138.6 35.35 139.5 ;
      RECT 27.89 138.6 29.77 139.5 ;
      RECT 17.35 138.6 19.23 139.5 ;
      RECT 14.25 138.6 16.13 139.5 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 ;
      POLYGON  0 0
               0 139.5         13.97 139.5         13.97 138.32         16.41 138.32
               16.41 139.5         17.07 139.5         17.07 138.32         19.51 138.32
               19.51 139.5         20.17 139.5         20.17 138.32         22.61 138.32
               22.61 139.5         23.89 139.5         23.89 138.32         26.33 138.32
               26.33 139.5         27.61 139.5         27.61 138.32         30.05 138.32
               30.05 139.5         33.19 139.5         33.19 138.32         35.63 138.32
               35.63 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via2 ;
      RECT 24.17 138.6 26.05 139.5 ;
      RECT 20.45 138.6 22.33 139.5 ;
      RECT 33.47 138.6 35.35 139.5 ;
      RECT 27.89 138.6 29.77 139.5 ;
      RECT 17.35 138.6 19.23 139.5 ;
      RECT 14.25 138.6 16.13 139.5 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 ;
      POLYGON  0 0
               0 139.5         13.97 139.5         13.97 138.32         16.41 138.32
               16.41 139.5         17.07 139.5         17.07 138.32         19.51 138.32
               19.51 139.5         20.17 139.5         20.17 138.32         22.61 138.32
               22.61 139.5         23.89 139.5         23.89 138.32         26.33 138.32
               26.33 139.5         27.61 139.5         27.61 138.32         30.05 138.32
               30.05 139.5         33.19 139.5         33.19 138.32         35.63 138.32
               35.63 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via3 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 ;
      POLYGON  0 139.5
               62.62 139.5         62.62 0         60.09 0         60.09 3.32
               2.53 3.32         2.53 0         0 0         0 139.5 ;
    LAYER metal5 ;
      RECT 0 92.26 62.62 139.5 ;
    LAYER metal6 ;
      RECT 0 92.26 62.62 139.5 ;
  END

END YA2GSD

MACRO ZMA2GSC
  CLASS PAD ;
  FOREIGN ZMA2GSC 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 34.1 BY 235.6 ;
  SYMMETRY X Y R90 ;
  SITE iocore_c ;

  PIN PD
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 9.29 234.08 11.17 234.98 ;
    LAYER metal2 ;
      RECT 9.29 234.08 11.17 234.98 ;
    LAYER metal3 ;
      RECT 9.29 234.08 11.17 234.98 ;
    END
  END PD

  PIN PU
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 5.57 234.08 7.45 234.98 ;
    LAYER metal2 ;
      RECT 5.57 234.08 7.45 234.98 ;
    LAYER metal3 ;
      RECT 5.57 234.08 7.45 234.98 ;
    END
  END PU

  PIN SR
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 30.99 234.08 32.87 234.98 ;
    LAYER metal2 ;
      RECT 30.99 234.08 32.87 234.98 ;
    LAYER metal3 ;
      RECT 30.99 234.08 32.87 234.98 ;
    END
  END SR

  PIN E
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 12.39 234.08 14.27 234.98 ;
    LAYER metal2 ;
      RECT 12.39 234.08 14.27 234.98 ;
    LAYER metal3 ;
      RECT 12.39 234.08 14.27 234.98 ;
    END
  END E

  PIN I
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 27.89 234.08 29.77 234.98 ;
    LAYER metal2 ;
      RECT 27.89 234.08 29.77 234.98 ;
    LAYER metal3 ;
      RECT 27.89 234.08 29.77 234.98 ;
    END
  END I

  PIN SMT
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 1.85 234.08 3.73 234.98 ;
    LAYER metal2 ;
      RECT 1.85 234.08 3.73 234.98 ;
    LAYER metal3 ;
      RECT 1.85 234.08 3.73 234.98 ;
    END
  END SMT

  PIN O
    DIRECTION OUTPUT ;
    PORT
    LAYER metal1 ;
      RECT 15.49 234.08 17.37 234.98 ;
    LAYER metal2 ;
      RECT 15.49 234.08 17.37 234.98 ;
    LAYER metal3 ;
      RECT 15.49 234.08 17.37 234.98 ;
    END
  END O

  PIN E2
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 18.59 234.08 20.47 234.98 ;
    LAYER metal2 ;
      RECT 18.59 234.08 20.47 234.98 ;
    LAYER metal3 ;
      RECT 18.59 234.08 20.47 234.98 ;
    END
  END E2

  PIN E4
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 24.79 234.08 26.67 234.98 ;
    LAYER metal2 ;
      RECT 24.79 234.08 26.67 234.98 ;
    LAYER metal3 ;
      RECT 24.79 234.08 26.67 234.98 ;
    END
  END E4

  PIN E8
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 21.69 234.08 23.57 234.98 ;
    LAYER metal2 ;
      RECT 21.69 234.08 23.57 234.98 ;
    LAYER metal3 ;
      RECT 21.69 234.08 23.57 234.98 ;
    END
  END E8

  PIN IO
    DIRECTION INOUT ;
    PORT
    LAYER metal1 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 ;
      RECT 1.91 0 32.19 4.3 ;
    END
  END IO

  OBS
    LAYER metal1 ;
      POLYGON  0 0
               0 234.98         1.61 234.98         1.61 233.84         3.97 233.84
               3.97 234.98         5.33 234.98         5.33 233.84         7.69 233.84
               7.69 234.98         9.05 234.98         9.05 233.84         11.41 233.84
               11.41 234.98         12.15 234.98         12.15 233.84         14.51 233.84
               14.51 234.98         15.25 234.98         15.25 233.84         17.61 233.84
               17.61 234.98         18.35 234.98         18.35 233.84         20.71 233.84
               20.71 234.98         21.45 234.98         21.45 233.84         23.81 233.84
               23.81 234.98         24.55 234.98         24.55 233.84         26.91 233.84
               26.91 234.98         27.65 234.98         27.65 233.84         30.01 233.84
               30.01 234.98         30.75 234.98         30.75 233.84         33.11 233.84
               33.11 234.98         34.1 234.98         34.1 0         32.47 0
               32.47 4.58         1.63 4.58         1.63 0         0 0 ;
    LAYER via ;
      RECT 27.89 234.08 29.77 234.98 ;
      RECT 1.85 234.08 3.73 234.98 ;
      RECT 30.99 234.08 32.87 234.98 ;
      RECT 12.39 234.08 14.27 234.98 ;
      RECT 24.79 234.08 26.67 234.98 ;
      RECT 9.29 234.08 11.17 234.98 ;
      RECT 15.49 234.08 17.37 234.98 ;
      RECT 21.69 234.08 23.57 234.98 ;
      RECT 18.59 234.08 20.47 234.98 ;
      RECT 5.57 234.08 7.45 234.98 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal2 ;
      POLYGON  0 0
               0 234.98         1.57 234.98         1.57 233.8         4.01 233.8
               4.01 234.98         5.29 234.98         5.29 233.8         7.73 233.8
               7.73 234.98         9.01 234.98         9.01 233.8         11.45 233.8
               11.45 234.98         12.11 234.98         12.11 233.8         14.55 233.8
               14.55 234.98         15.21 234.98         15.21 233.8         17.65 233.8
               17.65 234.98         18.31 234.98         18.31 233.8         20.75 233.8
               20.75 234.98         21.41 234.98         21.41 233.8         23.85 233.8
               23.85 234.98         24.51 234.98         24.51 233.8         26.95 233.8
               26.95 234.98         27.61 234.98         27.61 233.8         30.05 233.8
               30.05 234.98         30.71 234.98         30.71 233.8         33.15 233.8
               33.15 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via2 ;
      RECT 27.89 234.08 29.77 234.98 ;
      RECT 1.85 234.08 3.73 234.98 ;
      RECT 30.99 234.08 32.87 234.98 ;
      RECT 12.39 234.08 14.27 234.98 ;
      RECT 24.79 234.08 26.67 234.98 ;
      RECT 9.29 234.08 11.17 234.98 ;
      RECT 15.49 234.08 17.37 234.98 ;
      RECT 21.69 234.08 23.57 234.98 ;
      RECT 18.59 234.08 20.47 234.98 ;
      RECT 5.57 234.08 7.45 234.98 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal3 ;
      POLYGON  0 0
               0 234.98         1.57 234.98         1.57 233.8         4.01 233.8
               4.01 234.98         5.29 234.98         5.29 233.8         7.73 233.8
               7.73 234.98         9.01 234.98         9.01 233.8         11.45 233.8
               11.45 234.98         12.11 234.98         12.11 233.8         14.55 233.8
               14.55 234.98         15.21 234.98         15.21 233.8         17.65 233.8
               17.65 234.98         18.31 234.98         18.31 233.8         20.75 233.8
               20.75 234.98         21.41 234.98         21.41 233.8         23.85 233.8
               23.85 234.98         24.51 234.98         24.51 233.8         26.95 233.8
               26.95 234.98         27.61 234.98         27.61 233.8         30.05 233.8
               30.05 234.98         30.71 234.98         30.71 233.8         33.15 233.8
               33.15 234.98         34.1 234.98         34.1 0         32.51 0
               32.51 4.62         1.59 4.62         1.59 0         0 0 ;
    LAYER via3 ;
      RECT 1.91 0 32.19 4.3 ;
    LAYER metal4 ;
      POLYGON  0 234.98
               34.1 234.98         34.1 0         32.51 0         32.51 4.62
               1.59 4.62         1.59 0         0 0         0 234.98 ;
    LAYER metal5 ;
      RECT 0 155.59 34.1 234.98 ;
    LAYER metal6 ;
      RECT 0 155.59 34.1 234.98 ;
  END

END ZMA2GSC

MACRO ZMA2GSD
  CLASS PAD ;
  FOREIGN ZMA2GSD 0.000 0.000 ;
  ORIGIN 0 0 ;
  SIZE 62.62 BY 140.12 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;

  PIN PD
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 11.77 138.6 13.65 139.5 ;
    LAYER metal2 ;
      RECT 11.77 138.6 13.65 139.5 ;
    LAYER metal3 ;
      RECT 11.77 138.6 13.65 139.5 ;
    END
  END PD

  PIN PU
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 6.19 138.6 8.07 139.5 ;
    LAYER metal2 ;
      RECT 6.19 138.6 8.07 139.5 ;
    LAYER metal3 ;
      RECT 6.19 138.6 8.07 139.5 ;
    END
  END PU

  PIN SR
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 35.95 138.6 37.83 139.5 ;
    LAYER metal2 ;
      RECT 35.95 138.6 37.83 139.5 ;
    LAYER metal3 ;
      RECT 35.95 138.6 37.83 139.5 ;
    END
  END SR

  PIN E
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 41.53 138.6 43.41 139.5 ;
    LAYER metal2 ;
      RECT 41.53 138.6 43.41 139.5 ;
    LAYER metal3 ;
      RECT 41.53 138.6 43.41 139.5 ;
    END
  END E

  PIN I
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 32.23 138.6 34.11 139.5 ;
    LAYER metal2 ;
      RECT 32.23 138.6 34.11 139.5 ;
    LAYER metal3 ;
      RECT 32.23 138.6 34.11 139.5 ;
    END
  END I

  PIN SMT
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 1.85 138.6 3.73 139.5 ;
    LAYER metal2 ;
      RECT 1.85 138.6 3.73 139.5 ;
    LAYER metal3 ;
      RECT 1.85 138.6 3.73 139.5 ;
    END
  END SMT

  PIN O
    DIRECTION OUTPUT ;
    PORT
    LAYER metal1 ;
      RECT 17.97 138.6 19.85 139.5 ;
    LAYER metal2 ;
      RECT 17.97 138.6 19.85 139.5 ;
    LAYER metal3 ;
      RECT 17.97 138.6 19.85 139.5 ;
    END
  END O

  PIN E2
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 22.31 138.6 24.19 139.5 ;
    LAYER metal2 ;
      RECT 22.31 138.6 24.19 139.5 ;
    LAYER metal3 ;
      RECT 22.31 138.6 24.19 139.5 ;
    END
  END E2

  PIN E4
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 28.51 138.6 30.39 139.5 ;
    LAYER metal2 ;
      RECT 28.51 138.6 30.39 139.5 ;
    LAYER metal3 ;
      RECT 28.51 138.6 30.39 139.5 ;
    END
  END E4

  PIN E8
    DIRECTION INPUT ;
    PORT
    LAYER metal1 ;
      RECT 25.41 138.6 27.29 139.5 ;
    LAYER metal2 ;
      RECT 25.41 138.6 27.29 139.5 ;
    LAYER metal3 ;
      RECT 25.41 138.6 27.29 139.5 ;
    END
  END E8

  PIN IO
    DIRECTION INOUT ;
    PORT
    LAYER metal1 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 ;
      RECT 2.85 0 59.77 3 ;
    END
  END IO

  OBS
    LAYER metal1 ;
      POLYGON  0 0
               0 139.5         1.61 139.5         1.61 138.36         3.97 138.36
               3.97 139.5         5.95 139.5         5.95 138.36         8.31 138.36
               8.31 139.5         11.53 139.5         11.53 138.36         13.89 138.36
               13.89 139.5         17.73 139.5         17.73 138.36         20.09 138.36
               20.09 139.5         22.07 139.5         22.07 138.36         24.43 138.36
               24.43 139.5         25.17 139.5         25.17 138.36         27.53 138.36
               27.53 139.5         28.27 139.5         28.27 138.36         30.63 138.36
               30.63 139.5         31.99 139.5         31.99 138.36         34.35 138.36
               34.35 139.5         35.71 139.5         35.71 138.36         38.07 138.36
               38.07 139.5         41.29 139.5         41.29 138.36         43.65 138.36
               43.65 139.5         62.62 139.5         62.62 0         60.05 0
               60.05 3.28         2.57 3.28         2.57 0         0 0 ;
    LAYER via ;
      RECT 22.31 138.6 24.19 139.5 ;
      RECT 25.41 138.6 27.29 139.5 ;
      RECT 35.95 138.6 37.83 139.5 ;
      RECT 1.85 138.6 3.73 139.5 ;
      RECT 41.53 138.6 43.41 139.5 ;
      RECT 11.77 138.6 13.65 139.5 ;
      RECT 17.97 138.6 19.85 139.5 ;
      RECT 28.51 138.6 30.39 139.5 ;
      RECT 32.23 138.6 34.11 139.5 ;
      RECT 6.19 138.6 8.07 139.5 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal2 ;
      POLYGON  0 0
               0 139.5         1.57 139.5         1.57 138.32         4.01 138.32
               4.01 139.5         5.91 139.5         5.91 138.32         8.35 138.32
               8.35 139.5         11.49 139.5         11.49 138.32         13.93 138.32
               13.93 139.5         17.69 139.5         17.69 138.32         20.13 138.32
               20.13 139.5         22.03 139.5         22.03 138.32         24.47 138.32
               24.47 139.5         25.13 139.5         25.13 138.32         27.57 138.32
               27.57 139.5         28.23 139.5         28.23 138.32         30.67 138.32
               30.67 139.5         31.95 139.5         31.95 138.32         34.39 138.32
               34.39 139.5         35.67 139.5         35.67 138.32         38.11 138.32
               38.11 139.5         41.25 139.5         41.25 138.32         43.69 138.32
               43.69 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via2 ;
      RECT 22.31 138.6 24.19 139.5 ;
      RECT 25.41 138.6 27.29 139.5 ;
      RECT 35.95 138.6 37.83 139.5 ;
      RECT 1.85 138.6 3.73 139.5 ;
      RECT 41.53 138.6 43.41 139.5 ;
      RECT 11.77 138.6 13.65 139.5 ;
      RECT 17.97 138.6 19.85 139.5 ;
      RECT 28.51 138.6 30.39 139.5 ;
      RECT 32.23 138.6 34.11 139.5 ;
      RECT 6.19 138.6 8.07 139.5 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal3 ;
      POLYGON  0 0
               0 139.5         1.57 139.5         1.57 138.32         4.01 138.32
               4.01 139.5         5.91 139.5         5.91 138.32         8.35 138.32
               8.35 139.5         11.49 139.5         11.49 138.32         13.93 138.32
               13.93 139.5         17.69 139.5         17.69 138.32         20.13 138.32
               20.13 139.5         22.03 139.5         22.03 138.32         24.47 138.32
               24.47 139.5         25.13 139.5         25.13 138.32         27.57 138.32
               27.57 139.5         28.23 139.5         28.23 138.32         30.67 138.32
               30.67 139.5         31.95 139.5         31.95 138.32         34.39 138.32
               34.39 139.5         35.67 139.5         35.67 138.32         38.11 138.32
               38.11 139.5         41.25 139.5         41.25 138.32         43.69 138.32
               43.69 139.5         62.62 139.5         62.62 0         60.09 0
               60.09 3.32         2.53 3.32         2.53 0         0 0 ;
    LAYER via3 ;
      RECT 2.85 0 59.77 3 ;
    LAYER metal4 ;
      POLYGON  0 139.5
               62.62 139.5         62.62 0         60.09 0         60.09 3.32
               2.53 3.32         2.53 0         0 0         0 139.5 ;
    LAYER metal5 ;
      RECT 0 92.26 62.62 139.5 ;
    LAYER metal6 ;
      RECT 0 92.26 62.62 139.5 ;
  END

END ZMA2GSD

END LIBRARY
